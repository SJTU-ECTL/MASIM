module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 ;
  assign n25 = ( ~x0 & x1 ) | ( ~x0 & x2 ) | ( x1 & x2 ) ;
  assign n26 = ~x1 & n25 ;
  assign n27 = ~x0 & x1 ;
  assign n28 = n27 ^ n26 ^ x0 ;
  assign n29 = x3 | n28 ;
  assign n30 = x4 | n29 ;
  assign n31 = x5 | n30 ;
  assign n32 = x6 | n31 ;
  assign n33 = x7 | n32 ;
  assign n34 = x8 | n33 ;
  assign n35 = x9 | n34 ;
  assign n36 = x10 | n35 ;
  assign n37 = x22 & n35 ;
  assign n38 = n37 ^ n35 ^ x10 ;
  assign n39 = x22 & n32 ;
  assign n40 = ~x22 & n36 ;
  assign n41 = x11 | n36 ;
  assign n42 = x12 | n41 ;
  assign n43 = x22 & n31 ;
  assign n44 = n39 ^ n32 ^ x7 ;
  assign n45 = x13 | n42 ;
  assign n46 = x14 | n45 ;
  assign n47 = x15 | n46 ;
  assign n48 = x22 & n41 ;
  assign n49 = x22 & n29 ;
  assign n50 = x16 | n47 ;
  assign n51 = x22 & n42 ;
  assign n52 = n43 ^ n31 ^ x6 ;
  assign n53 = x22 & n50 ;
  assign n54 = x22 & n47 ;
  assign n55 = x17 | n50 ;
  assign n56 = n51 ^ n42 ^ x13 ;
  assign n57 = x22 & n55 ;
  assign n58 = x18 | n55 ;
  assign n59 = x22 & n58 ;
  assign n60 = n59 ^ n58 ^ x19 ;
  assign n61 = x19 | n58 ;
  assign n62 = n57 ^ n55 ^ x18 ;
  assign n63 = n60 & ~n62 ;
  assign n64 = n60 | n62 ;
  assign n65 = x22 & n61 ;
  assign n66 = x20 | n61 ;
  assign n67 = ~n60 & n62 ;
  assign n68 = n60 & n62 ;
  assign n69 = x22 & n66 ;
  assign n70 = n49 ^ n29 ^ x4 ;
  assign n71 = n53 ^ n50 ^ x17 ;
  assign n72 = n54 ^ n47 ^ x16 ;
  assign n73 = ~n71 & n72 ;
  assign n74 = n63 & n73 ;
  assign n75 = n48 ^ n41 ^ x12 ;
  assign n76 = n71 & ~n72 ;
  assign n77 = x22 & n34 ;
  assign n78 = n63 & n76 ;
  assign n79 = n77 ^ n34 ^ x9 ;
  assign n80 = x22 & n28 ;
  assign n81 = n65 ^ n61 ^ x20 ;
  assign n82 = ~x22 & n45 ;
  assign n83 = x22 & n46 ;
  assign n84 = n80 ^ n28 ^ x3 ;
  assign n85 = n83 ^ n46 ^ x15 ;
  assign n86 = n69 ^ n66 ^ x21 ;
  assign n87 = n71 | n72 ;
  assign n88 = n71 & n72 ;
  assign n89 = n63 & n88 ;
  assign n90 = n68 & n88 ;
  assign n91 = n63 & ~n87 ;
  assign n92 = n81 | n86 ;
  assign n93 = n81 & ~n86 ;
  assign n94 = n85 & ~n92 ;
  assign n95 = n67 & n88 ;
  assign n96 = ~n64 & n76 ;
  assign n97 = ~n81 & n86 ;
  assign n98 = n85 & n97 ;
  assign n99 = n85 | n92 ;
  assign n100 = ( n93 & n98 ) | ( n93 & n99 ) | ( n98 & n99 ) ;
  assign n101 = n94 & n96 ;
  assign n102 = n68 & ~n87 ;
  assign n103 = n67 & n76 ;
  assign n104 = n67 & n73 ;
  assign n105 = ~n85 & n93 ;
  assign n106 = n64 | n87 ;
  assign n107 = n68 & n76 ;
  assign n108 = n99 | n106 ;
  assign n109 = ( ~n100 & n106 ) | ( ~n100 & n108 ) | ( n106 & n108 ) ;
  assign n110 = ~n99 & n107 ;
  assign n111 = n101 | n110 ;
  assign n112 = n67 & ~n87 ;
  assign n113 = ~n64 & n73 ;
  assign n114 = n74 & n105 ;
  assign n115 = n78 & n105 ;
  assign n116 = ~n64 & n88 ;
  assign n117 = n98 & n116 ;
  assign n118 = ( n109 & n114 ) | ( n109 & ~n117 ) | ( n114 & ~n117 ) ;
  assign n119 = n81 & n86 ;
  assign n120 = ~n85 & n97 ;
  assign n121 = n68 & n73 ;
  assign n122 = n103 & n120 ;
  assign n123 = ~n114 & n118 ;
  assign n124 = ( n76 & n111 ) | ( n76 & n122 ) | ( n111 & n122 ) ;
  assign n125 = n94 & n95 ;
  assign n126 = n94 & n102 ;
  assign n127 = ( ~n115 & n123 ) | ( ~n115 & n126 ) | ( n123 & n126 ) ;
  assign n128 = ( ~n125 & n126 ) | ( ~n125 & n127 ) | ( n126 & n127 ) ;
  assign n129 = ~n126 & n128 ;
  assign n130 = n85 & n119 ;
  assign n131 = ~n90 & n93 ;
  assign n132 = n104 & n130 ;
  assign n133 = n95 & ~n99 ;
  assign n134 = ~n99 & n116 ;
  assign n135 = n96 & n98 ;
  assign n136 = n96 & ~n99 ;
  assign n137 = ~n99 & n104 ;
  assign n138 = n113 & n120 ;
  assign n139 = n89 & n130 ;
  assign n140 = ( n97 & n107 ) | ( n97 & n139 ) | ( n107 & n139 ) ;
  assign n141 = n102 & n130 ;
  assign n142 = ( ~n139 & n140 ) | ( ~n139 & n141 ) | ( n140 & n141 ) ;
  assign n143 = n104 & n120 ;
  assign n144 = ( n137 & ~n138 ) | ( n137 & n143 ) | ( ~n138 & n143 ) ;
  assign n145 = n139 | n142 ;
  assign n146 = n74 & n98 ;
  assign n147 = n89 & n120 ;
  assign n148 = n98 & n113 ;
  assign n149 = n134 | n148 ;
  assign n150 = ( ~n135 & n146 ) | ( ~n135 & n149 ) | ( n146 & n149 ) ;
  assign n151 = n135 | n150 ;
  assign n152 = ( ~n132 & n147 ) | ( ~n132 & n151 ) | ( n147 & n151 ) ;
  assign n153 = n132 | n152 ;
  assign n154 = ( n93 & ~n131 ) | ( n93 & n153 ) | ( ~n131 & n153 ) ;
  assign n155 = ( n133 & ~n136 ) | ( n133 & n154 ) | ( ~n136 & n154 ) ;
  assign n156 = n136 | n155 ;
  assign n157 = n125 | n139 ;
  assign n158 = n85 & n93 ;
  assign n159 = n102 & n158 ;
  assign n160 = n96 & n105 ;
  assign n161 = ~n85 & n119 ;
  assign n162 = n138 | n144 ;
  assign n163 = n102 & n161 ;
  assign n164 = n89 & n93 ;
  assign n165 = ( ~n126 & n160 ) | ( ~n126 & n162 ) | ( n160 & n162 ) ;
  assign n166 = n126 | n165 ;
  assign n167 = ( ~n92 & n102 ) | ( ~n92 & n159 ) | ( n102 & n159 ) ;
  assign n168 = n78 & n97 ;
  assign n169 = ( ~n122 & n143 ) | ( ~n122 & n157 ) | ( n143 & n157 ) ;
  assign n170 = n90 & n120 ;
  assign n171 = n122 | n169 ;
  assign n172 = ( n145 & ~n163 ) | ( n145 & n170 ) | ( ~n163 & n170 ) ;
  assign n173 = n98 & n112 ;
  assign n174 = ~n106 & n161 ;
  assign n175 = n96 & n120 ;
  assign n176 = n91 & n94 ;
  assign n177 = n74 & n130 ;
  assign n178 = n113 & n130 ;
  assign n179 = n107 & n120 ;
  assign n180 = n91 & n105 ;
  assign n181 = ~n106 & n120 ;
  assign n182 = n116 & n130 ;
  assign n183 = n89 & n105 ;
  assign n184 = n121 & n161 ;
  assign n185 = n176 | n177 ;
  assign n186 = n174 | n179 ;
  assign n187 = n105 & n113 ;
  assign n188 = n91 & n98 ;
  assign n189 = n90 & n161 ;
  assign n190 = n78 & n98 ;
  assign n191 = ( n173 & ~n178 ) | ( n173 & n190 ) | ( ~n178 & n190 ) ;
  assign n192 = n182 | n185 ;
  assign n193 = ( ~n181 & n186 ) | ( ~n181 & n192 ) | ( n186 & n192 ) ;
  assign n194 = n178 | n191 ;
  assign n195 = n181 | n193 ;
  assign n196 = n184 | n188 ;
  assign n197 = ( ~n183 & n189 ) | ( ~n183 & n194 ) | ( n189 & n194 ) ;
  assign n198 = ( ~n135 & n137 ) | ( ~n135 & n196 ) | ( n137 & n196 ) ;
  assign n199 = n135 | n198 ;
  assign n200 = n183 | n197 ;
  assign n201 = ( ~n195 & n199 ) | ( ~n195 & n200 ) | ( n199 & n200 ) ;
  assign n202 = n195 | n201 ;
  assign n203 = n89 & n158 ;
  assign n204 = ( ~n175 & n202 ) | ( ~n175 & n203 ) | ( n202 & n203 ) ;
  assign n205 = n175 | n204 ;
  assign n206 = n163 | n172 ;
  assign n207 = ( n180 & ~n187 ) | ( n180 & n205 ) | ( ~n187 & n205 ) ;
  assign n208 = n187 | n207 ;
  assign n209 = ( ~n110 & n160 ) | ( ~n110 & n208 ) | ( n160 & n208 ) ;
  assign n210 = n110 | n209 ;
  assign n211 = n105 & n121 ;
  assign n212 = n89 & n98 ;
  assign n213 = n105 & n112 ;
  assign n214 = n211 | n213 ;
  assign n215 = n179 | n212 ;
  assign n216 = n74 & n120 ;
  assign n217 = n90 & n158 ;
  assign n218 = n170 | n174 ;
  assign n219 = n216 | n218 ;
  assign n220 = n102 & n105 ;
  assign n221 = ~n99 & n121 ;
  assign n222 = ~n99 & n102 ;
  assign n223 = ( n200 & ~n211 ) | ( n200 & n212 ) | ( ~n211 & n212 ) ;
  assign n224 = n102 & n120 ;
  assign n225 = n217 | n221 ;
  assign n226 = n224 | n225 ;
  assign n227 = n98 & n102 ;
  assign n228 = ( n166 & n215 ) | ( n166 & ~n226 ) | ( n215 & ~n226 ) ;
  assign n229 = n113 & n161 ;
  assign n230 = n94 & ~n106 ;
  assign n231 = n96 & n158 ;
  assign n232 = n147 | n222 ;
  assign n233 = n94 & n113 ;
  assign n234 = ~n106 & n130 ;
  assign n235 = n78 & ~n99 ;
  assign n236 = n226 | n228 ;
  assign n237 = n113 & n158 ;
  assign n238 = ~n99 & n113 ;
  assign n239 = ( ~n183 & n231 ) | ( ~n183 & n236 ) | ( n231 & n236 ) ;
  assign n240 = ( ~n122 & n219 ) | ( ~n122 & n234 ) | ( n219 & n234 ) ;
  assign n241 = n122 | n240 ;
  assign n242 = ( ~n178 & n232 ) | ( ~n178 & n241 ) | ( n232 & n241 ) ;
  assign n243 = ( n182 & n214 ) | ( n182 & ~n229 ) | ( n214 & ~n229 ) ;
  assign n244 = n229 | n243 ;
  assign n245 = ( ~n174 & n222 ) | ( ~n174 & n244 ) | ( n222 & n244 ) ;
  assign n246 = n174 | n245 ;
  assign n247 = ( n230 & ~n235 ) | ( n230 & n246 ) | ( ~n235 & n246 ) ;
  assign n248 = n183 | n239 ;
  assign n249 = n178 | n242 ;
  assign n250 = n235 | n247 ;
  assign n251 = ( n133 & ~n233 ) | ( n133 & n249 ) | ( ~n233 & n249 ) ;
  assign n252 = ( n134 & ~n233 ) | ( n134 & n248 ) | ( ~n233 & n248 ) ;
  assign n253 = n211 | n223 ;
  assign n254 = n98 & n107 ;
  assign n255 = n91 & n120 ;
  assign n256 = n254 | n255 ;
  assign n257 = n108 & ~n233 ;
  assign n258 = n103 & n105 ;
  assign n259 = n125 | n258 ;
  assign n260 = ( n78 & n158 ) | ( n78 & n217 ) | ( n158 & n217 ) ;
  assign n261 = n89 & n94 ;
  assign n262 = n98 & n121 ;
  assign n263 = n235 | n256 ;
  assign n264 = n120 & n121 ;
  assign n265 = n264 ^ n262 ^ n261 ;
  assign n266 = n74 & n161 ;
  assign n267 = n216 | n262 ;
  assign n268 = n266 | n267 ;
  assign n269 = n263 | n265 ;
  assign n270 = n78 & n161 ;
  assign n271 = n98 & n104 ;
  assign n272 = n105 & n107 ;
  assign n273 = n116 & n120 ;
  assign n274 = n184 | n272 ;
  assign n275 = n138 | n272 ;
  assign n276 = n173 | n271 ;
  assign n277 = ( n251 & n257 ) | ( n251 & ~n269 ) | ( n257 & ~n269 ) ;
  assign n278 = ~n251 & n277 ;
  assign n279 = ( ~n212 & n276 ) | ( ~n212 & n278 ) | ( n276 & n278 ) ;
  assign n280 = ~n276 & n279 ;
  assign n281 = ( n260 & ~n273 ) | ( n260 & n275 ) | ( ~n273 & n275 ) ;
  assign n282 = ( ~n188 & n238 ) | ( ~n188 & n280 ) | ( n238 & n280 ) ;
  assign n283 = ( n95 & n119 ) | ( n95 & n274 ) | ( n119 & n274 ) ;
  assign n284 = n233 | n261 ;
  assign n285 = ( n180 & ~n259 ) | ( n180 & n284 ) | ( ~n259 & n284 ) ;
  assign n286 = n259 | n285 ;
  assign n287 = n227 | n270 ;
  assign n288 = ( n268 & n286 ) | ( n268 & ~n287 ) | ( n286 & ~n287 ) ;
  assign n289 = n287 | n288 ;
  assign n290 = n95 & n98 ;
  assign n291 = ~n238 & n282 ;
  assign n292 = ( n254 & n289 ) | ( n254 & ~n290 ) | ( n289 & ~n290 ) ;
  assign n293 = n290 | n292 ;
  assign n294 = ( ~n213 & n272 ) | ( ~n213 & n293 ) | ( n272 & n293 ) ;
  assign n295 = ( ~n110 & n213 ) | ( ~n110 & n294 ) | ( n213 & n294 ) ;
  assign n296 = ( ~n125 & n230 ) | ( ~n125 & n291 ) | ( n230 & n291 ) ;
  assign n297 = n273 | n281 ;
  assign n298 = n110 | n295 ;
  assign n299 = n104 & n105 ;
  assign n300 = n91 & ~n99 ;
  assign n301 = n89 & n161 ;
  assign n302 = n270 | n301 ;
  assign n303 = n107 & n158 ;
  assign n304 = n299 | n303 ;
  assign n305 = n300 ^ n190 ^ n179 ;
  assign n306 = n302 | n304 ;
  assign n307 = n94 & n112 ;
  assign n308 = ( n230 & n296 ) | ( n230 & ~n307 ) | ( n296 & ~n307 ) ;
  assign n309 = n107 & n130 ;
  assign n310 = n125 | n309 ;
  assign n311 = n91 & n161 ;
  assign n312 = n103 & n161 ;
  assign n313 = n306 | n310 ;
  assign n314 = n115 | n271 ;
  assign n315 = n266 | n312 ;
  assign n316 = n274 | n315 ;
  assign n317 = ( n283 & n313 ) | ( n283 & ~n316 ) | ( n313 & ~n316 ) ;
  assign n318 = n316 | n317 ;
  assign n319 = ( n180 & ~n229 ) | ( n180 & n311 ) | ( ~n229 & n311 ) ;
  assign n320 = n94 & n103 ;
  assign n321 = ( ~n177 & n254 ) | ( ~n177 & n318 ) | ( n254 & n318 ) ;
  assign n322 = ( n177 & ~n320 ) | ( n177 & n321 ) | ( ~n320 & n321 ) ;
  assign n323 = n305 | n314 ;
  assign n324 = n94 & n107 ;
  assign n325 = n89 & ~n99 ;
  assign n326 = n229 | n319 ;
  assign n327 = ~n230 & n308 ;
  assign n328 = n300 | n324 ;
  assign n329 = n170 | n315 ;
  assign n330 = ( ~n264 & n290 ) | ( ~n264 & n329 ) | ( n290 & n329 ) ;
  assign n331 = n320 | n322 ;
  assign n332 = n264 | n330 ;
  assign n333 = ( n176 & ~n305 ) | ( n176 & n327 ) | ( ~n305 & n327 ) ;
  assign n334 = ~n176 & n333 ;
  assign n335 = n91 & n130 ;
  assign n336 = n213 | n335 ;
  assign n337 = n331 | n336 ;
  assign n338 = ( n166 & ~n233 ) | ( n166 & n337 ) | ( ~n233 & n337 ) ;
  assign n339 = ( ~n237 & n258 ) | ( ~n237 & n328 ) | ( n258 & n328 ) ;
  assign n340 = n233 | n338 ;
  assign n341 = n237 | n339 ;
  assign n342 = ( n251 & ~n326 ) | ( n251 & n340 ) | ( ~n326 & n340 ) ;
  assign n343 = n78 & n158 ;
  assign n344 = ( ~n136 & n332 ) | ( ~n136 & n343 ) | ( n332 & n343 ) ;
  assign n345 = ( ~n136 & n324 ) | ( ~n136 & n344 ) | ( n324 & n344 ) ;
  assign n346 = n326 | n342 ;
  assign n347 = n136 | n345 ;
  assign n348 = n91 & n158 ;
  assign n349 = n107 & n161 ;
  assign n350 = ( n114 & ~n311 ) | ( n114 & n341 ) | ( ~n311 & n341 ) ;
  assign n351 = n311 | n350 ;
  assign n352 = n112 & n120 ;
  assign n353 = ~n106 & n158 ;
  assign n354 = n163 | n352 ;
  assign n355 = n94 | n158 ;
  assign n356 = n121 & n130 ;
  assign n357 = n103 & n130 ;
  assign n358 = n348 | n357 ;
  assign n359 = n90 & n94 ;
  assign n360 = n78 & n130 ;
  assign n361 = ( n116 & n355 ) | ( n116 & n359 ) | ( n355 & n359 ) ;
  assign n362 = n182 | n302 ;
  assign n363 = n262 | n360 ;
  assign n364 = ( ~n141 & n354 ) | ( ~n141 & n356 ) | ( n354 & n356 ) ;
  assign n365 = n141 | n364 ;
  assign n366 = n116 & n161 ;
  assign n367 = ( ~n147 & n353 ) | ( ~n147 & n365 ) | ( n353 & n365 ) ;
  assign n368 = n147 | n367 ;
  assign n369 = n74 & n158 ;
  assign n370 = n349 | n361 ;
  assign n371 = n227 | n366 ;
  assign n372 = ( n325 & n368 ) | ( n325 & ~n369 ) | ( n368 & ~n369 ) ;
  assign n373 = n369 | n372 ;
  assign n374 = ( n265 & ~n370 ) | ( n265 & n373 ) | ( ~n370 & n373 ) ;
  assign n375 = ( n253 & n371 ) | ( n253 & ~n373 ) | ( n371 & ~n373 ) ;
  assign n376 = n373 | n375 ;
  assign n377 = n370 | n374 ;
  assign n378 = n110 | n307 ;
  assign n379 = ( ~n177 & n353 ) | ( ~n177 & n358 ) | ( n353 & n358 ) ;
  assign n380 = n177 | n379 ;
  assign n381 = ( ~n315 & n378 ) | ( ~n315 & n380 ) | ( n378 & n380 ) ;
  assign n382 = ( ~n362 & n363 ) | ( ~n362 & n371 ) | ( n363 & n371 ) ;
  assign n383 = n224 | n264 ;
  assign n384 = n315 | n381 ;
  assign n385 = n362 | n382 ;
  assign n386 = ( n129 & ~n378 ) | ( n129 & n385 ) | ( ~n378 & n385 ) ;
  assign n387 = ~n385 & n386 ;
  assign n388 = n383 | n385 ;
  assign n389 = ~n99 & n103 ;
  assign n390 = ( n258 & n384 ) | ( n258 & ~n389 ) | ( n384 & ~n389 ) ;
  assign n391 = n389 | n390 ;
  assign n392 = n78 & n94 ;
  assign n393 = n94 & n104 ;
  assign n394 = n90 & ~n99 ;
  assign n395 = n112 & n158 ;
  assign n396 = n104 & n161 ;
  assign n397 = n121 & n158 ;
  assign n398 = n256 | n311 ;
  assign n399 = n105 & n116 ;
  assign n400 = n181 | n221 ;
  assign n401 = n178 | n309 ;
  assign n402 = ( ~n398 & n400 ) | ( ~n398 & n401 ) | ( n400 & n401 ) ;
  assign n403 = n398 | n402 ;
  assign n404 = n78 & n120 ;
  assign n405 = n104 | n112 ;
  assign n406 = ( n94 & n352 ) | ( n94 & n405 ) | ( n352 & n405 ) ;
  assign n407 = n224 | n397 ;
  assign n408 = n104 & n158 ;
  assign n409 = ( n143 & n273 ) | ( n143 & ~n407 ) | ( n273 & ~n407 ) ;
  assign n410 = n407 | n409 ;
  assign n411 = n116 & n158 ;
  assign n412 = n357 | n399 ;
  assign n413 = n404 | n412 ;
  assign n414 = ( ~n403 & n410 ) | ( ~n403 & n413 ) | ( n410 & n413 ) ;
  assign n415 = n403 | n414 ;
  assign n416 = n94 & n121 ;
  assign n417 = ( n94 & n116 ) | ( n94 & n416 ) | ( n116 & n416 ) ;
  assign n418 = ( n256 & ~n272 ) | ( n256 & n408 ) | ( ~n272 & n408 ) ;
  assign n419 = n94 & n116 ;
  assign n420 = ( n234 & ~n264 ) | ( n234 & n415 ) | ( ~n264 & n415 ) ;
  assign n421 = n264 | n420 ;
  assign n422 = ( ~n394 & n411 ) | ( ~n394 & n421 ) | ( n411 & n421 ) ;
  assign n423 = n394 | n422 ;
  assign n424 = ( n156 & n387 ) | ( n156 & ~n423 ) | ( n387 & ~n423 ) ;
  assign n425 = ~n156 & n424 ;
  assign n426 = n74 & n94 ;
  assign n427 = ( ~n163 & n396 ) | ( ~n163 & n425 ) | ( n396 & n425 ) ;
  assign n428 = n74 & ~n99 ;
  assign n429 = ~n396 & n427 ;
  assign n430 = ( n395 & ~n408 ) | ( n395 & n429 ) | ( ~n408 & n429 ) ;
  assign n431 = ~n395 & n430 ;
  assign n432 = n272 | n418 ;
  assign n433 = ~n99 & n112 ;
  assign n434 = ( n238 & n431 ) | ( n238 & ~n433 ) | ( n431 & ~n433 ) ;
  assign n435 = ( n238 & ~n393 ) | ( n238 & n434 ) | ( ~n393 & n434 ) ;
  assign n436 = ~n238 & n435 ;
  assign n437 = n224 | n404 ;
  assign n438 = n95 & n161 ;
  assign n439 = n335 | n438 ;
  assign n440 = n320 | n348 ;
  assign n441 = n90 & n98 ;
  assign n442 = n299 | n439 ;
  assign n443 = ( ~n122 & n437 ) | ( ~n122 & n442 ) | ( n437 & n442 ) ;
  assign n444 = n122 | n443 ;
  assign n445 = ( ~n389 & n397 ) | ( ~n389 & n441 ) | ( n397 & n441 ) ;
  assign n446 = n213 | n411 ;
  assign n447 = n105 & ~n106 ;
  assign n448 = n225 | n406 ;
  assign n449 = n389 | n445 ;
  assign n450 = n98 & ~n106 ;
  assign n451 = n366 | n440 ;
  assign n452 = ( n444 & ~n448 ) | ( n444 & n451 ) | ( ~n448 & n451 ) ;
  assign n453 = n448 | n452 ;
  assign n454 = ( n255 & ~n272 ) | ( n255 & n453 ) | ( ~n272 & n453 ) ;
  assign n455 = n272 | n454 ;
  assign n456 = ( n133 & ~n428 ) | ( n133 & n455 ) | ( ~n428 & n455 ) ;
  assign n457 = n428 | n456 ;
  assign n458 = n126 | n457 ;
  assign n459 = n98 & n103 ;
  assign n460 = n95 & n105 ;
  assign n461 = ( n210 & ~n310 ) | ( n210 & n458 ) | ( ~n310 & n458 ) ;
  assign n462 = n416 | n439 ;
  assign n463 = n310 | n461 ;
  assign n464 = ( ~n351 & n449 ) | ( ~n351 & n463 ) | ( n449 & n463 ) ;
  assign n465 = n351 | n464 ;
  assign n466 = ( n437 & n446 ) | ( n437 & ~n460 ) | ( n446 & ~n460 ) ;
  assign n467 = ( ~n231 & n396 ) | ( ~n231 & n459 ) | ( n396 & n459 ) ;
  assign n468 = n231 | n467 ;
  assign n469 = ( ~n270 & n465 ) | ( ~n270 & n468 ) | ( n465 & n468 ) ;
  assign n470 = n270 | n469 ;
  assign n471 = ( n356 & ~n357 ) | ( n356 & n470 ) | ( ~n357 & n470 ) ;
  assign n472 = n357 | n471 ;
  assign n473 = ( ~n139 & n227 ) | ( ~n139 & n472 ) | ( n227 & n472 ) ;
  assign n474 = n139 | n473 ;
  assign n475 = ( n408 & ~n450 ) | ( n408 & n474 ) | ( ~n450 & n474 ) ;
  assign n476 = n103 & n158 ;
  assign n477 = n250 | n457 ;
  assign n478 = n95 & n158 ;
  assign n479 = ( n416 & ~n450 ) | ( n416 & n475 ) | ( ~n450 & n475 ) ;
  assign n480 = n450 | n479 ;
  assign n481 = n90 & n105 ;
  assign n482 = n95 & n120 ;
  assign n483 = n459 | n482 ;
  assign n484 = n423 | n483 ;
  assign n485 = n216 | n312 ;
  assign n486 = n148 | n460 ;
  assign n487 = n303 | n438 ;
  assign n488 = n90 & n130 ;
  assign n489 = n227 | n481 ;
  assign n490 = ( n369 & ~n426 ) | ( n369 & n489 ) | ( ~n426 & n489 ) ;
  assign n491 = n183 | n488 ;
  assign n492 = n426 | n490 ;
  assign n493 = n324 | n491 ;
  assign n494 = ( n485 & ~n486 ) | ( n485 & n492 ) | ( ~n486 & n492 ) ;
  assign n495 = n486 | n494 ;
  assign n496 = ( ~n136 & n299 ) | ( ~n136 & n495 ) | ( n299 & n495 ) ;
  assign n497 = n136 | n496 ;
  assign n498 = ( n484 & n493 ) | ( n484 & ~n497 ) | ( n493 & ~n497 ) ;
  assign n499 = n497 | n498 ;
  assign n500 = ( ~n286 & n487 ) | ( ~n286 & n499 ) | ( n487 & n499 ) ;
  assign n501 = n286 | n500 ;
  assign n502 = n95 & n130 ;
  assign n503 = n290 | n359 ;
  assign n504 = ( n399 & ~n502 ) | ( n399 & n503 ) | ( ~n502 & n503 ) ;
  assign n505 = ( n90 & n120 ) | ( n90 & n217 ) | ( n120 & n217 ) ;
  assign n506 = n502 | n504 ;
  assign n507 = ( ~n203 & n325 ) | ( ~n203 & n506 ) | ( n325 & n506 ) ;
  assign n508 = n203 | n507 ;
  assign n509 = ( ~n136 & n302 ) | ( ~n136 & n508 ) | ( n302 & n508 ) ;
  assign n510 = ( n250 & ~n323 ) | ( n250 & n501 ) | ( ~n323 & n501 ) ;
  assign n511 = n96 & n161 ;
  assign n512 = n96 & n130 ;
  assign n513 = n112 & n130 ;
  assign n514 = n112 & n161 ;
  assign n515 = n323 | n510 ;
  assign n516 = n163 | n397 ;
  assign n517 = ( ~n141 & n512 ) | ( ~n141 & n515 ) | ( n512 & n515 ) ;
  assign n518 = n141 | n517 ;
  assign n519 = ( ~n175 & n220 ) | ( ~n175 & n518 ) | ( n220 & n518 ) ;
  assign n520 = n175 | n519 ;
  assign n521 = ( ~n101 & n238 ) | ( ~n101 & n520 ) | ( n238 & n520 ) ;
  assign n522 = ( n189 & ~n349 ) | ( n189 & n516 ) | ( ~n349 & n516 ) ;
  assign n523 = n460 | n466 ;
  assign n524 = n136 | n509 ;
  assign n525 = ( n196 & ~n483 ) | ( n196 & n524 ) | ( ~n483 & n524 ) ;
  assign n526 = n483 | n525 ;
  assign n527 = ( ~n125 & n496 ) | ( ~n125 & n526 ) | ( n496 & n526 ) ;
  assign n528 = n115 | n478 ;
  assign n529 = n302 | n528 ;
  assign n530 = n101 | n521 ;
  assign n531 = n125 | n527 ;
  assign n532 = n349 | n522 ;
  assign n533 = n266 | n478 ;
  assign n534 = n146 | n233 ;
  assign n535 = n369 | n502 ;
  assign n536 = n139 | n264 ;
  assign n537 = n159 | n231 ;
  assign n538 = n276 | n353 ;
  assign n539 = n115 | n212 ;
  assign n540 = n173 | n391 ;
  assign n541 = n126 | n273 ;
  assign n542 = n534 | n539 ;
  assign n543 = ( n533 & ~n538 ) | ( n533 & n542 ) | ( ~n538 & n542 ) ;
  assign n544 = n234 | n396 ;
  assign n545 = n535 | n544 ;
  assign n546 = ( n534 & n536 ) | ( n534 & ~n545 ) | ( n536 & ~n545 ) ;
  assign n547 = n538 | n543 ;
  assign n548 = ( n351 & ~n537 ) | ( n351 & n547 ) | ( ~n537 & n547 ) ;
  assign n549 = n159 | n174 ;
  assign n550 = ( ~n447 & n544 ) | ( ~n447 & n549 ) | ( n544 & n549 ) ;
  assign n551 = ( ~n540 & n541 ) | ( ~n540 & n545 ) | ( n541 & n545 ) ;
  assign n552 = n540 | n551 ;
  assign n553 = n537 | n548 ;
  assign n554 = n512 | n513 ;
  assign n555 = n366 | n514 ;
  assign n556 = n545 | n546 ;
  assign n557 = ( n101 & ~n110 ) | ( n101 & n553 ) | ( ~n110 & n553 ) ;
  assign n558 = n110 | n557 ;
  assign n559 = ( ~n477 & n508 ) | ( ~n477 & n558 ) | ( n508 & n558 ) ;
  assign n560 = n324 | n447 ;
  assign n561 = n477 | n559 ;
  assign n562 = ( ~n171 & n554 ) | ( ~n171 & n560 ) | ( n554 & n560 ) ;
  assign n563 = n447 | n550 ;
  assign n564 = n171 | n562 ;
  assign n565 = n147 | n555 ;
  assign n566 = n401 | n555 ;
  assign n567 = ( n529 & n564 ) | ( n529 & ~n566 ) | ( n564 & ~n566 ) ;
  assign n568 = n566 | n567 ;
  assign n569 = n300 | n488 ;
  assign n570 = ( ~n271 & n349 ) | ( ~n271 & n568 ) | ( n349 & n568 ) ;
  assign n571 = n271 | n570 ;
  assign n572 = ( ~n137 & n460 ) | ( ~n137 & n571 ) | ( n460 & n571 ) ;
  assign n573 = n137 | n572 ;
  assign n574 = n569 | n573 ;
  assign n575 = ( n326 & n552 ) | ( n326 & ~n574 ) | ( n552 & ~n574 ) ;
  assign n576 = n574 | n575 ;
  assign n577 = ( n433 & ~n450 ) | ( n433 & n576 ) | ( ~n450 & n576 ) ;
  assign n578 = n450 | n577 ;
  assign n579 = n196 | n574 ;
  assign n580 = n101 | n389 ;
  assign n581 = n122 | n237 ;
  assign n582 = n511 ^ n441 ^ n143 ;
  assign n583 = n218 | n582 ;
  assign n584 = n324 | n411 ;
  assign n585 = n135 | n393 ;
  assign n586 = n187 | n581 ;
  assign n587 = ( ~n583 & n584 ) | ( ~n583 & n585 ) | ( n584 & n585 ) ;
  assign n588 = n583 | n587 ;
  assign n589 = n538 | n580 ;
  assign n590 = ( n432 & ~n586 ) | ( n432 & n589 ) | ( ~n586 & n589 ) ;
  assign n591 = ( n192 & n432 ) | ( n192 & ~n588 ) | ( n432 & ~n588 ) ;
  assign n592 = n588 | n591 ;
  assign n593 = ( n168 & ~n324 ) | ( n168 & n395 ) | ( ~n324 & n395 ) ;
  assign n594 = n324 | n593 ;
  assign n595 = ( ~n132 & n182 ) | ( ~n132 & n563 ) | ( n182 & n563 ) ;
  assign n596 = n132 | n595 ;
  assign n597 = ( ~n132 & n323 ) | ( ~n132 & n592 ) | ( n323 & n592 ) ;
  assign n598 = n132 | n597 ;
  assign n599 = ( ~n262 & n488 ) | ( ~n262 & n598 ) | ( n488 & n598 ) ;
  assign n600 = ( n331 & ~n554 ) | ( n331 & n596 ) | ( ~n554 & n596 ) ;
  assign n601 = n554 | n600 ;
  assign n602 = ( n212 & ~n262 ) | ( n212 & n601 ) | ( ~n262 & n601 ) ;
  assign n603 = ( n231 & ~n262 ) | ( n231 & n599 ) | ( ~n262 & n599 ) ;
  assign n604 = n262 | n603 ;
  assign n605 = n586 | n590 ;
  assign n606 = n262 | n602 ;
  assign n607 = n482 | n582 ;
  assign n608 = ( n220 & ~n450 ) | ( n220 & n606 ) | ( ~n450 & n606 ) ;
  assign n609 = ( ~n137 & n325 ) | ( ~n137 & n607 ) | ( n325 & n607 ) ;
  assign n610 = n137 | n609 ;
  assign n611 = ( ~n532 & n563 ) | ( ~n532 & n605 ) | ( n563 & n605 ) ;
  assign n612 = ( ~n401 & n541 ) | ( ~n401 & n594 ) | ( n541 & n594 ) ;
  assign n613 = n401 | n612 ;
  assign n614 = n450 | n608 ;
  assign n615 = n532 | n611 ;
  assign n616 = ( ~n125 & n440 ) | ( ~n125 & n615 ) | ( n440 & n615 ) ;
  assign n617 = ( ~n233 & n531 ) | ( ~n233 & n616 ) | ( n531 & n616 ) ;
  assign n618 = ( ~n233 & n252 ) | ( ~n233 & n617 ) | ( n252 & n617 ) ;
  assign n619 = n233 | n618 ;
  assign n620 = ( n192 & ~n511 ) | ( n192 & n619 ) | ( ~n511 & n619 ) ;
  assign n621 = ( n124 & n487 ) | ( n124 & ~n613 ) | ( n487 & ~n613 ) ;
  assign n622 = n511 | n620 ;
  assign n623 = ( n335 & ~n352 ) | ( n335 & n622 ) | ( ~n352 & n622 ) ;
  assign n624 = n613 | n621 ;
  assign n625 = n164 | n343 ;
  assign n626 = n594 | n625 ;
  assign n627 = ( n346 & n532 ) | ( n346 & ~n626 ) | ( n532 & ~n626 ) ;
  assign n628 = n125 | n616 ;
  assign n629 = n352 | n623 ;
  assign n630 = ( ~n394 & n478 ) | ( ~n394 & n629 ) | ( n478 & n629 ) ;
  assign n631 = ( ~n307 & n394 ) | ( ~n307 & n630 ) | ( n394 & n630 ) ;
  assign n632 = n307 | n631 ;
  assign n633 = n626 | n627 ;
  assign n634 = n235 | n360 ;
  assign n635 = n217 ^ n177 ^ n163 ;
  assign n636 = n175 | n634 ;
  assign n637 = n182 | n404 ;
  assign n638 = ( n86 & n511 ) | ( n86 & n636 ) | ( n511 & n636 ) ;
  assign n639 = ( n635 & n637 ) | ( n635 & ~n638 ) | ( n637 & ~n638 ) ;
  assign n640 = n638 | n639 ;
  assign n641 = n356 ^ n222 ^ n220 ;
  assign n642 = n139 | n235 ;
  assign n643 = ( ~n492 & n640 ) | ( ~n492 & n641 ) | ( n640 & n641 ) ;
  assign n644 = n132 | n290 ;
  assign n645 = ( ~n565 & n635 ) | ( ~n565 & n642 ) | ( n635 & n642 ) ;
  assign n646 = n492 | n643 ;
  assign n647 = n565 | n645 ;
  assign n648 = ( n254 & ~n264 ) | ( n254 & n646 ) | ( ~n264 & n646 ) ;
  assign n649 = n512 ^ n459 ^ n349 ;
  assign n650 = n235 | n585 ;
  assign n651 = n238 | n304 ;
  assign n652 = n274 | n649 ;
  assign n653 = ( n149 & n650 ) | ( n149 & ~n651 ) | ( n650 & ~n651 ) ;
  assign n654 = n651 | n653 ;
  assign n655 = ( ~n560 & n641 ) | ( ~n560 & n652 ) | ( n641 & n652 ) ;
  assign n656 = n180 | n399 ;
  assign n657 = n644 | n656 ;
  assign n658 = ( n505 & n649 ) | ( n505 & ~n657 ) | ( n649 & ~n657 ) ;
  assign n659 = n264 | n648 ;
  assign n660 = n560 | n655 ;
  assign n661 = ( ~n110 & n399 ) | ( ~n110 & n659 ) | ( n399 & n659 ) ;
  assign n662 = n132 | n394 ;
  assign n663 = ( ~n396 & n580 ) | ( ~n396 & n662 ) | ( n580 & n662 ) ;
  assign n664 = n129 & ~n656 ;
  assign n665 = n537 | n654 ;
  assign n666 = ( ~n580 & n664 ) | ( ~n580 & n665 ) | ( n664 & n665 ) ;
  assign n667 = n141 | n146 ;
  assign n668 = ( n267 & n579 ) | ( n267 & ~n667 ) | ( n579 & ~n667 ) ;
  assign n669 = n667 | n668 ;
  assign n670 = n394 | n636 ;
  assign n671 = n110 | n661 ;
  assign n672 = n396 | n663 ;
  assign n673 = ~n665 & n666 ;
  assign n674 = ( n665 & n669 ) | ( n665 & ~n671 ) | ( n669 & ~n671 ) ;
  assign n675 = n189 | n395 ;
  assign n676 = n657 | n658 ;
  assign n677 = n179 | n211 ;
  assign n678 = n671 | n674 ;
  assign n679 = n417 | n677 ;
  assign n680 = ( n353 & n678 ) | ( n353 & ~n679 ) | ( n678 & ~n679 ) ;
  assign n681 = n679 | n680 ;
  assign n682 = ( ~n160 & n675 ) | ( ~n160 & n681 ) | ( n675 & n681 ) ;
  assign n683 = ( n160 & ~n284 ) | ( n160 & n682 ) | ( ~n284 & n682 ) ;
  assign n684 = n284 | n683 ;
  assign n685 = n349 | n644 ;
  assign n686 = ( ~n462 & n626 ) | ( ~n462 & n685 ) | ( n626 & n685 ) ;
  assign n687 = n462 | n686 ;
  assign n688 = n271 | n441 ;
  assign n689 = n254 | n670 ;
  assign n690 = n644 | n667 ;
  assign n691 = n264 | n348 ;
  assign n692 = n528 | n670 ;
  assign n693 = n188 | n312 ;
  assign n694 = n656 | n693 ;
  assign n695 = n357 | n488 ;
  assign n696 = ( ~n147 & n323 ) | ( ~n147 & n689 ) | ( n323 & n689 ) ;
  assign n697 = n298 | n502 ;
  assign n698 = n426 | n433 ;
  assign n699 = n135 | n148 ;
  assign n700 = n667 | n699 ;
  assign n701 = n298 | n528 ;
  assign n702 = n400 | n462 ;
  assign n703 = ( ~n695 & n698 ) | ( ~n695 & n700 ) | ( n698 & n700 ) ;
  assign n704 = n695 | n703 ;
  assign n705 = ( ~n688 & n692 ) | ( ~n688 & n704 ) | ( n692 & n704 ) ;
  assign n706 = n688 | n705 ;
  assign n707 = ( ~n136 & n237 ) | ( ~n136 & n706 ) | ( n237 & n706 ) ;
  assign n708 = n136 | n707 ;
  assign n709 = ( ~n359 & n428 ) | ( ~n359 & n708 ) | ( n428 & n708 ) ;
  assign n710 = ( n307 & ~n359 ) | ( n307 & n709 ) | ( ~n359 & n709 ) ;
  assign n711 = n359 | n710 ;
  assign n712 = ( n356 & n633 ) | ( n356 & ~n711 ) | ( n633 & ~n711 ) ;
  assign n713 = n711 | n712 ;
  assign n714 = ( ~n139 & n459 ) | ( ~n139 & n713 ) | ( n459 & n713 ) ;
  assign n715 = n301 | n481 ;
  assign n716 = n139 | n714 ;
  assign n717 = ( n101 & ~n460 ) | ( n101 & n716 ) | ( ~n460 & n716 ) ;
  assign n718 = ( n679 & ~n691 ) | ( n679 & n711 ) | ( ~n691 & n711 ) ;
  assign n719 = n691 | n718 ;
  assign n720 = n229 | n514 ;
  assign n721 = n139 | n389 ;
  assign n722 = ( n693 & n715 ) | ( n693 & ~n721 ) | ( n715 & ~n721 ) ;
  assign n723 = n721 | n722 ;
  assign n724 = n720 | n723 ;
  assign n725 = ( n697 & n719 ) | ( n697 & ~n724 ) | ( n719 & ~n724 ) ;
  assign n726 = n724 | n725 ;
  assign n727 = ( n300 & ~n309 ) | ( n300 & n513 ) | ( ~n309 & n513 ) ;
  assign n728 = n309 | n727 ;
  assign n729 = ( ~n138 & n482 ) | ( ~n138 & n726 ) | ( n482 & n726 ) ;
  assign n730 = ( n687 & ~n704 ) | ( n687 & n728 ) | ( ~n704 & n728 ) ;
  assign n731 = ( ~n310 & n487 ) | ( ~n310 & n694 ) | ( n487 & n694 ) ;
  assign n732 = n310 | n731 ;
  assign n733 = n704 | n730 ;
  assign n734 = n108 & ~n146 ;
  assign n735 = ~n693 & n734 ;
  assign n736 = ( n189 & ~n270 ) | ( n189 & n733 ) | ( ~n270 & n733 ) ;
  assign n737 = ( n554 & ~n698 ) | ( n554 & n735 ) | ( ~n698 & n735 ) ;
  assign n738 = n147 | n696 ;
  assign n739 = n138 | n729 ;
  assign n740 = ( n303 & ~n450 ) | ( n303 & n739 ) | ( ~n450 & n739 ) ;
  assign n741 = n450 | n740 ;
  assign n742 = n270 | n736 ;
  assign n743 = ( ~n181 & n369 ) | ( ~n181 & n742 ) | ( n369 & n742 ) ;
  assign n744 = n460 | n717 ;
  assign n745 = n181 | n743 ;
  assign n746 = ( ~n159 & n187 ) | ( ~n159 & n741 ) | ( n187 & n741 ) ;
  assign n747 = ( n137 & ~n399 ) | ( n137 & n745 ) | ( ~n399 & n745 ) ;
  assign n748 = n167 | n746 ;
  assign n749 = ~n554 & n737 ;
  assign n750 = n132 | n359 ;
  assign n751 = n211 | n450 ;
  assign n752 = n135 | n141 ;
  assign n753 = n138 | n441 ;
  assign n754 = n178 | n419 ;
  assign n755 = n180 | n369 ;
  assign n756 = ( n184 & n320 ) | ( n184 & ~n750 ) | ( n320 & ~n750 ) ;
  assign n757 = n750 | n756 ;
  assign n758 = n133 | n261 ;
  assign n759 = n751 | n758 ;
  assign n760 = ( ~n101 & n274 ) | ( ~n101 & n759 ) | ( n274 & n759 ) ;
  assign n761 = n101 | n760 ;
  assign n762 = n220 | n476 ;
  assign n763 = ( n218 & ~n476 ) | ( n218 & n752 ) | ( ~n476 & n752 ) ;
  assign n764 = ( n137 & ~n755 ) | ( n137 & n762 ) | ( ~n755 & n762 ) ;
  assign n765 = ( n638 & ~n753 ) | ( n638 & n757 ) | ( ~n753 & n757 ) ;
  assign n766 = n755 | n764 ;
  assign n767 = n476 | n763 ;
  assign n768 = n366 | n482 ;
  assign n769 = n754 | n761 ;
  assign n770 = ( n449 & n768 ) | ( n449 & ~n769 ) | ( n768 & ~n769 ) ;
  assign n771 = n769 | n770 ;
  assign n772 = n126 | n416 ;
  assign n773 = n266 | n482 ;
  assign n774 = ( ~n406 & n766 ) | ( ~n406 & n773 ) | ( n766 & n773 ) ;
  assign n775 = ( ~n392 & n406 ) | ( ~n392 & n774 ) | ( n406 & n774 ) ;
  assign n776 = n586 | n772 ;
  assign n777 = ( ~n122 & n143 ) | ( ~n122 & n771 ) | ( n143 & n771 ) ;
  assign n778 = n392 | n775 ;
  assign n779 = ( n423 & ~n776 ) | ( n423 & n778 ) | ( ~n776 & n778 ) ;
  assign n780 = n776 | n779 ;
  assign n781 = n753 | n765 ;
  assign n782 = n122 | n777 ;
  assign n783 = ( n114 & ~n173 ) | ( n114 & n782 ) | ( ~n173 & n782 ) ;
  assign n784 = n173 | n783 ;
  assign n785 = n143 | n352 ;
  assign n786 = ( n647 & ~n780 ) | ( n647 & n781 ) | ( ~n780 & n781 ) ;
  assign n787 = n780 | n786 ;
  assign n788 = n216 | n502 ;
  assign n789 = ( n173 & ~n585 ) | ( n173 & n788 ) | ( ~n585 & n788 ) ;
  assign n790 = n585 | n789 ;
  assign n791 = ( n354 & ~n762 ) | ( n354 & n790 ) | ( ~n762 & n790 ) ;
  assign n792 = ( ~n216 & n304 ) | ( ~n216 & n787 ) | ( n304 & n787 ) ;
  assign n793 = ( ~n148 & n182 ) | ( ~n148 & n781 ) | ( n182 & n781 ) ;
  assign n794 = n762 | n791 ;
  assign n795 = n148 | n793 ;
  assign n796 = n354 | n795 ;
  assign n797 = n301 | n762 ;
  assign n798 = n216 | n792 ;
  assign n799 = ( ~n133 & n491 ) | ( ~n133 & n798 ) | ( n491 & n798 ) ;
  assign n800 = n114 | n356 ;
  assign n801 = ( ~n189 & n767 ) | ( ~n189 & n800 ) | ( n767 & n800 ) ;
  assign n802 = n189 | n801 ;
  assign n803 = ( n702 & ~n796 ) | ( n702 & n802 ) | ( ~n796 & n802 ) ;
  assign n804 = n796 | n803 ;
  assign n805 = n232 | n393 ;
  assign n806 = ( n263 & ~n578 ) | ( n263 & n805 ) | ( ~n578 & n805 ) ;
  assign n807 = ( ~n393 & n578 ) | ( ~n393 & n804 ) | ( n578 & n804 ) ;
  assign n808 = n578 | n806 ;
  assign n809 = n229 | n404 ;
  assign n810 = ( ~n230 & n232 ) | ( ~n230 & n809 ) | ( n232 & n809 ) ;
  assign n811 = n230 | n810 ;
  assign n812 = n676 | n811 ;
  assign n813 = ( n761 & n797 ) | ( n761 & ~n812 ) | ( n797 & ~n812 ) ;
  assign n814 = n812 | n813 ;
  assign n815 = n238 | n255 ;
  assign n816 = n110 | n394 ;
  assign n817 = ( ~n139 & n360 ) | ( ~n139 & n488 ) | ( n360 & n488 ) ;
  assign n818 = ( n189 & ~n227 ) | ( n189 & n814 ) | ( ~n227 & n814 ) ;
  assign n819 = ( n538 & ~n560 ) | ( n538 & n816 ) | ( ~n560 & n816 ) ;
  assign n820 = n560 | n819 ;
  assign n821 = ( ~n159 & n348 ) | ( ~n159 & n794 ) | ( n348 & n794 ) ;
  assign n822 = n117 | n180 ;
  assign n823 = n216 | n357 ;
  assign n824 = ( ~n538 & n701 ) | ( ~n538 & n815 ) | ( n701 & n815 ) ;
  assign n825 = n538 | n824 ;
  assign n826 = ( n290 & ~n428 ) | ( n290 & n476 ) | ( ~n428 & n476 ) ;
  assign n827 = n139 | n817 ;
  assign n828 = n227 | n818 ;
  assign n829 = ( n438 & ~n514 ) | ( n438 & n823 ) | ( ~n514 & n823 ) ;
  assign n830 = ( n468 & ~n795 ) | ( n468 & n825 ) | ( ~n795 & n825 ) ;
  assign n831 = n514 | n829 ;
  assign n832 = ( n751 & n822 ) | ( n751 & ~n831 ) | ( n822 & ~n831 ) ;
  assign n833 = n795 | n830 ;
  assign n834 = n831 | n832 ;
  assign n835 = ( n135 & ~n138 ) | ( n135 & n262 ) | ( ~n138 & n262 ) ;
  assign n836 = ( ~n159 & n261 ) | ( ~n159 & n821 ) | ( n261 & n821 ) ;
  assign n837 = n159 | n836 ;
  assign n838 = ( ~n772 & n785 ) | ( ~n772 & n820 ) | ( n785 & n820 ) ;
  assign n839 = n772 | n838 ;
  assign n840 = n428 | n826 ;
  assign n841 = ( ~n827 & n834 ) | ( ~n827 & n840 ) | ( n834 & n840 ) ;
  assign n842 = ( n310 & ~n772 ) | ( n310 & n840 ) | ( ~n772 & n840 ) ;
  assign n843 = n772 | n842 ;
  assign n844 = ( ~n138 & n399 ) | ( ~n138 & n747 ) | ( n399 & n747 ) ;
  assign n845 = n138 | n835 ;
  assign n846 = n138 | n844 ;
  assign n847 = n138 | n203 ;
  assign n848 = ( n101 & ~n299 ) | ( n101 & n847 ) | ( ~n299 & n847 ) ;
  assign n849 = ( ~n311 & n511 ) | ( ~n311 & n846 ) | ( n511 & n846 ) ;
  assign n850 = n827 | n841 ;
  assign n851 = ( n221 & ~n359 ) | ( n221 & n839 ) | ( ~n359 & n839 ) ;
  assign n852 = n299 | n848 ;
  assign n853 = ( ~n220 & n751 ) | ( ~n220 & n852 ) | ( n751 & n852 ) ;
  assign n854 = n126 | n751 ;
  assign n855 = ( n210 & ~n815 ) | ( n210 & n854 ) | ( ~n815 & n854 ) ;
  assign n856 = n815 | n855 ;
  assign n857 = ( n377 & ~n672 ) | ( n377 & n827 ) | ( ~n672 & n827 ) ;
  assign n858 = n672 | n857 ;
  assign n859 = ( n122 & ~n136 ) | ( n122 & n858 ) | ( ~n136 & n858 ) ;
  assign n860 = ( ~n234 & n476 ) | ( ~n234 & n513 ) | ( n476 & n513 ) ;
  assign n861 = n136 | n859 ;
  assign n862 = n234 | n860 ;
  assign n863 = ( ~n313 & n856 ) | ( ~n313 & n862 ) | ( n856 & n862 ) ;
  assign n864 = n313 | n863 ;
  assign n865 = ( n561 & n845 ) | ( n561 & ~n862 ) | ( n845 & ~n862 ) ;
  assign n866 = ( ~n720 & n861 ) | ( ~n720 & n864 ) | ( n861 & n864 ) ;
  assign n867 = n141 | n273 ;
  assign n868 = ( n114 & ~n221 ) | ( n114 & n867 ) | ( ~n221 & n867 ) ;
  assign n869 = n221 | n868 ;
  assign n870 = n862 | n865 ;
  assign n871 = n146 | n290 ;
  assign n872 = ( n137 & ~n426 ) | ( n137 & n850 ) | ( ~n426 & n850 ) ;
  assign n873 = ( ~n404 & n459 ) | ( ~n404 & n871 ) | ( n459 & n871 ) ;
  assign n874 = n404 | n873 ;
  assign n875 = n310 | n404 ;
  assign n876 = n426 | n872 ;
  assign n877 = n233 | n310 ;
  assign n878 = ( n252 & ~n837 ) | ( n252 & n877 ) | ( ~n837 & n877 ) ;
  assign n879 = ( ~n378 & n869 ) | ( ~n378 & n876 ) | ( n869 & n876 ) ;
  assign n880 = n359 | n851 ;
  assign n881 = n378 | n879 ;
  assign n882 = ( ~n811 & n845 ) | ( ~n811 & n881 ) | ( n845 & n881 ) ;
  assign n883 = n311 | n849 ;
  assign n884 = n183 | n476 ;
  assign n885 = n811 | n882 ;
  assign n886 = ( ~n542 & n628 ) | ( ~n542 & n885 ) | ( n628 & n885 ) ;
  assign n887 = n542 | n886 ;
  assign n888 = ( n190 & ~n264 ) | ( n190 & n887 ) | ( ~n264 & n887 ) ;
  assign n889 = n264 | n888 ;
  assign n890 = ( n160 & ~n183 ) | ( n160 & n889 ) | ( ~n183 & n889 ) ;
  assign n891 = n220 | n853 ;
  assign n892 = n218 | n542 ;
  assign n893 = ( n183 & ~n433 ) | ( n183 & n890 ) | ( ~n433 & n890 ) ;
  assign n894 = n134 | n227 ;
  assign n895 = n558 | n894 ;
  assign n896 = n233 | n254 ;
  assign n897 = ( n190 & ~n352 ) | ( n190 & n896 ) | ( ~n352 & n896 ) ;
  assign n898 = n352 | n897 ;
  assign n899 = ( ~n304 & n876 ) | ( ~n304 & n895 ) | ( n876 & n895 ) ;
  assign n900 = n304 | n899 ;
  assign n901 = n224 | n234 ;
  assign n902 = ( n348 & n447 ) | ( n348 & ~n481 ) | ( n447 & ~n481 ) ;
  assign n903 = ( ~n126 & n898 ) | ( ~n126 & n901 ) | ( n898 & n901 ) ;
  assign n904 = n337 | n894 ;
  assign n905 = n481 | n902 ;
  assign n906 = ( ~n410 & n904 ) | ( ~n410 & n905 ) | ( n904 & n905 ) ;
  assign n907 = n126 | n903 ;
  assign n908 = n410 | n906 ;
  assign n909 = ( n634 & ~n698 ) | ( n634 & n907 ) | ( ~n698 & n907 ) ;
  assign n910 = n698 | n909 ;
  assign n911 = ( n315 & ~n400 ) | ( n315 & n910 ) | ( ~n400 & n910 ) ;
  assign n912 = n400 | n911 ;
  assign n913 = ( ~n148 & n311 ) | ( ~n148 & n912 ) | ( n311 & n912 ) ;
  assign n914 = n101 | n419 ;
  assign n915 = ( n874 & ~n894 ) | ( n874 & n914 ) | ( ~n894 & n914 ) ;
  assign n916 = n894 | n915 ;
  assign n917 = n450 ^ n179 ^ n136 ;
  assign n918 = n304 | n917 ;
  assign n919 = ( ~n267 & n413 ) | ( ~n267 & n917 ) | ( n413 & n917 ) ;
  assign n920 = n148 | n913 ;
  assign n921 = ( n203 & ~n481 ) | ( n203 & n920 ) | ( ~n481 & n920 ) ;
  assign n922 = n481 | n921 ;
  assign n923 = n267 | n919 ;
  assign n924 = ( n914 & ~n922 ) | ( n914 & n923 ) | ( ~n922 & n923 ) ;
  assign n925 = n922 | n924 ;
  assign n926 = ( ~n573 & n802 ) | ( ~n573 & n925 ) | ( n802 & n925 ) ;
  assign n927 = ( n173 & n212 ) | ( n173 & ~n357 ) | ( n212 & ~n357 ) ;
  assign n928 = n573 | n926 ;
  assign n929 = n264 | n488 ;
  assign n930 = ( n335 & ~n720 ) | ( n335 & n929 ) | ( ~n720 & n929 ) ;
  assign n931 = n720 | n930 ;
  assign n932 = n586 | n931 ;
  assign n933 = ( n869 & n918 ) | ( n869 & ~n932 ) | ( n918 & ~n932 ) ;
  assign n934 = n357 | n927 ;
  assign n935 = ~n493 & n734 ;
  assign n936 = n932 | n933 ;
  assign n937 = n187 | n395 ;
  assign n938 = ( ~n934 & n935 ) | ( ~n934 & n937 ) | ( n935 & n937 ) ;
  assign n939 = ~n937 & n938 ;
  assign n940 = ( n728 & ~n907 ) | ( n728 & n939 ) | ( ~n907 & n939 ) ;
  assign n941 = ~n728 & n940 ;
  assign n942 = n117 | n311 ;
  assign n943 = n217 | n222 ;
  assign n944 = ( n934 & n942 ) | ( n934 & ~n943 ) | ( n942 & ~n943 ) ;
  assign n945 = n114 | n180 ;
  assign n946 = n943 | n944 ;
  assign n947 = n392 | n945 ;
  assign n948 = n675 | n947 ;
  assign n949 = ( n556 & n891 ) | ( n556 & ~n948 ) | ( n891 & ~n948 ) ;
  assign n950 = n948 | n949 ;
  assign n951 = ( ~n908 & n946 ) | ( ~n908 & n948 ) | ( n946 & n948 ) ;
  assign n952 = n908 | n951 ;
  assign n953 = ( ~n323 & n861 ) | ( ~n323 & n952 ) | ( n861 & n952 ) ;
  assign n954 = ( ~n133 & n323 ) | ( ~n133 & n953 ) | ( n323 & n953 ) ;
  assign n955 = ( ~n187 & n227 ) | ( ~n187 & n459 ) | ( n227 & n459 ) ;
  assign n956 = n493 | n754 ;
  assign n957 = n187 | n955 ;
  assign n958 = ( n352 & ~n411 ) | ( n352 & n957 ) | ( ~n411 & n957 ) ;
  assign n959 = n411 | n958 ;
  assign n960 = ( n189 & ~n482 ) | ( n189 & n936 ) | ( ~n482 & n936 ) ;
  assign n961 = n176 | n901 ;
  assign n962 = ( ~n234 & n356 ) | ( ~n234 & n478 ) | ( n356 & n478 ) ;
  assign n963 = n117 | n175 ;
  assign n964 = ( n961 & n962 ) | ( n961 & ~n963 ) | ( n962 & ~n963 ) ;
  assign n965 = n963 | n964 ;
  assign n966 = n482 | n960 ;
  assign n967 = ( ~n160 & n230 ) | ( ~n160 & n965 ) | ( n230 & n965 ) ;
  assign n968 = ( ~n217 & n392 ) | ( ~n217 & n966 ) | ( n392 & n966 ) ;
  assign n969 = n160 | n967 ;
  assign n970 = n217 | n968 ;
  assign n971 = ( ~n672 & n749 ) | ( ~n672 & n969 ) | ( n749 & n969 ) ;
  assign n972 = ~n969 & n971 ;
  assign n973 = n956 | n959 ;
  assign n974 = ( n626 & ~n837 ) | ( n626 & n972 ) | ( ~n837 & n972 ) ;
  assign n975 = ~n968 & n974 ;
  assign n976 = n359 | n392 ;
  assign n977 = n541 | n976 ;
  assign n978 = n883 | n977 ;
  assign n979 = ~n217 & n975 ;
  assign n980 = ( ~n366 & n626 ) | ( ~n366 & n979 ) | ( n626 & n979 ) ;
  assign n981 = ~n626 & n980 ;
  assign n982 = ( ~n784 & n959 ) | ( ~n784 & n978 ) | ( n959 & n978 ) ;
  assign n983 = n784 | n982 ;
  assign n984 = ( n163 & n258 ) | ( n163 & ~n359 ) | ( n258 & ~n359 ) ;
  assign n985 = n359 | n984 ;
  assign n986 = n147 | n884 ;
  assign n987 = n173 | n325 ;
  assign n988 = ( n843 & n946 ) | ( n843 & ~n985 ) | ( n946 & ~n985 ) ;
  assign n989 = n177 | n513 ;
  assign n990 = ( n833 & ~n970 ) | ( n833 & n989 ) | ( ~n970 & n989 ) ;
  assign n991 = n970 | n990 ;
  assign n992 = ( ~n170 & n986 ) | ( ~n170 & n991 ) | ( n986 & n991 ) ;
  assign n993 = n986 | n987 ;
  assign n994 = ( ~n360 & n969 ) | ( ~n360 & n983 ) | ( n969 & n983 ) ;
  assign n995 = n117 | n273 ;
  assign n996 = n203 | n369 ;
  assign n997 = ( n85 & n995 ) | ( n85 & n996 ) | ( n995 & n996 ) ;
  assign n998 = ( ~n309 & n523 ) | ( ~n309 & n997 ) | ( n523 & n997 ) ;
  assign n999 = n309 | n998 ;
  assign n1000 = ( n660 & n892 ) | ( n660 & ~n999 ) | ( n892 & ~n999 ) ;
  assign n1001 = ( n754 & ~n785 ) | ( n754 & n999 ) | ( ~n785 & n999 ) ;
  assign n1002 = n300 | n478 ;
  assign n1003 = n785 | n1001 ;
  assign n1004 = n393 | n997 ;
  assign n1005 = ( n124 & ~n993 ) | ( n124 & n1004 ) | ( ~n993 & n1004 ) ;
  assign n1006 = n999 | n1000 ;
  assign n1007 = ( ~n391 & n970 ) | ( ~n391 & n1006 ) | ( n970 & n1006 ) ;
  assign n1008 = ( n628 & ~n1002 ) | ( n628 & n1003 ) | ( ~n1002 & n1003 ) ;
  assign n1009 = n1002 | n1008 ;
  assign n1010 = ( n156 & ~n931 ) | ( n156 & n1009 ) | ( ~n931 & n1009 ) ;
  assign n1011 = n993 | n1005 ;
  assign n1012 = n391 | n1007 ;
  assign n1013 = ( n614 & ~n719 ) | ( n614 & n1011 ) | ( ~n719 & n1011 ) ;
  assign n1014 = n719 | n1013 ;
  assign n1015 = n159 | n397 ;
  assign n1016 = n393 | n807 ;
  assign n1017 = n211 | n1015 ;
  assign n1018 = n117 | n408 ;
  assign n1019 = n220 | n396 ;
  assign n1020 = n528 | n1017 ;
  assign n1021 = n720 | n866 ;
  assign n1022 = ( n255 & ~n514 ) | ( n255 & n1014 ) | ( ~n514 & n1014 ) ;
  assign n1023 = ( ~n266 & n459 ) | ( ~n266 & n1021 ) | ( n459 & n1021 ) ;
  assign n1024 = n514 | n1022 ;
  assign n1025 = ( ~n408 & n459 ) | ( ~n408 & n1024 ) | ( n459 & n1024 ) ;
  assign n1026 = n272 | n514 ;
  assign n1027 = n1019 | n1026 ;
  assign n1028 = ( n225 & ~n1020 ) | ( n225 & n1027 ) | ( ~n1020 & n1027 ) ;
  assign n1029 = n1020 | n1028 ;
  assign n1030 = n160 | n213 ;
  assign n1031 = ( ~n133 & n1016 ) | ( ~n133 & n1018 ) | ( n1016 & n1018 ) ;
  assign n1032 = n1018 | n1030 ;
  assign n1033 = ( n447 & ~n460 ) | ( n447 & n1032 ) | ( ~n460 & n1032 ) ;
  assign n1034 = n460 | n1033 ;
  assign n1035 = n315 | n993 ;
  assign n1036 = ( ~n378 & n738 ) | ( ~n378 & n1034 ) | ( n738 & n1034 ) ;
  assign n1037 = n985 | n988 ;
  assign n1038 = n378 | n1036 ;
  assign n1039 = ( ~n303 & n426 ) | ( ~n303 & n1038 ) | ( n426 & n1038 ) ;
  assign n1040 = ( ~n400 & n950 ) | ( ~n400 & n1037 ) | ( n950 & n1037 ) ;
  assign n1041 = ~n267 & n734 ;
  assign n1042 = n266 | n1023 ;
  assign n1043 = ( n315 & n1029 ) | ( n315 & ~n1034 ) | ( n1029 & ~n1034 ) ;
  assign n1044 = n296 & ~n1043 ;
  assign n1045 = ~n230 & n1044 ;
  assign n1046 = ( ~n307 & n1034 ) | ( ~n307 & n1045 ) | ( n1034 & n1045 ) ;
  assign n1047 = ~n1002 & n1041 ;
  assign n1048 = ~n747 & n1046 ;
  assign n1049 = n303 | n1017 ;
  assign n1050 = n164 | n1049 ;
  assign n1051 = n189 | n440 ;
  assign n1052 = n303 | n1039 ;
  assign n1053 = n875 | n1052 ;
  assign n1054 = ( ~n164 & n1051 ) | ( ~n164 & n1053 ) | ( n1051 & n1053 ) ;
  assign n1055 = n164 | n1054 ;
  assign n1056 = n266 | n1017 ;
  assign n1057 = ( n347 & ~n784 ) | ( n347 & n1055 ) | ( ~n784 & n1055 ) ;
  assign n1058 = n784 | n1057 ;
  assign n1059 = n230 | n270 ;
  assign n1060 = ( ~n320 & n349 ) | ( ~n320 & n1059 ) | ( n349 & n1059 ) ;
  assign n1061 = n320 | n1060 ;
  assign n1062 = ~n1034 & n1048 ;
  assign n1063 = n147 | n311 ;
  assign n1064 = n1047 & ~n1063 ;
  assign n1065 = ( ~n335 & n1026 ) | ( ~n335 & n1061 ) | ( n1026 & n1061 ) ;
  assign n1066 = n335 | n1065 ;
  assign n1067 = ( ~n950 & n973 ) | ( ~n950 & n1066 ) | ( n973 & n1066 ) ;
  assign n1068 = n950 | n1067 ;
  assign n1069 = ( ~n266 & n1052 ) | ( ~n266 & n1068 ) | ( n1052 & n1068 ) ;
  assign n1070 = n266 | n1069 ;
  assign n1071 = n335 | n1063 ;
  assign n1072 = ( ~n315 & n644 ) | ( ~n315 & n1071 ) | ( n644 & n1071 ) ;
  assign n1073 = n315 | n1072 ;
  assign n1074 = ( ~n396 & n483 ) | ( ~n396 & n1073 ) | ( n483 & n1073 ) ;
  assign n1075 = n396 | n1074 ;
  assign n1076 = ( n168 & ~n212 ) | ( n168 & n1075 ) | ( ~n212 & n1075 ) ;
  assign n1077 = ( n349 & ~n1056 ) | ( n349 & n1063 ) | ( ~n1056 & n1063 ) ;
  assign n1078 = n1056 | n1077 ;
  assign n1079 = ( ~n366 & n985 ) | ( ~n366 & n1078 ) | ( n985 & n1078 ) ;
  assign n1080 = n366 | n1079 ;
  assign n1081 = ( ~n187 & n213 ) | ( ~n187 & n1080 ) | ( n213 & n1080 ) ;
  assign n1082 = n584 | n914 ;
  assign n1083 = n187 | n1081 ;
  assign n1084 = ( n394 & ~n433 ) | ( n394 & n1083 ) | ( ~n433 & n1083 ) ;
  assign n1085 = n433 | n1084 ;
  assign n1086 = ( n297 & ~n369 ) | ( n297 & n584 ) | ( ~n369 & n584 ) ;
  assign n1087 = n369 | n1086 ;
  assign n1088 = ( ~n440 & n1002 ) | ( ~n440 & n1087 ) | ( n1002 & n1087 ) ;
  assign n1089 = n218 | n1085 ;
  assign n1090 = ( ~n440 & n487 ) | ( ~n440 & n1089 ) | ( n487 & n1089 ) ;
  assign n1091 = n440 | n1088 ;
  assign n1092 = n440 | n1090 ;
  assign n1093 = n1053 | n1059 ;
  assign n1094 = n541 | n1002 ;
  assign n1095 = n122 | n481 ;
  assign n1096 = n541 | n1095 ;
  assign n1097 = ( n815 & ~n1093 ) | ( n815 & n1096 ) | ( ~n1093 & n1096 ) ;
  assign n1098 = n212 | n1076 ;
  assign n1099 = n1093 | n1097 ;
  assign n1100 = ( n624 & n644 ) | ( n624 & ~n778 ) | ( n644 & ~n778 ) ;
  assign n1101 = n187 | n188 ;
  assign n1102 = n388 | n644 ;
  assign n1103 = ( n483 & ~n1095 ) | ( n483 & n1102 ) | ( ~n1095 & n1102 ) ;
  assign n1104 = n1095 | n1103 ;
  assign n1105 = n181 | n699 ;
  assign n1106 = n261 | n397 ;
  assign n1107 = n837 | n878 ;
  assign n1108 = n393 | n699 ;
  assign n1109 = n401 | n1098 ;
  assign n1110 = ( ~n371 & n614 ) | ( ~n371 & n1108 ) | ( n614 & n1108 ) ;
  assign n1111 = ( ~n206 & n1027 ) | ( ~n206 & n1104 ) | ( n1027 & n1104 ) ;
  assign n1112 = ( n963 & n1095 ) | ( n963 & ~n1105 ) | ( n1095 & ~n1105 ) ;
  assign n1113 = n141 | n311 ;
  assign n1114 = n963 | n1106 ;
  assign n1115 = n1105 | n1112 ;
  assign n1116 = ( ~n366 & n1101 ) | ( ~n366 & n1113 ) | ( n1101 & n1113 ) ;
  assign n1117 = ( n297 & n1050 ) | ( n297 & ~n1115 ) | ( n1050 & ~n1115 ) ;
  assign n1118 = n1115 | n1117 ;
  assign n1119 = n366 | n1098 ;
  assign n1120 = n366 | n1116 ;
  assign n1121 = ( n610 & ~n1099 ) | ( n610 & n1120 ) | ( ~n1099 & n1120 ) ;
  assign n1122 = n309 | n502 ;
  assign n1123 = n1099 | n1121 ;
  assign n1124 = ( n734 & ~n837 ) | ( n734 & n1123 ) | ( ~n837 & n1123 ) ;
  assign n1125 = ( ~n654 & n1120 ) | ( ~n654 & n1122 ) | ( n1120 & n1122 ) ;
  assign n1126 = n654 | n1125 ;
  assign n1127 = ( ~n416 & n1114 ) | ( ~n416 & n1126 ) | ( n1114 & n1126 ) ;
  assign n1128 = n419 ^ n203 ^ n133 ;
  assign n1129 = n734 & ~n1128 ;
  assign n1130 = ( n497 & ~n1085 ) | ( n497 & n1129 ) | ( ~n1085 & n1129 ) ;
  assign n1131 = ( ~n676 & n1123 ) | ( ~n676 & n1124 ) | ( n1123 & n1124 ) ;
  assign n1132 = ~n497 & n1130 ;
  assign n1133 = ~n1123 & n1131 ;
  assign n1134 = ( ~n416 & n1094 ) | ( ~n416 & n1127 ) | ( n1094 & n1127 ) ;
  assign n1135 = n139 | n146 ;
  assign n1136 = ( ~n411 & n460 ) | ( ~n411 & n1135 ) | ( n460 & n1135 ) ;
  assign n1137 = n411 | n1136 ;
  assign n1138 = ( ~n353 & n438 ) | ( ~n353 & n1137 ) | ( n438 & n1137 ) ;
  assign n1139 = n353 | n1138 ;
  assign n1140 = n931 | n1010 ;
  assign n1141 = ( ~n115 & n325 ) | ( ~n115 & n1139 ) | ( n325 & n1139 ) ;
  assign n1142 = ( ~n438 & n989 ) | ( ~n438 & n1140 ) | ( n989 & n1140 ) ;
  assign n1143 = n438 | n1142 ;
  assign n1144 = n115 | n1141 ;
  assign n1145 = ( n114 & ~n1128 ) | ( n114 & n1144 ) | ( ~n1128 & n1144 ) ;
  assign n1146 = n1128 | n1145 ;
  assign n1147 = ( ~n184 & n483 ) | ( ~n184 & n1146 ) | ( n483 & n1146 ) ;
  assign n1148 = n184 | n1147 ;
  assign n1149 = n174 | n441 ;
  assign n1150 = n388 | n1149 ;
  assign n1151 = ( ~n416 & n447 ) | ( ~n416 & n1148 ) | ( n447 & n1148 ) ;
  assign n1152 = ( n179 & ~n514 ) | ( n179 & n870 ) | ( ~n514 & n870 ) ;
  assign n1153 = n514 | n1152 ;
  assign n1154 = ( ~n416 & n1134 ) | ( ~n416 & n1151 ) | ( n1134 & n1151 ) ;
  assign n1155 = n416 | n1151 ;
  assign n1156 = n326 | n1155 ;
  assign n1157 = n348 | n528 ;
  assign n1158 = n922 | n1144 ;
  assign n1159 = n348 | n394 ;
  assign n1160 = ( ~n395 & n1149 ) | ( ~n395 & n1159 ) | ( n1149 & n1159 ) ;
  assign n1161 = n395 | n1160 ;
  assign n1162 = ( n343 & ~n785 ) | ( n343 & n1161 ) | ( ~n785 & n1161 ) ;
  assign n1163 = n785 | n1162 ;
  assign n1164 = ( ~n532 & n900 ) | ( ~n532 & n1163 ) | ( n900 & n1163 ) ;
  assign n1165 = ( n511 & ~n514 ) | ( n511 & n1158 ) | ( ~n514 & n1158 ) ;
  assign n1166 = ( ~n676 & n1064 ) | ( ~n676 & n1163 ) | ( n1064 & n1163 ) ;
  assign n1167 = ~n1163 & n1166 ;
  assign n1168 = ( ~n369 & n476 ) | ( ~n369 & n1157 ) | ( n476 & n1157 ) ;
  assign n1169 = n416 | n1154 ;
  assign n1170 = n671 | n1149 ;
  assign n1171 = ( ~n174 & n347 ) | ( ~n174 & n1169 ) | ( n347 & n1169 ) ;
  assign n1172 = n514 | n1165 ;
  assign n1173 = ( n1066 & ~n1156 ) | ( n1066 & n1170 ) | ( ~n1156 & n1170 ) ;
  assign n1174 = n174 | n1171 ;
  assign n1175 = ( ~n270 & n512 ) | ( ~n270 & n1174 ) | ( n512 & n1174 ) ;
  assign n1176 = n270 | n1175 ;
  assign n1177 = ( ~n147 & n182 ) | ( ~n147 & n1176 ) | ( n182 & n1176 ) ;
  assign n1178 = n147 | n1177 ;
  assign n1179 = n1156 | n1173 ;
  assign n1180 = ( ~n224 & n476 ) | ( ~n224 & n1178 ) | ( n476 & n1178 ) ;
  assign n1181 = ( ~n148 & n290 ) | ( ~n148 & n1179 ) | ( n290 & n1179 ) ;
  assign n1182 = n148 | n1181 ;
  assign n1183 = ( n148 & ~n159 ) | ( n148 & n1012 ) | ( ~n159 & n1012 ) ;
  assign n1184 = n753 | n815 ;
  assign n1185 = n532 | n1164 ;
  assign n1186 = n148 | n213 ;
  assign n1187 = ( ~n133 & n273 ) | ( ~n133 & n1186 ) | ( n273 & n1186 ) ;
  assign n1188 = n133 | n1187 ;
  assign n1189 = ( ~n175 & n320 ) | ( ~n175 & n356 ) | ( n320 & n356 ) ;
  assign n1190 = n175 | n1189 ;
  assign n1191 = ( ~n170 & n408 ) | ( ~n170 & n1190 ) | ( n408 & n1190 ) ;
  assign n1192 = n176 | n428 ;
  assign n1193 = n170 | n1191 ;
  assign n1194 = ( ~n723 & n1188 ) | ( ~n723 & n1193 ) | ( n1188 & n1193 ) ;
  assign n1195 = n723 | n1194 ;
  assign n1196 = ( n511 & ~n753 ) | ( n511 & n931 ) | ( ~n753 & n931 ) ;
  assign n1197 = n753 | n1196 ;
  assign n1198 = ( ~n125 & n585 ) | ( ~n125 & n1195 ) | ( n585 & n1195 ) ;
  assign n1199 = n125 | n1198 ;
  assign n1200 = ( ~n937 & n1059 ) | ( ~n937 & n1199 ) | ( n1059 & n1199 ) ;
  assign n1201 = n937 | n1200 ;
  assign n1202 = n450 | n482 ;
  assign n1203 = ( n184 & ~n399 ) | ( n184 & n1202 ) | ( ~n399 & n1202 ) ;
  assign n1204 = n125 | n560 ;
  assign n1205 = ( n753 & ~n778 ) | ( n753 & n1204 ) | ( ~n778 & n1204 ) ;
  assign n1206 = ( n175 & ~n481 ) | ( n175 & n1192 ) | ( ~n481 & n1192 ) ;
  assign n1207 = n399 | n1203 ;
  assign n1208 = ( ~n263 & n976 ) | ( ~n263 & n1207 ) | ( n976 & n1207 ) ;
  assign n1209 = n263 | n1208 ;
  assign n1210 = n133 | n300 ;
  assign n1211 = n778 | n1205 ;
  assign n1212 = ( ~n558 & n1201 ) | ( ~n558 & n1209 ) | ( n1201 & n1209 ) ;
  assign n1213 = n481 | n1206 ;
  assign n1214 = n558 | n1212 ;
  assign n1215 = ( n532 & n1197 ) | ( n532 & ~n1213 ) | ( n1197 & ~n1213 ) ;
  assign n1216 = ( ~n1106 & n1195 ) | ( ~n1106 & n1211 ) | ( n1195 & n1211 ) ;
  assign n1217 = n1106 | n1216 ;
  assign n1218 = ( n311 & ~n679 ) | ( n311 & n1217 ) | ( ~n679 & n1217 ) ;
  assign n1219 = n679 | n1218 ;
  assign n1220 = n1213 | n1215 ;
  assign n1221 = ( n356 & ~n357 ) | ( n356 & n1220 ) | ( ~n357 & n1220 ) ;
  assign n1222 = n357 | n1221 ;
  assign n1223 = ( n353 & ~n677 ) | ( n353 & n1222 ) | ( ~n677 & n1222 ) ;
  assign n1224 = ( ~n426 & n677 ) | ( ~n426 & n1223 ) | ( n677 & n1223 ) ;
  assign n1225 = n426 | n1224 ;
  assign n1226 = ( n1113 & ~n1210 ) | ( n1113 & n1225 ) | ( ~n1210 & n1225 ) ;
  assign n1227 = n1210 | n1226 ;
  assign n1228 = n1209 | n1227 ;
  assign n1229 = ( n999 & n1035 ) | ( n999 & ~n1228 ) | ( n1035 & ~n1228 ) ;
  assign n1230 = n1228 | n1229 ;
  assign n1231 = ( ~n216 & n564 ) | ( ~n216 & n1230 ) | ( n564 & n1230 ) ;
  assign n1232 = n216 | n1231 ;
  assign n1233 = ( ~n778 & n1100 ) | ( ~n778 & n1225 ) | ( n1100 & n1225 ) ;
  assign n1234 = n778 | n1233 ;
  assign n1235 = ( n114 & ~n394 ) | ( n114 & n1232 ) | ( ~n394 & n1232 ) ;
  assign n1236 = ( ~n441 & n468 ) | ( ~n441 & n928 ) | ( n468 & n928 ) ;
  assign n1237 = ( n356 & ~n360 ) | ( n356 & n1143 ) | ( ~n360 & n1143 ) ;
  assign n1238 = n360 | n1237 ;
  assign n1239 = n369 | n1168 ;
  assign n1240 = ( ~n175 & n273 ) | ( ~n175 & n1238 ) | ( n273 & n1238 ) ;
  assign n1241 = ( ~n400 & n604 ) | ( ~n400 & n1040 ) | ( n604 & n1040 ) ;
  assign n1242 = n441 | n1236 ;
  assign n1243 = ( n230 & ~n299 ) | ( n230 & n1242 ) | ( ~n299 & n1242 ) ;
  assign n1244 = n230 | n233 ;
  assign n1245 = n175 | n1240 ;
  assign n1246 = n261 | n301 ;
  assign n1247 = n433 | n893 ;
  assign n1248 = n136 | n433 ;
  assign n1249 = ( ~n307 & n604 ) | ( ~n307 & n1246 ) | ( n604 & n1246 ) ;
  assign n1250 = n307 | n1249 ;
  assign n1251 = n413 | n1250 ;
  assign n1252 = n408 | n1025 ;
  assign n1253 = n378 | n1106 ;
  assign n1254 = ( ~n720 & n1132 ) | ( ~n720 & n1251 ) | ( n1132 & n1251 ) ;
  assign n1255 = n976 | n1128 ;
  assign n1256 = ~n1251 & n1254 ;
  assign n1257 = n312 | n408 ;
  assign n1258 = ( n178 & ~n441 ) | ( n178 & n488 ) | ( ~n441 & n488 ) ;
  assign n1259 = ( n238 & ~n513 ) | ( n238 & n1257 ) | ( ~n513 & n1257 ) ;
  assign n1260 = n513 | n1259 ;
  assign n1261 = ( ~n273 & n356 ) | ( ~n273 & n1256 ) | ( n356 & n1256 ) ;
  assign n1262 = ~n356 & n1261 ;
  assign n1263 = ( ~n117 & n212 ) | ( ~n117 & n1262 ) | ( n212 & n1262 ) ;
  assign n1264 = ( n212 & ~n290 ) | ( n212 & n1263 ) | ( ~n290 & n1263 ) ;
  assign n1265 = n220 | n1248 ;
  assign n1266 = ( ~n187 & n416 ) | ( ~n187 & n1265 ) | ( n416 & n1265 ) ;
  assign n1267 = n187 | n1266 ;
  assign n1268 = ( ~n1253 & n1255 ) | ( ~n1253 & n1267 ) | ( n1255 & n1267 ) ;
  assign n1269 = ( n732 & ~n905 ) | ( n732 & n1267 ) | ( ~n905 & n1267 ) ;
  assign n1270 = n441 | n1258 ;
  assign n1271 = ( ~n117 & n395 ) | ( ~n117 & n1270 ) | ( n395 & n1270 ) ;
  assign n1272 = n117 | n1271 ;
  assign n1273 = n1253 | n1268 ;
  assign n1274 = ( n1107 & ~n1260 ) | ( n1107 & n1272 ) | ( ~n1260 & n1272 ) ;
  assign n1275 = n182 | n800 ;
  assign n1276 = ( ~n258 & n408 ) | ( ~n258 & n460 ) | ( n408 & n460 ) ;
  assign n1277 = n905 | n1269 ;
  assign n1278 = ( n800 & ~n985 ) | ( n800 & n1272 ) | ( ~n985 & n1272 ) ;
  assign n1279 = ( n361 & ~n773 ) | ( n361 & n1275 ) | ( ~n773 & n1275 ) ;
  assign n1280 = n258 | n1276 ;
  assign n1281 = ( ~n945 & n1239 ) | ( ~n945 & n1280 ) | ( n1239 & n1280 ) ;
  assign n1282 = n945 | n1281 ;
  assign n1283 = n1260 | n1274 ;
  assign n1284 = ( ~n720 & n1155 ) | ( ~n720 & n1283 ) | ( n1155 & n1283 ) ;
  assign n1285 = ( ~n181 & n1244 ) | ( ~n181 & n1280 ) | ( n1244 & n1280 ) ;
  assign n1286 = n181 | n1285 ;
  assign n1287 = ( ~n1213 & n1273 ) | ( ~n1213 & n1286 ) | ( n1273 & n1286 ) ;
  assign n1288 = n985 | n1278 ;
  assign n1289 = ( n1030 & ~n1213 ) | ( n1030 & n1287 ) | ( ~n1213 & n1287 ) ;
  assign n1290 = n720 | n1284 ;
  assign n1291 = ( n189 & ~n273 ) | ( n189 & n1290 ) | ( ~n273 & n1290 ) ;
  assign n1292 = n273 | n1291 ;
  assign n1293 = ( ~n255 & n369 ) | ( ~n255 & n1292 ) | ( n369 & n1292 ) ;
  assign n1294 = n255 | n1293 ;
  assign n1295 = ( n222 & ~n272 ) | ( n222 & n1294 ) | ( ~n272 & n1294 ) ;
  assign n1296 = ( ~n272 & n300 ) | ( ~n272 & n1295 ) | ( n300 & n1295 ) ;
  assign n1297 = n272 | n1296 ;
  assign n1298 = n1213 | n1289 ;
  assign n1299 = ( n221 & ~n426 ) | ( n221 & n1298 ) | ( ~n426 & n1298 ) ;
  assign n1300 = n426 | n1299 ;
  assign n1301 = ( ~n931 & n1167 ) | ( ~n931 & n1300 ) | ( n1167 & n1300 ) ;
  assign n1302 = ( n134 & ~n360 ) | ( n134 & n394 ) | ( ~n360 & n394 ) ;
  assign n1303 = n360 | n1302 ;
  assign n1304 = ~n1300 & n1301 ;
  assign n1305 = ( ~n237 & n478 ) | ( ~n237 & n828 ) | ( n478 & n828 ) ;
  assign n1306 = n237 | n1305 ;
  assign n1307 = ( n331 & ~n511 ) | ( n331 & n1304 ) | ( ~n511 & n1304 ) ;
  assign n1308 = ~n331 & n1307 ;
  assign n1309 = ( ~n234 & n255 ) | ( ~n234 & n1308 ) | ( n255 & n1308 ) ;
  assign n1310 = n206 | n1111 ;
  assign n1311 = n146 | n513 ;
  assign n1312 = ~n255 & n1309 ;
  assign n1313 = ( n101 & ~n117 ) | ( n101 & n1312 ) | ( ~n117 & n1312 ) ;
  assign n1314 = n184 | n229 ;
  assign n1315 = n502 ^ n255 ^ n188 ;
  assign n1316 = n773 | n1279 ;
  assign n1317 = ( ~n115 & n1303 ) | ( ~n115 & n1315 ) | ( n1303 & n1315 ) ;
  assign n1318 = n115 | n1317 ;
  assign n1319 = ( n1213 & ~n1316 ) | ( n1213 & n1318 ) | ( ~n1316 & n1318 ) ;
  assign n1320 = n1316 | n1319 ;
  assign n1321 = ( ~n216 & n299 ) | ( ~n216 & n1320 ) | ( n299 & n1320 ) ;
  assign n1322 = n216 | n1321 ;
  assign n1323 = ( n378 & ~n647 ) | ( n378 & n1322 ) | ( ~n647 & n1322 ) ;
  assign n1324 = ( n831 & ~n1311 ) | ( n831 & n1315 ) | ( ~n1311 & n1315 ) ;
  assign n1325 = n1311 | n1324 ;
  assign n1326 = ( ~n1150 & n1314 ) | ( ~n1150 & n1325 ) | ( n1314 & n1325 ) ;
  assign n1327 = n1150 | n1326 ;
  assign n1328 = ( n349 & ~n356 ) | ( n349 & n1327 ) | ( ~n356 & n1327 ) ;
  assign n1329 = ~n101 & n1313 ;
  assign n1330 = n647 | n1323 ;
  assign n1331 = n110 | n125 ;
  assign n1332 = n356 | n1328 ;
  assign n1333 = ( n177 & ~n234 ) | ( n177 & n1332 ) | ( ~n234 & n1332 ) ;
  assign n1334 = n234 | n1333 ;
  assign n1335 = ( n1234 & n1286 ) | ( n1234 & ~n1318 ) | ( n1286 & ~n1318 ) ;
  assign n1336 = n511 | n1334 ;
  assign n1337 = ( n206 & ~n1109 ) | ( n206 & n1336 ) | ( ~n1109 & n1336 ) ;
  assign n1338 = n1109 | n1337 ;
  assign n1339 = n1318 | n1335 ;
  assign n1340 = ( ~n216 & n941 ) | ( ~n216 & n1321 ) | ( n941 & n1321 ) ;
  assign n1341 = ( n189 & ~n512 ) | ( n189 & n1338 ) | ( ~n512 & n1338 ) ;
  assign n1342 = ~n1321 & n1340 ;
  assign n1343 = n108 & ~n1334 ;
  assign n1344 = ( ~n125 & n1306 ) | ( ~n125 & n1342 ) | ( n1306 & n1342 ) ;
  assign n1345 = ( n149 & ~n880 ) | ( n149 & n1343 ) | ( ~n880 & n1343 ) ;
  assign n1346 = ~n1306 & n1344 ;
  assign n1347 = ( n135 & ~n441 ) | ( n135 & n1346 ) | ( ~n441 & n1346 ) ;
  assign n1348 = ~n135 & n1347 ;
  assign n1349 = ( ~n137 & n1306 ) | ( ~n137 & n1331 ) | ( n1306 & n1331 ) ;
  assign n1350 = ~n149 & n1345 ;
  assign n1351 = ( n891 & ~n1286 ) | ( n891 & n1350 ) | ( ~n1286 & n1350 ) ;
  assign n1352 = ~n891 & n1351 ;
  assign n1353 = ( ~n136 & n238 ) | ( ~n136 & n1348 ) | ( n238 & n1348 ) ;
  assign n1354 = ( n132 & ~n488 ) | ( n132 & n1058 ) | ( ~n488 & n1058 ) ;
  assign n1355 = ( ~n634 & n884 ) | ( ~n634 & n1277 ) | ( n884 & n1277 ) ;
  assign n1356 = n349 | n773 ;
  assign n1357 = n234 | n393 ;
  assign n1358 = ( n460 & ~n634 ) | ( n460 & n1355 ) | ( ~n634 & n1355 ) ;
  assign n1359 = n634 | n1358 ;
  assign n1360 = ( ~n149 & n1356 ) | ( ~n149 & n1359 ) | ( n1356 & n1359 ) ;
  assign n1361 = n132 | n229 ;
  assign n1362 = n311 | n976 ;
  assign n1363 = ( ~n989 & n1359 ) | ( ~n989 & n1362 ) | ( n1359 & n1362 ) ;
  assign n1364 = n139 | n262 ;
  assign n1365 = ( n179 & ~n426 ) | ( n179 & n1364 ) | ( ~n426 & n1364 ) ;
  assign n1366 = n426 | n1365 ;
  assign n1367 = ( ~n335 & n343 ) | ( ~n335 & n1366 ) | ( n343 & n1366 ) ;
  assign n1368 = n335 | n1367 ;
  assign n1369 = ( ~n1082 & n1361 ) | ( ~n1082 & n1368 ) | ( n1361 & n1368 ) ;
  assign n1370 = n1082 | n1369 ;
  assign n1371 = ( n182 & ~n357 ) | ( n182 & n1370 ) | ( ~n357 & n1370 ) ;
  assign n1372 = n357 | n1371 ;
  assign n1373 = ( n224 & ~n271 ) | ( n224 & n1372 ) | ( ~n271 & n1372 ) ;
  assign n1374 = n271 | n1373 ;
  assign n1375 = ( n115 & ~n307 ) | ( n115 & n1374 ) | ( ~n307 & n1374 ) ;
  assign n1376 = n307 | n1375 ;
  assign n1377 = n181 | n217 ;
  assign n1378 = ( n1357 & n1376 ) | ( n1357 & ~n1377 ) | ( n1376 & ~n1377 ) ;
  assign n1379 = n1377 | n1378 ;
  assign n1380 = n468 | n1379 ;
  assign n1381 = ( n376 & n1184 ) | ( n376 & ~n1380 ) | ( n1184 & ~n1380 ) ;
  assign n1382 = n360 | n994 ;
  assign n1383 = n149 | n1360 ;
  assign n1384 = ( n1092 & n1260 ) | ( n1092 & ~n1376 ) | ( n1260 & ~n1376 ) ;
  assign n1385 = n1380 | n1381 ;
  assign n1386 = ( n331 & ~n349 ) | ( n331 & n1385 ) | ( ~n349 & n1385 ) ;
  assign n1387 = n989 | n1363 ;
  assign n1388 = n1376 | n1384 ;
  assign n1389 = ( ~n199 & n468 ) | ( ~n199 & n1388 ) | ( n468 & n1388 ) ;
  assign n1390 = n199 | n1389 ;
  assign n1391 = ( ~n141 & n309 ) | ( ~n141 & n1390 ) | ( n309 & n1390 ) ;
  assign n1392 = ( ~n1193 & n1379 ) | ( ~n1193 & n1387 ) | ( n1379 & n1387 ) ;
  assign n1393 = ( ~n149 & n376 ) | ( ~n149 & n1300 ) | ( n376 & n1300 ) ;
  assign n1394 = n149 | n1393 ;
  assign n1395 = n1193 | n1392 ;
  assign n1396 = ( ~n270 & n353 ) | ( ~n270 & n1395 ) | ( n353 & n1395 ) ;
  assign n1397 = n141 | n1391 ;
  assign n1398 = n270 | n1396 ;
  assign n1399 = n349 | n1386 ;
  assign n1400 = ( ~n146 & n360 ) | ( ~n146 & n1399 ) | ( n360 & n1399 ) ;
  assign n1401 = ( n199 & ~n444 ) | ( n199 & n1394 ) | ( ~n444 & n1394 ) ;
  assign n1402 = n444 | n1401 ;
  assign n1403 = ( n173 & ~n482 ) | ( n173 & n1397 ) | ( ~n482 & n1397 ) ;
  assign n1404 = ( ~n311 & n989 ) | ( ~n311 & n1402 ) | ( n989 & n1402 ) ;
  assign n1405 = n311 | n1404 ;
  assign n1406 = ( n262 & ~n482 ) | ( n262 & n1405 ) | ( ~n482 & n1405 ) ;
  assign n1407 = ( ~n299 & n996 ) | ( ~n299 & n1398 ) | ( n996 & n1398 ) ;
  assign n1408 = ( ~n488 & n512 ) | ( ~n488 & n1341 ) | ( n512 & n1341 ) ;
  assign n1409 = n488 | n1408 ;
  assign n1410 = ( n220 & ~n450 ) | ( n220 & n1118 ) | ( ~n450 & n1118 ) ;
  assign n1411 = ~n212 & n1264 ;
  assign n1412 = n137 | n1349 ;
  assign n1413 = n488 | n1354 ;
  assign n1414 = ( n212 & ~n481 ) | ( n212 & n1413 ) | ( ~n481 & n1413 ) ;
  assign n1415 = ( n221 & ~n481 ) | ( n221 & n1414 ) | ( ~n481 & n1414 ) ;
  assign n1416 = n481 | n1415 ;
  assign n1417 = n146 | n1400 ;
  assign n1418 = ( ~n180 & n395 ) | ( ~n180 & n1417 ) | ( n395 & n1417 ) ;
  assign n1419 = n180 | n1418 ;
  assign n1420 = ( ~n110 & n220 ) | ( ~n110 & n1419 ) | ( n220 & n1419 ) ;
  assign n1421 = n110 | n1420 ;
  assign n1422 = n482 | n1403 ;
  assign n1423 = ( n395 & ~n428 ) | ( n395 & n1422 ) | ( ~n428 & n1422 ) ;
  assign n1424 = ( ~n211 & n395 ) | ( ~n211 & n1091 ) | ( n395 & n1091 ) ;
  assign n1425 = ( ~n211 & n325 ) | ( ~n211 & n1424 ) | ( n325 & n1424 ) ;
  assign n1426 = n211 | n1425 ;
  assign n1427 = ( n673 & ~n1300 ) | ( n673 & n1426 ) | ( ~n1300 & n1426 ) ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1429 = ( ~n371 & n690 ) | ( ~n371 & n1426 ) | ( n690 & n1426 ) ;
  assign n1430 = n371 | n1429 ;
  assign n1431 = ( ~n213 & n221 ) | ( ~n213 & n512 ) | ( n221 & n512 ) ;
  assign n1432 = n213 | n1431 ;
  assign n1433 = ( ~n1250 & n1383 ) | ( ~n1250 & n1432 ) | ( n1383 & n1432 ) ;
  assign n1434 = n1250 | n1433 ;
  assign n1435 = n482 | n1406 ;
  assign n1436 = ( n1288 & n1368 ) | ( n1288 & ~n1412 ) | ( n1368 & ~n1412 ) ;
  assign n1437 = n1412 | n1436 ;
  assign n1438 = ( ~n276 & n1126 ) | ( ~n276 & n1437 ) | ( n1126 & n1437 ) ;
  assign n1439 = n276 | n1438 ;
  assign n1440 = ( ~n203 & n396 ) | ( ~n203 & n1439 ) | ( n396 & n1439 ) ;
  assign n1441 = ( n178 & ~n502 ) | ( n178 & n1434 ) | ( ~n502 & n1434 ) ;
  assign n1442 = n502 | n1441 ;
  assign n1443 = ( n224 & ~n581 ) | ( n224 & n1442 ) | ( ~n581 & n1442 ) ;
  assign n1444 = n581 | n1443 ;
  assign n1445 = ( n203 & ~n416 ) | ( n203 & n1440 ) | ( ~n416 & n1440 ) ;
  assign n1446 = n416 | n1445 ;
  assign n1447 = ( ~n159 & n235 ) | ( ~n159 & n1042 ) | ( n235 & n1042 ) ;
  assign n1448 = ( ~n159 & n307 ) | ( ~n159 & n1447 ) | ( n307 & n1447 ) ;
  assign n1449 = ( n883 & n1330 ) | ( n883 & ~n1432 ) | ( n1330 & ~n1432 ) ;
  assign n1450 = n1432 | n1449 ;
  assign n1451 = ( n184 & ~n301 ) | ( n184 & n1450 ) | ( ~n301 & n1450 ) ;
  assign n1452 = n371 | n1110 ;
  assign n1453 = ( n254 & ~n419 ) | ( n254 & n1153 ) | ( ~n419 & n1153 ) ;
  assign n1454 = ( n231 & ~n254 ) | ( n231 & n981 ) | ( ~n254 & n981 ) ;
  assign n1455 = ~n231 & n1454 ;
  assign n1456 = ( n133 & ~n211 ) | ( n133 & n1455 ) | ( ~n211 & n1455 ) ;
  assign n1457 = ( ~n301 & n399 ) | ( ~n301 & n1062 ) | ( n399 & n1062 ) ;
  assign n1458 = ~n399 & n1457 ;
  assign n1459 = ( n182 & ~n187 ) | ( n182 & n1458 ) | ( ~n187 & n1458 ) ;
  assign n1460 = ( ~n271 & n301 ) | ( ~n271 & n1339 ) | ( n301 & n1339 ) ;
  assign n1461 = ( ~n237 & n271 ) | ( ~n237 & n1460 ) | ( n271 & n1460 ) ;
  assign n1462 = ( ~n182 & n335 ) | ( ~n182 & n1185 ) | ( n335 & n1185 ) ;
  assign n1463 = n182 | n1462 ;
  assign n1464 = ( n179 & ~n188 ) | ( n179 & n1463 ) | ( ~n188 & n1463 ) ;
  assign n1465 = n400 | n1241 ;
  assign n1466 = ( ~n188 & n512 ) | ( ~n188 & n1465 ) | ( n512 & n1465 ) ;
  assign n1467 = ( ~n884 & n1248 ) | ( ~n884 & n1352 ) | ( n1248 & n1352 ) ;
  assign n1468 = ~n1248 & n1467 ;
  assign n1469 = ( n392 & ~n428 ) | ( n392 & n916 ) | ( ~n428 & n916 ) ;
  assign n1470 = n428 | n1469 ;
  assign n1471 = n610 | n1470 ;
  assign n1472 = ( n334 & ~n1248 ) | ( n334 & n1471 ) | ( ~n1248 & n1471 ) ;
  assign n1473 = ~n1471 & n1472 ;
  assign n1474 = ( ~n229 & n512 ) | ( ~n229 & n1473 ) | ( n512 & n1473 ) ;
  assign n1475 = ~n512 & n1474 ;
  assign n1476 = ( ~n224 & n352 ) | ( ~n224 & n1475 ) | ( n352 & n1475 ) ;
  assign n1477 = ~n352 & n1476 ;
  assign n1478 = ( ~n237 & n884 ) | ( ~n237 & n1428 ) | ( n884 & n1428 ) ;
  assign n1479 = ~n884 & n1478 ;
  assign n1480 = ( n271 & ~n303 ) | ( n271 & n392 ) | ( ~n303 & n392 ) ;
  assign n1481 = n303 | n1480 ;
  assign n1482 = ( n335 & ~n393 ) | ( n335 & n1481 ) | ( ~n393 & n1481 ) ;
  assign n1483 = n393 | n1482 ;
  assign n1484 = ( ~n1172 & n1412 ) | ( ~n1172 & n1483 ) | ( n1412 & n1483 ) ;
  assign n1485 = n1172 | n1484 ;
  assign n1486 = ( ~n400 & n1214 ) | ( ~n400 & n1248 ) | ( n1214 & n1248 ) ;
  assign n1487 = n400 | n1486 ;
  assign n1488 = ( n163 & ~n178 ) | ( n163 & n1487 ) | ( ~n178 & n1487 ) ;
  assign n1489 = ( n134 & ~n178 ) | ( n134 & n1488 ) | ( ~n178 & n1488 ) ;
  assign n1490 = ( n1430 & n1432 ) | ( n1430 & ~n1483 ) | ( n1432 & ~n1483 ) ;
  assign n1491 = n1483 | n1490 ;
  assign n1492 = ( ~n126 & n210 ) | ( ~n126 & n1491 ) | ( n210 & n1491 ) ;
  assign n1493 = n126 | n1492 ;
  assign n1494 = ( ~n634 & n1260 ) | ( ~n634 & n1493 ) | ( n1260 & n1493 ) ;
  assign n1495 = n634 | n1494 ;
  assign n1496 = ( n163 & ~n264 ) | ( n163 & n1495 ) | ( ~n264 & n1495 ) ;
  assign n1497 = n264 | n1496 ;
  assign n1498 = ( n216 & ~n419 ) | ( n216 & n1497 ) | ( ~n419 & n1497 ) ;
  assign n1499 = ( ~n254 & n411 ) | ( ~n254 & n1435 ) | ( n411 & n1435 ) ;
  assign n1500 = n254 | n1499 ;
  assign n1501 = ( ~n115 & n447 ) | ( ~n115 & n1500 ) | ( n447 & n1500 ) ;
  assign n1502 = n115 | n1501 ;
  assign n1503 = ( n179 & ~n271 ) | ( n179 & n1382 ) | ( ~n271 & n1382 ) ;
  assign n1504 = n271 | n1503 ;
  assign n1505 = ( ~n258 & n447 ) | ( ~n258 & n1504 ) | ( n447 & n1504 ) ;
  assign n1506 = ( n233 & ~n258 ) | ( n233 & n1505 ) | ( ~n258 & n1505 ) ;
  assign n1507 = n301 | n1451 ;
  assign n1508 = ( ~n177 & n396 ) | ( ~n177 & n1219 ) | ( n396 & n1219 ) ;
  assign n1509 = n188 | n1464 ;
  assign n1510 = n237 | n1461 ;
  assign n1511 = n170 | n992 ;
  assign n1512 = ( ~n178 & n182 ) | ( ~n178 & n1485 ) | ( n182 & n1485 ) ;
  assign n1513 = ( ~n177 & n393 ) | ( ~n177 & n1070 ) | ( n393 & n1070 ) ;
  assign n1514 = n213 | n231 ;
  assign n1515 = ( ~n312 & n396 ) | ( ~n312 & n1507 ) | ( n396 & n1507 ) ;
  assign n1516 = ( n190 & ~n399 ) | ( n190 & n1511 ) | ( ~n399 & n1511 ) ;
  assign n1517 = n177 | n1508 ;
  assign n1518 = ( n238 & ~n411 ) | ( n238 & n1509 ) | ( ~n411 & n1509 ) ;
  assign n1519 = n312 | n1515 ;
  assign n1520 = ( n348 & ~n450 ) | ( n348 & n1519 ) | ( ~n450 & n1519 ) ;
  assign n1521 = ( n231 & ~n450 ) | ( n231 & n1520 ) | ( ~n450 & n1520 ) ;
  assign n1522 = n237 | n399 ;
  assign n1523 = n178 | n1512 ;
  assign n1524 = ( ~n348 & n1015 ) | ( ~n348 & n1523 ) | ( n1015 & n1523 ) ;
  assign n1525 = ( n160 & n937 ) | ( n160 & ~n1522 ) | ( n937 & ~n1522 ) ;
  assign n1526 = n450 | n1521 ;
  assign n1527 = n1522 | n1525 ;
  assign n1528 = ( n808 & n1470 ) | ( n808 & ~n1527 ) | ( n1470 & ~n1527 ) ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = n224 | n1180 ;
  assign n1531 = ( ~n411 & n1514 ) | ( ~n411 & n1527 ) | ( n1514 & n1527 ) ;
  assign n1532 = n411 | n1531 ;
  assign n1533 = ( n1227 & n1452 ) | ( n1227 & ~n1532 ) | ( n1452 & ~n1532 ) ;
  assign n1534 = n1532 | n1533 ;
  assign n1535 = ( n178 & ~n634 ) | ( n178 & n1534 ) | ( ~n634 & n1534 ) ;
  assign n1536 = n634 | n1535 ;
  assign n1537 = ( ~n139 & n170 ) | ( ~n139 & n1536 ) | ( n170 & n1536 ) ;
  assign n1538 = n139 | n1537 ;
  assign n1539 = ( ~n181 & n224 ) | ( ~n181 & n1538 ) | ( n224 & n1538 ) ;
  assign n1540 = n399 | n1516 ;
  assign n1541 = n181 | n1539 ;
  assign n1542 = n411 | n1518 ;
  assign n1543 = ( ~n177 & n396 ) | ( ~n177 & n1133 ) | ( n396 & n1133 ) ;
  assign n1544 = ( n126 & ~n389 ) | ( n126 & n1542 ) | ( ~n389 & n1542 ) ;
  assign n1545 = ( ~n146 & n190 ) | ( ~n146 & n1517 ) | ( n190 & n1517 ) ;
  assign n1546 = n146 | n1545 ;
  assign n1547 = n450 | n1410 ;
  assign n1548 = n178 | n1489 ;
  assign n1549 = ~n396 & n1543 ;
  assign n1550 = ( n343 & ~n460 ) | ( n343 & n1546 ) | ( ~n460 & n1546 ) ;
  assign n1551 = ( ~n428 & n460 ) | ( ~n428 & n1550 ) | ( n460 & n1550 ) ;
  assign n1552 = n177 | n1513 ;
  assign n1553 = ( ~n880 & n1310 ) | ( ~n880 & n1532 ) | ( n1310 & n1532 ) ;
  assign n1554 = n299 | n1407 ;
  assign n1555 = n299 | n1532 ;
  assign n1556 = n122 | n1555 ;
  assign n1557 = n299 | n1243 ;
  assign n1558 = n222 | n392 ;
  assign n1559 = ( ~n880 & n1119 ) | ( ~n880 & n1556 ) | ( n1119 & n1556 ) ;
  assign n1560 = n1192 | n1547 ;
  assign n1561 = n1282 | n1547 ;
  assign n1562 = ( n276 & ~n785 ) | ( n276 & n1561 ) | ( ~n785 & n1561 ) ;
  assign n1563 = n785 | n1562 ;
  assign n1564 = n159 | n1183 ;
  assign n1565 = ( ~n160 & n325 ) | ( ~n160 & n1564 ) | ( n325 & n1564 ) ;
  assign n1566 = ( n160 & ~n419 ) | ( n160 & n1565 ) | ( ~n419 & n1565 ) ;
  assign n1567 = n261 | n325 ;
  assign n1568 = n880 | n1553 ;
  assign n1569 = n235 | n426 ;
  assign n1570 = ( n880 & ~n1558 ) | ( n880 & n1567 ) | ( ~n1558 & n1567 ) ;
  assign n1571 = n1558 | n1570 ;
  assign n1572 = ( n325 & ~n428 ) | ( n325 & n1444 ) | ( ~n428 & n1444 ) ;
  assign n1573 = ( ~n1560 & n1569 ) | ( ~n1560 & n1571 ) | ( n1569 & n1571 ) ;
  assign n1574 = n1560 | n1573 ;
  assign n1575 = n880 | n1559 ;
  assign n1576 = n1556 | n1571 ;
  assign n1577 = ( ~n1282 & n1325 ) | ( ~n1282 & n1575 ) | ( n1325 & n1575 ) ;
  assign n1578 = n1282 | n1577 ;
  assign n1579 = ( ~n182 & n343 ) | ( ~n182 & n1578 ) | ( n343 & n1578 ) ;
  assign n1580 = ( ~n137 & n343 ) | ( ~n137 & n1252 ) | ( n343 & n1252 ) ;
  assign n1581 = ( n989 & ~n1050 ) | ( n989 & n1568 ) | ( ~n1050 & n1568 ) ;
  assign n1582 = ( ~n312 & n1050 ) | ( ~n312 & n1581 ) | ( n1050 & n1581 ) ;
  assign n1583 = ( n137 & ~n392 ) | ( n137 & n1580 ) | ( ~n392 & n1580 ) ;
  assign n1584 = n312 | n1582 ;
  assign n1585 = ( ~n188 & n1050 ) | ( ~n188 & n1529 ) | ( n1050 & n1529 ) ;
  assign n1586 = n182 | n1579 ;
  assign n1587 = n392 | n1583 ;
  assign n1588 = n133 | n799 ;
  assign n1589 = ( ~n389 & n426 ) | ( ~n389 & n1588 ) | ( n426 & n1588 ) ;
  assign n1590 = ( n995 & ~n1409 ) | ( n995 & n1576 ) | ( ~n1409 & n1576 ) ;
  assign n1591 = ( ~n389 & n393 ) | ( ~n389 & n1477 ) | ( n393 & n1477 ) ;
  assign n1592 = ( n261 & ~n389 ) | ( n261 & n1544 ) | ( ~n389 & n1544 ) ;
  assign n1593 = ~n393 & n1591 ;
  assign n1594 = ( n320 & ~n426 ) | ( n320 & n1593 ) | ( ~n426 & n1593 ) ;
  assign n1595 = ~n320 & n1594 ;
  assign n1596 = ~n182 & n1459 ;
  assign n1597 = ( n133 & ~n394 ) | ( n133 & n1031 ) | ( ~n394 & n1031 ) ;
  assign n1598 = n133 | n954 ;
  assign n1599 = n419 | n1453 ;
  assign n1600 = ~n238 & n1353 ;
  assign n1601 = n394 | n1235 ;
  assign n1602 = ~n133 & n1456 ;
  assign n1603 = ( ~n348 & n428 ) | ( ~n348 & n1524 ) | ( n428 & n1524 ) ;
  assign n1604 = n348 | n1603 ;
  assign n1605 = n389 | n1592 ;
  assign n1606 = n428 | n1551 ;
  assign n1607 = ( n188 & ~n389 ) | ( n188 & n1466 ) | ( ~n389 & n1466 ) ;
  assign n1608 = n389 | n1607 ;
  assign n1609 = n419 | n1566 ;
  assign n1610 = n389 | n1589 ;
  assign n1611 = ( ~n159 & n478 ) | ( ~n159 & n1468 ) | ( n478 & n1468 ) ;
  assign n1612 = ~n478 & n1611 ;
  assign n1613 = ( ~n217 & n238 ) | ( ~n217 & n1612 ) | ( n238 & n1612 ) ;
  assign n1614 = n394 | n1597 ;
  assign n1615 = ( n238 & ~n419 ) | ( n238 & n1613 ) | ( ~n419 & n1613 ) ;
  assign n1616 = ~n238 & n1615 ;
  assign n1617 = n428 | n1423 ;
  assign n1618 = ( n222 & ~n394 ) | ( n222 & n1479 ) | ( ~n394 & n1479 ) ;
  assign n1619 = ( ~n137 & n222 ) | ( ~n137 & n1618 ) | ( n222 & n1618 ) ;
  assign n1620 = ~n222 & n1619 ;
  assign n1621 = ( ~n348 & n478 ) | ( ~n348 & n1182 ) | ( n478 & n1182 ) ;
  assign n1622 = n348 | n1621 ;
  assign n1623 = ( ~n258 & n303 ) | ( ~n258 & n1622 ) | ( n303 & n1622 ) ;
  assign n1624 = ( n137 & ~n258 ) | ( n137 & n1623 ) | ( ~n258 & n1623 ) ;
  assign n1625 = n258 | n1624 ;
  assign n1626 = n419 | n1498 ;
  assign n1627 = n428 | n1572 ;
  assign n1628 = n188 | n1585 ;
  assign n1629 = ( ~n188 & n258 ) | ( ~n188 & n1245 ) | ( n258 & n1245 ) ;
  assign n1630 = n188 | n1629 ;
  assign n1631 = n258 | n1506 ;
  assign n1632 = n159 | n1448 ;
  assign n1633 = ( n217 & ~n389 ) | ( n217 & n1541 ) | ( ~n389 & n1541 ) ;
  assign n1634 = n389 | n1633 ;
  assign n1635 = ~x22 & n30 ;
  assign n1636 = n1635 ^ x5 ^ 1'b0 ;
  assign n1637 = n1602 ^ n1596 ^ 1'b0 ;
  assign n1638 = n1596 & n1602 ;
  assign n1639 = n1600 & ~n1638 ;
  assign n1640 = n1602 | n1636 ;
  assign n1641 = ( n70 & ~n436 ) | ( n70 & n1602 ) | ( ~n436 & n1602 ) ;
  assign n1642 = n436 & n1636 ;
  assign n1643 = n1637 | n1639 ;
  assign n1644 = n1642 ^ n1636 ^ n1602 ;
  assign n1645 = n1602 ^ n52 ^ 1'b0 ;
  assign n1646 = n84 & n1637 ;
  assign n1647 = n1643 ^ n1638 ^ n1600 ;
  assign n1648 = ~n1646 & n1647 ;
  assign n1649 = n1640 ^ n436 ^ 1'b0 ;
  assign n1650 = ( n1640 & n1645 ) | ( n1640 & ~n1649 ) | ( n1645 & ~n1649 ) ;
  assign n1651 = n1650 ^ n1648 ^ 1'b0 ;
  assign n1652 = ( n84 & ~n1602 ) | ( n84 & n1641 ) | ( ~n1602 & n1641 ) ;
  assign n1653 = n1602 | n1652 ;
  assign n1654 = n82 ^ x14 ^ 1'b0 ;
  assign n1655 = ~n70 & n436 ;
  assign n1656 = n1637 | n1647 ;
  assign n1657 = ( n436 & n1644 ) | ( n436 & ~n1655 ) | ( n1644 & ~n1655 ) ;
  assign n1658 = ( ~n1646 & n1653 ) | ( ~n1646 & n1657 ) | ( n1653 & n1657 ) ;
  assign n1659 = n1648 & ~n1650 ;
  assign n1660 = n1651 & n1658 ;
  assign n1661 = ( n84 & ~n1643 ) | ( n84 & n1660 ) | ( ~n1643 & n1660 ) ;
  assign n1662 = ( n84 & n1656 ) | ( n84 & ~n1660 ) | ( n1656 & ~n1660 ) ;
  assign n1663 = ~n1661 & n1662 ;
  assign n1664 = n1637 & ~n1639 ;
  assign n1665 = ( n70 & ~n1663 ) | ( n70 & n1664 ) | ( ~n1663 & n1664 ) ;
  assign n1666 = n1637 & ~n1647 ;
  assign n1667 = ( n70 & n1663 ) | ( n70 & ~n1666 ) | ( n1663 & ~n1666 ) ;
  assign n1668 = ~n1637 & n1654 ;
  assign n1669 = ~n1665 & n1667 ;
  assign n1670 = ( n1651 & n1658 ) | ( n1651 & ~n1669 ) | ( n1658 & ~n1669 ) ;
  assign n1671 = ( n1643 & n1645 ) | ( n1643 & n1656 ) | ( n1645 & n1656 ) ;
  assign n1672 = n1668 ^ n1647 ^ 1'b0 ;
  assign n1673 = n1643 ^ n70 ^ 1'b0 ;
  assign n1674 = ( n1643 & n1656 ) | ( n1643 & ~n1673 ) | ( n1656 & ~n1673 ) ;
  assign n1675 = ( n1639 & n1647 ) | ( n1639 & n1672 ) | ( n1647 & n1672 ) ;
  assign n1676 = n44 & ~n1664 ;
  assign n1677 = ( n1636 & ~n1666 ) | ( n1636 & n1674 ) | ( ~n1666 & n1674 ) ;
  assign n1678 = ~x22 & n33 ;
  assign n1679 = ( n1636 & n1664 ) | ( n1636 & ~n1674 ) | ( n1664 & ~n1674 ) ;
  assign n1680 = n1677 & ~n1679 ;
  assign n1681 = n44 | n1666 ;
  assign n1682 = ~n1669 & n1670 ;
  assign n1683 = ( n1671 & n1676 ) | ( n1671 & ~n1681 ) | ( n1676 & ~n1681 ) ;
  assign n1684 = n52 | n1602 ;
  assign n1685 = n1684 ^ n436 ^ 1'b0 ;
  assign n1686 = n1602 ^ n44 ^ 1'b0 ;
  assign n1687 = ( n1684 & ~n1685 ) | ( n1684 & n1686 ) | ( ~n1685 & n1686 ) ;
  assign n1688 = n1687 ^ n1680 ^ n1659 ;
  assign n1689 = ( n1659 & n1680 ) | ( n1659 & ~n1687 ) | ( n1680 & ~n1687 ) ;
  assign n1690 = ( n1643 & n1656 ) | ( n1643 & n1686 ) | ( n1656 & n1686 ) ;
  assign n1691 = n1601 ^ n1600 ^ 1'b0 ;
  assign n1692 = n84 & ~n1691 ;
  assign n1693 = ( n1682 & n1688 ) | ( n1682 & ~n1692 ) | ( n1688 & ~n1692 ) ;
  assign n1694 = n1555 | n1563 ;
  assign n1695 = n1678 ^ x8 ^ 1'b0 ;
  assign n1696 = ~n1599 & n1601 ;
  assign n1697 = ( n1599 & n1600 ) | ( n1599 & ~n1696 ) | ( n1600 & ~n1696 ) ;
  assign n1698 = ~n1691 & n1697 ;
  assign n1699 = n1691 & n1697 ;
  assign n1700 = n1699 ^ n84 ^ 1'b0 ;
  assign n1701 = ( n1599 & n1600 ) | ( n1599 & n1698 ) | ( n1600 & n1698 ) ;
  assign n1702 = ( n84 & ~n1600 ) | ( n84 & n1601 ) | ( ~n1600 & n1601 ) ;
  assign n1703 = n1599 & ~n1702 ;
  assign n1704 = n1695 ^ n1602 ^ 1'b0 ;
  assign n1705 = n1691 | n1701 ;
  assign n1706 = n1691 & ~n1701 ;
  assign n1707 = n44 | n1602 ;
  assign n1708 = n1707 ^ n436 ^ 1'b0 ;
  assign n1709 = ( n1704 & n1707 ) | ( n1704 & ~n1708 ) | ( n1707 & ~n1708 ) ;
  assign n1710 = n1709 ^ n1703 ^ 1'b0 ;
  assign n1711 = ( n1599 & n1601 ) | ( n1599 & n1654 ) | ( n1601 & n1654 ) ;
  assign n1712 = ( n1699 & ~n1700 ) | ( n1699 & n1706 ) | ( ~n1700 & n1706 ) ;
  assign n1713 = ( n70 & n1705 ) | ( n70 & ~n1712 ) | ( n1705 & ~n1712 ) ;
  assign n1714 = ( n70 & n1698 ) | ( n70 & n1712 ) | ( n1698 & n1712 ) ;
  assign n1715 = n1713 & ~n1714 ;
  assign n1716 = n1666 | n1695 ;
  assign n1717 = ~n1691 & n1711 ;
  assign n1718 = n1717 ^ n1711 ^ n1599 ;
  assign n1719 = ~n1664 & n1695 ;
  assign n1720 = ( n1690 & ~n1716 ) | ( n1690 & n1719 ) | ( ~n1716 & n1719 ) ;
  assign n1721 = n1643 ^ n1636 ^ 1'b0 ;
  assign n1722 = ( n1643 & n1656 ) | ( n1643 & ~n1721 ) | ( n1656 & ~n1721 ) ;
  assign n1723 = ( n52 & n1664 ) | ( n52 & ~n1722 ) | ( n1664 & ~n1722 ) ;
  assign n1724 = ( n52 & ~n1666 ) | ( n52 & n1722 ) | ( ~n1666 & n1722 ) ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = n1725 ^ n1715 ^ n1710 ;
  assign n1727 = ( ~n1689 & n1693 ) | ( ~n1689 & n1726 ) | ( n1693 & n1726 ) ;
  assign n1728 = ( ~n84 & n684 ) | ( ~n84 & n1599 ) | ( n684 & n1599 ) ;
  assign n1729 = n684 | n1599 ;
  assign n1730 = n1599 ^ n684 ^ 1'b0 ;
  assign n1731 = ( ~n1710 & n1715 ) | ( ~n1710 & n1725 ) | ( n1715 & n1725 ) ;
  assign n1732 = ( n1598 & ~n1728 ) | ( n1598 & n1730 ) | ( ~n1728 & n1730 ) ;
  assign n1733 = n1732 ^ n1729 ^ n1728 ;
  assign n1734 = n1732 & ~n1733 ;
  assign n1735 = n1703 & ~n1709 ;
  assign n1736 = n1735 ^ n1734 ^ n1731 ;
  assign n1737 = ( n1731 & n1734 ) | ( n1731 & n1735 ) | ( n1734 & n1735 ) ;
  assign n1738 = n1699 ^ n70 ^ 1'b0 ;
  assign n1739 = n1602 | n1695 ;
  assign n1740 = n1739 ^ n436 ^ 1'b0 ;
  assign n1741 = n1602 ^ n79 ^ 1'b0 ;
  assign n1742 = ( n1699 & n1706 ) | ( n1699 & ~n1738 ) | ( n1706 & ~n1738 ) ;
  assign n1743 = ( n1739 & ~n1740 ) | ( n1739 & n1741 ) | ( ~n1740 & n1741 ) ;
  assign n1744 = ( n1636 & n1698 ) | ( n1636 & n1742 ) | ( n1698 & n1742 ) ;
  assign n1745 = ( n1643 & n1656 ) | ( n1643 & n1741 ) | ( n1656 & n1741 ) ;
  assign n1746 = ( n1636 & n1705 ) | ( n1636 & ~n1742 ) | ( n1705 & ~n1742 ) ;
  assign n1747 = ( n1643 & n1656 ) | ( n1643 & n1704 ) | ( n1656 & n1704 ) ;
  assign n1748 = ~n1744 & n1746 ;
  assign n1749 = n1748 ^ n1743 ^ n1683 ;
  assign n1750 = ( n1727 & ~n1736 ) | ( n1727 & n1749 ) | ( ~n1736 & n1749 ) ;
  assign n1751 = n38 | n1666 ;
  assign n1752 = ( n1683 & ~n1743 ) | ( n1683 & n1748 ) | ( ~n1743 & n1748 ) ;
  assign n1753 = n79 & ~n1664 ;
  assign n1754 = n79 | n1666 ;
  assign n1755 = n38 & ~n1664 ;
  assign n1756 = ( n1747 & n1753 ) | ( n1747 & ~n1754 ) | ( n1753 & ~n1754 ) ;
  assign n1757 = ( n1745 & ~n1751 ) | ( n1745 & n1755 ) | ( ~n1751 & n1755 ) ;
  assign n1758 = n1699 ^ n1636 ^ 1'b0 ;
  assign n1759 = ~n1598 & n1729 ;
  assign n1760 = n1730 | n1759 ;
  assign n1761 = n1760 ^ n1729 ^ n1598 ;
  assign n1762 = n1730 | n1761 ;
  assign n1763 = n1760 ^ n84 ^ 1'b0 ;
  assign n1764 = n1602 ^ n38 ^ 1'b0 ;
  assign n1765 = n1730 & ~n1759 ;
  assign n1766 = ( n1699 & n1706 ) | ( n1699 & ~n1758 ) | ( n1706 & ~n1758 ) ;
  assign n1767 = n79 | n1602 ;
  assign n1768 = ( n52 & n1705 ) | ( n52 & ~n1766 ) | ( n1705 & ~n1766 ) ;
  assign n1769 = ( n52 & n1698 ) | ( n52 & n1766 ) | ( n1698 & n1766 ) ;
  assign n1770 = n1767 ^ n436 ^ 1'b0 ;
  assign n1771 = ( n1760 & n1762 ) | ( n1760 & ~n1763 ) | ( n1762 & ~n1763 ) ;
  assign n1772 = n1730 & ~n1761 ;
  assign n1773 = n1768 & ~n1769 ;
  assign n1774 = ( n70 & n1765 ) | ( n70 & ~n1771 ) | ( n1765 & ~n1771 ) ;
  assign n1775 = ( n1764 & n1767 ) | ( n1764 & ~n1770 ) | ( n1767 & ~n1770 ) ;
  assign n1776 = n40 ^ x11 ^ 1'b0 ;
  assign n1777 = ( n70 & n1771 ) | ( n70 & ~n1772 ) | ( n1771 & ~n1772 ) ;
  assign n1778 = ~n1774 & n1777 ;
  assign n1779 = ( n1643 & n1656 ) | ( n1643 & n1764 ) | ( n1656 & n1764 ) ;
  assign n1780 = ( n1720 & n1773 ) | ( n1720 & n1778 ) | ( n1773 & n1778 ) ;
  assign n1781 = n1778 ^ n1773 ^ n1720 ;
  assign n1782 = n1775 ^ n1733 ^ 1'b0 ;
  assign n1783 = n1782 ^ n1781 ^ n1752 ;
  assign n1784 = ( ~n1737 & n1750 ) | ( ~n1737 & n1783 ) | ( n1750 & n1783 ) ;
  assign n1785 = n75 & ~n1664 ;
  assign n1786 = n1666 | n1776 ;
  assign n1787 = ( n1654 & n1730 ) | ( n1654 & n1759 ) | ( n1730 & n1759 ) ;
  assign n1788 = ~n1664 & n1776 ;
  assign n1789 = ( n1779 & ~n1786 ) | ( n1779 & n1788 ) | ( ~n1786 & n1788 ) ;
  assign n1790 = n1733 & ~n1775 ;
  assign n1791 = n1776 ^ n1602 ^ 1'b0 ;
  assign n1792 = ( n1643 & n1656 ) | ( n1643 & n1791 ) | ( n1656 & n1791 ) ;
  assign n1793 = ( n1752 & n1781 ) | ( n1752 & ~n1782 ) | ( n1781 & ~n1782 ) ;
  assign n1794 = n75 | n1666 ;
  assign n1795 = ( n1785 & n1792 ) | ( n1785 & ~n1794 ) | ( n1792 & ~n1794 ) ;
  assign n1796 = n38 | n1602 ;
  assign n1797 = n1796 ^ n436 ^ 1'b0 ;
  assign n1798 = ( n1791 & n1796 ) | ( n1791 & ~n1797 ) | ( n1796 & ~n1797 ) ;
  assign n1799 = n1602 ^ n75 ^ 1'b0 ;
  assign n1800 = ( n1643 & n1656 ) | ( n1643 & n1799 ) | ( n1656 & n1799 ) ;
  assign n1801 = n56 | n1666 ;
  assign n1802 = n56 & ~n1664 ;
  assign n1803 = ( n1800 & ~n1801 ) | ( n1800 & n1802 ) | ( ~n1801 & n1802 ) ;
  assign n1804 = n1602 ^ n56 ^ 1'b0 ;
  assign n1805 = ( n1643 & n1656 ) | ( n1643 & n1804 ) | ( n1656 & n1804 ) ;
  assign n1806 = n1602 | n1776 ;
  assign n1807 = n1654 | n1666 ;
  assign n1808 = n1654 & ~n1664 ;
  assign n1809 = ( n1805 & ~n1807 ) | ( n1805 & n1808 ) | ( ~n1807 & n1808 ) ;
  assign n1810 = n1699 ^ n52 ^ 1'b0 ;
  assign n1811 = ( n1699 & n1706 ) | ( n1699 & ~n1810 ) | ( n1706 & ~n1810 ) ;
  assign n1812 = ( n44 & n1698 ) | ( n44 & n1811 ) | ( n1698 & n1811 ) ;
  assign n1813 = ( n44 & n1705 ) | ( n44 & ~n1811 ) | ( n1705 & ~n1811 ) ;
  assign n1814 = n1806 ^ n436 ^ 1'b0 ;
  assign n1815 = ( n1799 & n1806 ) | ( n1799 & ~n1814 ) | ( n1806 & ~n1814 ) ;
  assign n1816 = n1614 ^ n1598 ^ 1'b0 ;
  assign n1817 = ~n1812 & n1813 ;
  assign n1818 = n84 & n1816 ;
  assign n1819 = n1817 ^ n1798 ^ n1756 ;
  assign n1820 = ( n1756 & ~n1798 ) | ( n1756 & n1817 ) | ( ~n1798 & n1817 ) ;
  assign n1821 = n1760 ^ n70 ^ 1'b0 ;
  assign n1822 = ( n1760 & n1762 ) | ( n1760 & ~n1821 ) | ( n1762 & ~n1821 ) ;
  assign n1823 = ( n1636 & ~n1772 ) | ( n1636 & n1822 ) | ( ~n1772 & n1822 ) ;
  assign n1824 = ( n1636 & n1765 ) | ( n1636 & ~n1822 ) | ( n1765 & ~n1822 ) ;
  assign n1825 = n1823 & ~n1824 ;
  assign n1826 = ( n1790 & n1818 ) | ( n1790 & n1825 ) | ( n1818 & n1825 ) ;
  assign n1827 = n1825 ^ n1818 ^ n1790 ;
  assign n1828 = n1827 ^ n1819 ^ n1780 ;
  assign n1829 = ( n1780 & ~n1819 ) | ( n1780 & n1827 ) | ( ~n1819 & n1827 ) ;
  assign n1830 = ( n1784 & ~n1793 ) | ( n1784 & n1828 ) | ( ~n1793 & n1828 ) ;
  assign n1831 = n1598 | n1614 ;
  assign n1832 = n1699 ^ n44 ^ 1'b0 ;
  assign n1833 = ( n1699 & n1706 ) | ( n1699 & ~n1832 ) | ( n1706 & ~n1832 ) ;
  assign n1834 = ~n1574 & n1831 ;
  assign n1835 = ( n1695 & n1705 ) | ( n1695 & ~n1833 ) | ( n1705 & ~n1833 ) ;
  assign n1836 = n1760 ^ n1636 ^ 1'b0 ;
  assign n1837 = ( n1760 & n1762 ) | ( n1760 & ~n1836 ) | ( n1762 & ~n1836 ) ;
  assign n1838 = n1816 | n1834 ;
  assign n1839 = ( n52 & n1765 ) | ( n52 & ~n1837 ) | ( n1765 & ~n1837 ) ;
  assign n1840 = ( n1695 & n1698 ) | ( n1695 & n1833 ) | ( n1698 & n1833 ) ;
  assign n1841 = ( n52 & ~n1772 ) | ( n52 & n1837 ) | ( ~n1772 & n1837 ) ;
  assign n1842 = n1835 & ~n1840 ;
  assign n1843 = ( n84 & n1598 ) | ( n84 & n1614 ) | ( n1598 & n1614 ) ;
  assign n1844 = n1574 & ~n1843 ;
  assign n1845 = n75 | n1602 ;
  assign n1846 = n1838 ^ n1831 ^ n1574 ;
  assign n1847 = n1845 ^ n436 ^ 1'b0 ;
  assign n1848 = ( n1804 & n1845 ) | ( n1804 & ~n1847 ) | ( n1845 & ~n1847 ) ;
  assign n1849 = ~n1815 & n1844 ;
  assign n1850 = n1816 & ~n1846 ;
  assign n1851 = n1844 ^ n1815 ^ 1'b0 ;
  assign n1852 = n1574 | n1694 ;
  assign n1853 = n1694 ^ n1574 ^ 1'b0 ;
  assign n1854 = ( n1654 & n1816 ) | ( n1654 & n1834 ) | ( n1816 & n1834 ) ;
  assign n1855 = ~n1839 & n1841 ;
  assign n1856 = ( n1757 & n1842 ) | ( n1757 & n1855 ) | ( n1842 & n1855 ) ;
  assign n1857 = n1855 ^ n1842 ^ n1757 ;
  assign n1858 = n1816 | n1846 ;
  assign n1859 = n1838 ^ n84 ^ 1'b0 ;
  assign n1860 = n1816 & ~n1834 ;
  assign n1861 = ( n1838 & n1858 ) | ( n1838 & ~n1859 ) | ( n1858 & ~n1859 ) ;
  assign n1862 = ( n70 & ~n1850 ) | ( n70 & n1861 ) | ( ~n1850 & n1861 ) ;
  assign n1863 = ( n70 & n1860 ) | ( n70 & ~n1861 ) | ( n1860 & ~n1861 ) ;
  assign n1864 = n1862 & ~n1863 ;
  assign n1865 = ( n1820 & ~n1851 ) | ( n1820 & n1864 ) | ( ~n1851 & n1864 ) ;
  assign n1866 = n1864 ^ n1851 ^ n1820 ;
  assign n1867 = n1866 ^ n1857 ^ n1826 ;
  assign n1868 = ( ~n1829 & n1830 ) | ( ~n1829 & n1867 ) | ( n1830 & n1867 ) ;
  assign n1869 = n1760 ^ n52 ^ 1'b0 ;
  assign n1870 = n1699 ^ n1695 ^ 1'b0 ;
  assign n1871 = ( ~n84 & n1409 ) | ( ~n84 & n1853 ) | ( n1409 & n1853 ) ;
  assign n1872 = ( n1826 & n1857 ) | ( n1826 & ~n1866 ) | ( n1857 & ~n1866 ) ;
  assign n1873 = ( n1699 & n1706 ) | ( n1699 & ~n1870 ) | ( n1706 & ~n1870 ) ;
  assign n1874 = ( n79 & n1705 ) | ( n79 & ~n1873 ) | ( n1705 & ~n1873 ) ;
  assign n1875 = ( n79 & n1698 ) | ( n79 & n1873 ) | ( n1698 & n1873 ) ;
  assign n1876 = n1874 & ~n1875 ;
  assign n1877 = ( n1760 & n1762 ) | ( n1760 & ~n1869 ) | ( n1762 & ~n1869 ) ;
  assign n1878 = n1853 & ~n1871 ;
  assign n1879 = ( n44 & n1765 ) | ( n44 & ~n1877 ) | ( n1765 & ~n1877 ) ;
  assign n1880 = ( n44 & ~n1772 ) | ( n44 & n1877 ) | ( ~n1772 & n1877 ) ;
  assign n1881 = ~n1879 & n1880 ;
  assign n1882 = n1881 ^ n1876 ^ n1849 ;
  assign n1883 = ( n1856 & n1878 ) | ( n1856 & n1882 ) | ( n1878 & n1882 ) ;
  assign n1884 = n1882 ^ n1878 ^ n1856 ;
  assign n1885 = n1838 ^ n70 ^ 1'b0 ;
  assign n1886 = ( n1838 & n1858 ) | ( n1838 & ~n1885 ) | ( n1858 & ~n1885 ) ;
  assign n1887 = ( n1636 & ~n1850 ) | ( n1636 & n1886 ) | ( ~n1850 & n1886 ) ;
  assign n1888 = ( n1636 & n1860 ) | ( n1636 & ~n1886 ) | ( n1860 & ~n1886 ) ;
  assign n1889 = n1887 & ~n1888 ;
  assign n1890 = ( n1789 & ~n1848 ) | ( n1789 & n1889 ) | ( ~n1848 & n1889 ) ;
  assign n1891 = ( n1849 & n1876 ) | ( n1849 & n1881 ) | ( n1876 & n1881 ) ;
  assign n1892 = n1889 ^ n1848 ^ n1789 ;
  assign n1893 = ( n1865 & n1884 ) | ( n1865 & ~n1892 ) | ( n1884 & ~n1892 ) ;
  assign n1894 = n1892 ^ n1884 ^ n1865 ;
  assign n1895 = ( n1868 & ~n1872 ) | ( n1868 & n1894 ) | ( ~n1872 & n1894 ) ;
  assign n1896 = n1838 ^ n1636 ^ 1'b0 ;
  assign n1897 = ( n1838 & n1858 ) | ( n1838 & ~n1896 ) | ( n1858 & ~n1896 ) ;
  assign n1898 = ( n52 & n1860 ) | ( n52 & ~n1897 ) | ( n1860 & ~n1897 ) ;
  assign n1899 = ( n52 & ~n1850 ) | ( n52 & n1897 ) | ( ~n1850 & n1897 ) ;
  assign n1900 = n1699 ^ n79 ^ 1'b0 ;
  assign n1901 = ( n1699 & n1706 ) | ( n1699 & ~n1900 ) | ( n1706 & ~n1900 ) ;
  assign n1902 = ( n38 & n1698 ) | ( n38 & n1901 ) | ( n1698 & n1901 ) ;
  assign n1903 = ( n38 & n1705 ) | ( n38 & ~n1901 ) | ( n1705 & ~n1901 ) ;
  assign n1904 = ~n1902 & n1903 ;
  assign n1905 = n436 & ~n1654 ;
  assign n1906 = ( n436 & n1602 ) | ( n436 & ~n1905 ) | ( n1602 & ~n1905 ) ;
  assign n1907 = n1760 ^ n44 ^ 1'b0 ;
  assign n1908 = ~n1898 & n1899 ;
  assign n1909 = ( n1760 & n1762 ) | ( n1760 & ~n1907 ) | ( n1762 & ~n1907 ) ;
  assign n1910 = ( n1695 & n1765 ) | ( n1695 & ~n1909 ) | ( n1765 & ~n1909 ) ;
  assign n1911 = ( n1695 & ~n1772 ) | ( n1695 & n1909 ) | ( ~n1772 & n1909 ) ;
  assign n1912 = ~n1910 & n1911 ;
  assign n1913 = n1912 ^ n1908 ^ n1904 ;
  assign n1914 = ( n1904 & n1908 ) | ( n1904 & n1912 ) | ( n1908 & n1912 ) ;
  assign n1915 = ( n1890 & n1891 ) | ( n1890 & n1913 ) | ( n1891 & n1913 ) ;
  assign n1916 = n1913 ^ n1891 ^ n1890 ;
  assign n1917 = n1852 ^ n84 ^ 1'b0 ;
  assign n1918 = n1409 | n1853 ;
  assign n1919 = n1654 ^ n1602 ^ 1'b0 ;
  assign n1920 = ( n1852 & ~n1917 ) | ( n1852 & n1918 ) | ( ~n1917 & n1918 ) ;
  assign n1921 = n70 & n1853 ;
  assign n1922 = ( ~n1853 & n1920 ) | ( ~n1853 & n1921 ) | ( n1920 & n1921 ) ;
  assign n1923 = n56 | n1602 ;
  assign n1924 = n1923 ^ n436 ^ 1'b0 ;
  assign n1925 = ( n1919 & n1923 ) | ( n1919 & ~n1924 ) | ( n1923 & ~n1924 ) ;
  assign n1926 = n1925 ^ n1409 ^ 1'b0 ;
  assign n1927 = n1926 ^ n1922 ^ n1795 ;
  assign n1928 = ( n1795 & n1922 ) | ( n1795 & ~n1926 ) | ( n1922 & ~n1926 ) ;
  assign n1929 = n1927 ^ n1916 ^ n1883 ;
  assign n1930 = ( ~n1893 & n1895 ) | ( ~n1893 & n1929 ) | ( n1895 & n1929 ) ;
  assign n1931 = ( n1883 & n1916 ) | ( n1883 & ~n1927 ) | ( n1916 & ~n1927 ) ;
  assign n1932 = ~n1636 & n1853 ;
  assign n1933 = ~n70 & n1918 ;
  assign n1934 = n1409 & ~n1925 ;
  assign n1935 = n70 & n1852 ;
  assign n1936 = ( ~n1932 & n1933 ) | ( ~n1932 & n1935 ) | ( n1933 & n1935 ) ;
  assign n1937 = ( n1914 & n1934 ) | ( n1914 & n1936 ) | ( n1934 & n1936 ) ;
  assign n1938 = n1936 ^ n1934 ^ n1914 ;
  assign n1939 = n1699 ^ n38 ^ 1'b0 ;
  assign n1940 = ( n1699 & n1706 ) | ( n1699 & ~n1939 ) | ( n1706 & ~n1939 ) ;
  assign n1941 = n1699 ^ n75 ^ 1'b0 ;
  assign n1942 = n84 & n1409 ;
  assign n1943 = ( n1699 & n1706 ) | ( n1699 & ~n1941 ) | ( n1706 & ~n1941 ) ;
  assign n1944 = n1942 ^ n1906 ^ n1803 ;
  assign n1945 = ( n1803 & ~n1906 ) | ( n1803 & n1942 ) | ( ~n1906 & n1942 ) ;
  assign n1946 = ( n1698 & n1776 ) | ( n1698 & n1940 ) | ( n1776 & n1940 ) ;
  assign n1947 = ( n1705 & n1776 ) | ( n1705 & ~n1940 ) | ( n1776 & ~n1940 ) ;
  assign n1948 = ~n1946 & n1947 ;
  assign n1949 = n1776 ^ n1699 ^ 1'b0 ;
  assign n1950 = ( n1699 & n1706 ) | ( n1699 & ~n1949 ) | ( n1706 & ~n1949 ) ;
  assign n1951 = n1699 ^ n56 ^ 1'b0 ;
  assign n1952 = ( n1699 & n1706 ) | ( n1699 & ~n1951 ) | ( n1706 & ~n1951 ) ;
  assign n1953 = ( n56 & n1698 ) | ( n56 & n1943 ) | ( n1698 & n1943 ) ;
  assign n1954 = ( n1654 & n1698 ) | ( n1654 & n1952 ) | ( n1698 & n1952 ) ;
  assign n1955 = ( n56 & n1705 ) | ( n56 & ~n1943 ) | ( n1705 & ~n1943 ) ;
  assign n1956 = ~n1953 & n1955 ;
  assign n1957 = n1838 ^ n52 ^ 1'b0 ;
  assign n1958 = ( n1654 & n1705 ) | ( n1654 & ~n1952 ) | ( n1705 & ~n1952 ) ;
  assign n1959 = ~n1954 & n1958 ;
  assign n1960 = ( n1838 & n1858 ) | ( n1838 & ~n1957 ) | ( n1858 & ~n1957 ) ;
  assign n1961 = ( n44 & n1860 ) | ( n44 & ~n1960 ) | ( n1860 & ~n1960 ) ;
  assign n1962 = ( n75 & n1705 ) | ( n75 & ~n1950 ) | ( n1705 & ~n1950 ) ;
  assign n1963 = ( n44 & ~n1850 ) | ( n44 & n1960 ) | ( ~n1850 & n1960 ) ;
  assign n1964 = ~n1961 & n1963 ;
  assign n1965 = n1760 ^ n1695 ^ 1'b0 ;
  assign n1966 = ( n1760 & n1762 ) | ( n1760 & ~n1965 ) | ( n1762 & ~n1965 ) ;
  assign n1967 = ( n75 & n1698 ) | ( n75 & n1950 ) | ( n1698 & n1950 ) ;
  assign n1968 = ( n79 & n1765 ) | ( n79 & ~n1966 ) | ( n1765 & ~n1966 ) ;
  assign n1969 = ( n79 & ~n1772 ) | ( n79 & n1966 ) | ( ~n1772 & n1966 ) ;
  assign n1970 = ~n1968 & n1969 ;
  assign n1971 = n1970 ^ n1964 ^ n1948 ;
  assign n1972 = ( n1948 & n1964 ) | ( n1948 & n1970 ) | ( n1964 & n1970 ) ;
  assign n1973 = n1971 ^ n1944 ^ n1928 ;
  assign n1974 = n1973 ^ n1938 ^ n1915 ;
  assign n1975 = n1962 & ~n1967 ;
  assign n1976 = n1974 ^ n1931 ^ n1930 ;
  assign n1977 = ( n1915 & n1938 ) | ( n1915 & ~n1973 ) | ( n1938 & ~n1973 ) ;
  assign n1978 = ( n1930 & ~n1931 ) | ( n1930 & n1974 ) | ( ~n1931 & n1974 ) ;
  assign n1979 = ( n1928 & ~n1944 ) | ( n1928 & n1971 ) | ( ~n1944 & n1971 ) ;
  assign n1980 = n1760 ^ n79 ^ 1'b0 ;
  assign n1981 = ( n1760 & n1762 ) | ( n1760 & ~n1980 ) | ( n1762 & ~n1980 ) ;
  assign n1982 = n52 & n1853 ;
  assign n1983 = n1852 ^ n1636 ^ 1'b0 ;
  assign n1984 = ( n1852 & n1918 ) | ( n1852 & ~n1983 ) | ( n1918 & ~n1983 ) ;
  assign n1985 = ( ~n1853 & n1982 ) | ( ~n1853 & n1984 ) | ( n1982 & n1984 ) ;
  assign n1986 = n1985 ^ n1972 ^ n1945 ;
  assign n1987 = ( n1945 & n1972 ) | ( n1945 & n1985 ) | ( n1972 & n1985 ) ;
  assign n1988 = n1838 ^ n44 ^ 1'b0 ;
  assign n1989 = ( n1838 & n1858 ) | ( n1838 & ~n1988 ) | ( n1858 & ~n1988 ) ;
  assign n1990 = ( n1695 & ~n1850 ) | ( n1695 & n1989 ) | ( ~n1850 & n1989 ) ;
  assign n1991 = ( n1695 & n1860 ) | ( n1695 & ~n1989 ) | ( n1860 & ~n1989 ) ;
  assign n1992 = n1990 & ~n1991 ;
  assign n1993 = ( n38 & n1765 ) | ( n38 & ~n1981 ) | ( n1765 & ~n1981 ) ;
  assign n1994 = ( n38 & ~n1772 ) | ( n38 & n1981 ) | ( ~n1772 & n1981 ) ;
  assign n1995 = ~n1993 & n1994 ;
  assign n1996 = ( n1975 & n1992 ) | ( n1975 & n1995 ) | ( n1992 & n1995 ) ;
  assign n1997 = n1995 ^ n1992 ^ n1975 ;
  assign n1998 = n70 & n1409 ;
  assign n1999 = ( ~n1602 & n1809 ) | ( ~n1602 & n1998 ) | ( n1809 & n1998 ) ;
  assign n2000 = n1998 ^ n1809 ^ n1602 ;
  assign n2001 = n2000 ^ n1997 ^ n1937 ;
  assign n2002 = ( n1937 & n1997 ) | ( n1937 & ~n2000 ) | ( n1997 & ~n2000 ) ;
  assign n2003 = n2001 ^ n1986 ^ n1979 ;
  assign n2004 = ( ~n1977 & n1978 ) | ( ~n1977 & n2003 ) | ( n1978 & n2003 ) ;
  assign n2005 = n2003 ^ n1978 ^ n1977 ;
  assign n2006 = n1838 ^ n1695 ^ 1'b0 ;
  assign n2007 = ( n1838 & n1858 ) | ( n1838 & ~n2006 ) | ( n1858 & ~n2006 ) ;
  assign n2008 = ( n79 & ~n1850 ) | ( n79 & n2007 ) | ( ~n1850 & n2007 ) ;
  assign n2009 = ( n1979 & n1986 ) | ( n1979 & ~n2001 ) | ( n1986 & ~n2001 ) ;
  assign n2010 = ( n79 & n1860 ) | ( n79 & ~n2007 ) | ( n1860 & ~n2007 ) ;
  assign n2011 = n2008 & ~n2010 ;
  assign n2012 = n1760 ^ n38 ^ 1'b0 ;
  assign n2013 = ( n1760 & n1762 ) | ( n1760 & ~n2012 ) | ( n1762 & ~n2012 ) ;
  assign n2014 = n1976 ^ n1247 ^ 1'b0 ;
  assign n2015 = ~n1247 & n1976 ;
  assign n2016 = ( ~n1772 & n1776 ) | ( ~n1772 & n2013 ) | ( n1776 & n2013 ) ;
  assign n2017 = ( n1765 & n1776 ) | ( n1765 & ~n2013 ) | ( n1776 & ~n2013 ) ;
  assign n2018 = n2015 ^ n2005 ^ n1606 ;
  assign n2019 = n2016 & ~n2017 ;
  assign n2020 = ( ~n1606 & n2005 ) | ( ~n1606 & n2015 ) | ( n2005 & n2015 ) ;
  assign n2021 = n1409 & n1636 ;
  assign n2022 = ( ~n1602 & n1675 ) | ( ~n1602 & n2021 ) | ( n1675 & n2021 ) ;
  assign n2023 = n52 & n1409 ;
  assign n2024 = n2021 ^ n1675 ^ n1602 ;
  assign n2025 = n2019 ^ n2011 ^ n1956 ;
  assign n2026 = ( n1956 & n2011 ) | ( n1956 & n2019 ) | ( n2011 & n2019 ) ;
  assign n2027 = ~n44 & n1853 ;
  assign n2028 = n2025 ^ n2024 ^ n1987 ;
  assign n2029 = ( n1987 & ~n2024 ) | ( n1987 & n2025 ) | ( ~n2024 & n2025 ) ;
  assign n2030 = ~n52 & n1918 ;
  assign n2031 = n52 & n1852 ;
  assign n2032 = ( ~n2027 & n2030 ) | ( ~n2027 & n2031 ) | ( n2030 & n2031 ) ;
  assign n2033 = ( n1602 & ~n1647 ) | ( n1602 & n2023 ) | ( ~n1647 & n2023 ) ;
  assign n2034 = n2032 ^ n1999 ^ n1996 ;
  assign n2035 = n2023 ^ n1647 ^ n1602 ;
  assign n2036 = n2034 ^ n2028 ^ n2002 ;
  assign n2037 = ( n2004 & ~n2009 ) | ( n2004 & n2036 ) | ( ~n2009 & n2036 ) ;
  assign n2038 = n2036 ^ n2009 ^ n2004 ;
  assign n2039 = n1776 ^ n1760 ^ 1'b0 ;
  assign n2040 = ( n1760 & n1762 ) | ( n1760 & ~n2039 ) | ( n1762 & ~n2039 ) ;
  assign n2041 = ( n1329 & n2020 ) | ( n1329 & n2038 ) | ( n2020 & n2038 ) ;
  assign n2042 = n2038 ^ n2020 ^ n1329 ;
  assign n2043 = ( n75 & n1765 ) | ( n75 & ~n2040 ) | ( n1765 & ~n2040 ) ;
  assign n2044 = ( n1996 & n1999 ) | ( n1996 & n2032 ) | ( n1999 & n2032 ) ;
  assign n2045 = ( n75 & ~n1772 ) | ( n75 & n2040 ) | ( ~n1772 & n2040 ) ;
  assign n2046 = ~n2043 & n2045 ;
  assign n2047 = ( n2022 & ~n2035 ) | ( n2022 & n2046 ) | ( ~n2035 & n2046 ) ;
  assign n2048 = ( n2002 & ~n2028 ) | ( n2002 & n2034 ) | ( ~n2028 & n2034 ) ;
  assign n2049 = n2046 ^ n2035 ^ n2022 ;
  assign n2050 = n1760 ^ n56 ^ 1'b0 ;
  assign n2051 = ( n1760 & n1762 ) | ( n1760 & ~n2050 ) | ( n1762 & ~n2050 ) ;
  assign n2052 = n1760 ^ n75 ^ 1'b0 ;
  assign n2053 = ( n1760 & n1762 ) | ( n1760 & ~n2052 ) | ( n1762 & ~n2052 ) ;
  assign n2054 = n1852 ^ n1695 ^ 1'b0 ;
  assign n2055 = n79 & n1853 ;
  assign n2056 = ( n1852 & n1918 ) | ( n1852 & ~n2054 ) | ( n1918 & ~n2054 ) ;
  assign n2057 = ( ~n1853 & n2055 ) | ( ~n1853 & n2056 ) | ( n2055 & n2056 ) ;
  assign n2058 = ( n1654 & n1765 ) | ( n1654 & ~n2051 ) | ( n1765 & ~n2051 ) ;
  assign n2059 = ( n1654 & ~n1772 ) | ( n1654 & n2051 ) | ( ~n1772 & n2051 ) ;
  assign n2060 = ( n56 & n1765 ) | ( n56 & ~n2053 ) | ( n1765 & ~n2053 ) ;
  assign n2061 = ~n2058 & n2059 ;
  assign n2062 = ~n1654 & n1846 ;
  assign n2063 = ( ~n1850 & n1854 ) | ( ~n1850 & n2062 ) | ( n1854 & n2062 ) ;
  assign n2064 = ( n56 & ~n1772 ) | ( n56 & n2053 ) | ( ~n1772 & n2053 ) ;
  assign n2065 = ~n2060 & n2064 ;
  assign n2066 = ~n1654 & n1761 ;
  assign n2067 = n44 & n1852 ;
  assign n2068 = ( ~n1772 & n1787 ) | ( ~n1772 & n2066 ) | ( n1787 & n2066 ) ;
  assign n2069 = ~n44 & n1918 ;
  assign n2070 = ~n1695 & n1853 ;
  assign n2071 = ( n2067 & n2069 ) | ( n2067 & ~n2070 ) | ( n2069 & ~n2070 ) ;
  assign n2072 = n1838 ^ n79 ^ 1'b0 ;
  assign n2073 = ( n1838 & n1858 ) | ( n1838 & ~n2072 ) | ( n1858 & ~n2072 ) ;
  assign n2074 = ( n38 & ~n1850 ) | ( n38 & n2073 ) | ( ~n1850 & n2073 ) ;
  assign n2075 = ( n38 & n1860 ) | ( n38 & ~n2073 ) | ( n1860 & ~n2073 ) ;
  assign n2076 = n2074 & ~n2075 ;
  assign n2077 = ( n1959 & n2071 ) | ( n1959 & n2076 ) | ( n2071 & n2076 ) ;
  assign n2078 = n2076 ^ n2071 ^ n1959 ;
  assign n2079 = n1838 ^ n75 ^ 1'b0 ;
  assign n2080 = ( n2026 & n2044 ) | ( n2026 & n2078 ) | ( n2044 & n2078 ) ;
  assign n2081 = n2078 ^ n2044 ^ n2026 ;
  assign n2082 = ( n1838 & n1858 ) | ( n1838 & ~n2079 ) | ( n1858 & ~n2079 ) ;
  assign n2083 = ( n56 & n1860 ) | ( n56 & ~n2082 ) | ( n1860 & ~n2082 ) ;
  assign n2084 = ( n56 & ~n1850 ) | ( n56 & n2082 ) | ( ~n1850 & n2082 ) ;
  assign n2085 = n1838 ^ n1776 ^ 1'b0 ;
  assign n2086 = ~n2083 & n2084 ;
  assign n2087 = ( n1838 & n1858 ) | ( n1838 & ~n2085 ) | ( n1858 & ~n2085 ) ;
  assign n2088 = ( n75 & ~n1850 ) | ( n75 & n2087 ) | ( ~n1850 & n2087 ) ;
  assign n2089 = ( n75 & n1860 ) | ( n75 & ~n2087 ) | ( n1860 & ~n2087 ) ;
  assign n2090 = n2088 & ~n2089 ;
  assign n2091 = n2081 ^ n2049 ^ n2029 ;
  assign n2092 = ( n2029 & ~n2049 ) | ( n2029 & n2081 ) | ( ~n2049 & n2081 ) ;
  assign n2093 = n2091 ^ n2048 ^ n2037 ;
  assign n2094 = ( ~n1605 & n2041 ) | ( ~n1605 & n2093 ) | ( n2041 & n2093 ) ;
  assign n2095 = n2093 ^ n2041 ^ n1605 ;
  assign n2096 = n1838 ^ n38 ^ 1'b0 ;
  assign n2097 = ( n1838 & n1858 ) | ( n1838 & ~n2096 ) | ( n1858 & ~n2096 ) ;
  assign n2098 = ( n1776 & n1860 ) | ( n1776 & ~n2097 ) | ( n1860 & ~n2097 ) ;
  assign n2099 = ( n1776 & ~n1850 ) | ( n1776 & n2097 ) | ( ~n1850 & n2097 ) ;
  assign n2100 = ~n2098 & n2099 ;
  assign n2101 = n44 & n1409 ;
  assign n2102 = ( n2037 & ~n2048 ) | ( n2037 & n2091 ) | ( ~n2048 & n2091 ) ;
  assign n2103 = ( n1718 & n2065 ) | ( n1718 & ~n2101 ) | ( n2065 & ~n2101 ) ;
  assign n2104 = n2101 ^ n2065 ^ n1718 ;
  assign n2105 = ( n2033 & n2057 ) | ( n2033 & n2100 ) | ( n2057 & n2100 ) ;
  assign n2106 = n2100 ^ n2057 ^ n2033 ;
  assign n2107 = n1838 ^ n56 ^ 1'b0 ;
  assign n2108 = n2106 ^ n2104 ^ n2077 ;
  assign n2109 = n2108 ^ n2080 ^ n2047 ;
  assign n2110 = ( n1838 & n1858 ) | ( n1838 & ~n2107 ) | ( n1858 & ~n2107 ) ;
  assign n2111 = n2109 ^ n2102 ^ n2092 ;
  assign n2112 = ( n1654 & ~n1850 ) | ( n1654 & n2110 ) | ( ~n1850 & n2110 ) ;
  assign n2113 = ( n2077 & ~n2104 ) | ( n2077 & n2106 ) | ( ~n2104 & n2106 ) ;
  assign n2114 = ( n1654 & n1860 ) | ( n1654 & ~n2110 ) | ( n1860 & ~n2110 ) ;
  assign n2115 = ( n2047 & n2080 ) | ( n2047 & ~n2108 ) | ( n2080 & ~n2108 ) ;
  assign n2116 = n2112 & ~n2114 ;
  assign n2117 = n2111 ^ n2094 ^ n1416 ;
  assign n2118 = ( ~n2092 & n2102 ) | ( ~n2092 & n2109 ) | ( n2102 & n2109 ) ;
  assign n2119 = ( ~n1416 & n2094 ) | ( ~n1416 & n2111 ) | ( n2094 & n2111 ) ;
  assign n2120 = n1409 & n1695 ;
  assign n2121 = ~n79 & n1918 ;
  assign n2122 = ( ~n1701 & n2101 ) | ( ~n1701 & n2120 ) | ( n2101 & n2120 ) ;
  assign n2123 = n79 & n1852 ;
  assign n2124 = ~n38 & n1853 ;
  assign n2125 = ( n2121 & n2123 ) | ( n2121 & ~n2124 ) | ( n2123 & ~n2124 ) ;
  assign n2126 = n1695 ^ n44 ^ 1'b0 ;
  assign n2127 = ( n2061 & n2090 ) | ( n2061 & n2125 ) | ( n2090 & n2125 ) ;
  assign n2128 = n2125 ^ n2090 ^ n2061 ;
  assign n2129 = n1409 & n2126 ;
  assign n2130 = n2129 ^ n1701 ^ 1'b0 ;
  assign n2131 = n2130 ^ n2105 ^ n2103 ;
  assign n2132 = ( n2103 & n2105 ) | ( n2103 & ~n2130 ) | ( n2105 & ~n2130 ) ;
  assign n2133 = n2131 ^ n2128 ^ n2113 ;
  assign n2134 = n2133 ^ n2118 ^ n2115 ;
  assign n2135 = n2134 ^ n2119 ^ n1510 ;
  assign n2136 = ( ~n1510 & n2119 ) | ( ~n1510 & n2134 ) | ( n2119 & n2134 ) ;
  assign n2137 = n1852 ^ n1776 ^ 1'b0 ;
  assign n2138 = n75 & n1853 ;
  assign n2139 = ( n1852 & n1918 ) | ( n1852 & ~n2137 ) | ( n1918 & ~n2137 ) ;
  assign n2140 = ( ~n1853 & n2138 ) | ( ~n1853 & n2139 ) | ( n2138 & n2139 ) ;
  assign n2141 = n79 & n1409 ;
  assign n2142 = ( ~n2115 & n2118 ) | ( ~n2115 & n2133 ) | ( n2118 & n2133 ) ;
  assign n2143 = n1852 ^ n75 ^ 1'b0 ;
  assign n2144 = ( n1852 & n1918 ) | ( n1852 & ~n2143 ) | ( n1918 & ~n2143 ) ;
  assign n2145 = n56 & n1853 ;
  assign n2146 = ( ~n1853 & n2144 ) | ( ~n1853 & n2145 ) | ( n2144 & n2145 ) ;
  assign n2147 = ( n2113 & n2128 ) | ( n2113 & ~n2131 ) | ( n2128 & ~n2131 ) ;
  assign n2148 = ~n1776 & n1853 ;
  assign n2149 = ~n38 & n1918 ;
  assign n2150 = n38 & n1852 ;
  assign n2151 = ( ~n2148 & n2149 ) | ( ~n2148 & n2150 ) | ( n2149 & n2150 ) ;
  assign n2152 = ( n2068 & n2086 ) | ( n2068 & ~n2141 ) | ( n2086 & ~n2141 ) ;
  assign n2153 = n2152 ^ n2140 ^ n2116 ;
  assign n2154 = ( n2116 & n2140 ) | ( n2116 & n2152 ) | ( n2140 & n2152 ) ;
  assign n2155 = n38 & n1409 ;
  assign n2156 = n2151 ^ n2127 ^ n2122 ;
  assign n2157 = ( n2122 & n2127 ) | ( n2122 & n2151 ) | ( n2127 & n2151 ) ;
  assign n2158 = n1409 & n1776 ;
  assign n2159 = ( n2063 & n2146 ) | ( n2063 & ~n2158 ) | ( n2146 & ~n2158 ) ;
  assign n2160 = n2158 ^ n2146 ^ n2063 ;
  assign n2161 = n2141 ^ n2086 ^ n2068 ;
  assign n2162 = n2161 ^ n2156 ^ n2132 ;
  assign n2163 = n2162 ^ n2147 ^ n2142 ;
  assign n2164 = ( n2142 & ~n2147 ) | ( n2142 & n2162 ) | ( ~n2147 & n2162 ) ;
  assign n2165 = n2155 ^ n2141 ^ n1761 ;
  assign n2166 = ( n2153 & n2157 ) | ( n2153 & ~n2165 ) | ( n2157 & ~n2165 ) ;
  assign n2167 = ( n2132 & n2156 ) | ( n2132 & ~n2161 ) | ( n2156 & ~n2161 ) ;
  assign n2168 = ( ~n1761 & n2141 ) | ( ~n1761 & n2155 ) | ( n2141 & n2155 ) ;
  assign n2169 = n2163 ^ n2136 ^ n1604 ;
  assign n2170 = n2168 ^ n2160 ^ n2154 ;
  assign n2171 = n2165 ^ n2157 ^ n2153 ;
  assign n2172 = n2171 ^ n2167 ^ n2164 ;
  assign n2173 = ( ~n1604 & n2136 ) | ( ~n1604 & n2163 ) | ( n2136 & n2163 ) ;
  assign n2174 = n2173 ^ n2172 ^ n1411 ;
  assign n2175 = ( n2164 & ~n2167 ) | ( n2164 & n2171 ) | ( ~n2167 & n2171 ) ;
  assign n2176 = n2175 ^ n2170 ^ n2166 ;
  assign n2177 = ( n1411 & n2172 ) | ( n1411 & n2173 ) | ( n2172 & n2173 ) ;
  assign n2178 = ( ~n1608 & n2176 ) | ( ~n1608 & n2177 ) | ( n2176 & n2177 ) ;
  assign n2179 = ( n2154 & ~n2160 ) | ( n2154 & n2168 ) | ( ~n2160 & n2168 ) ;
  assign n2180 = ( ~n2166 & n2170 ) | ( ~n2166 & n2175 ) | ( n2170 & n2175 ) ;
  assign n2181 = n2177 ^ n2176 ^ n1608 ;
  assign n2182 = n52 ^ n44 ^ 1'b0 ;
  assign n2183 = n75 & n1409 ;
  assign n2184 = n2183 ^ n2158 ^ n1846 ;
  assign n2185 = ( ~n1846 & n2158 ) | ( ~n1846 & n2183 ) | ( n2158 & n2183 ) ;
  assign n2186 = n1654 & n1853 ;
  assign n2187 = n1852 ^ n56 ^ 1'b0 ;
  assign n2188 = ( n1852 & n1918 ) | ( n1852 & ~n2187 ) | ( n1918 & ~n2187 ) ;
  assign n2189 = ( ~n1853 & n2186 ) | ( ~n1853 & n2188 ) | ( n2186 & n2188 ) ;
  assign n2190 = n2189 ^ n2184 ^ n2159 ;
  assign n2191 = ( n2159 & ~n2184 ) | ( n2159 & n2189 ) | ( ~n2184 & n2189 ) ;
  assign n2192 = n2186 ^ n1654 ^ n1409 ;
  assign n2193 = ( n1409 & n1852 ) | ( n1409 & n2192 ) | ( n1852 & n2192 ) ;
  assign n2194 = n56 & n1409 ;
  assign n2195 = ( n2185 & n2193 ) | ( n2185 & ~n2194 ) | ( n2193 & ~n2194 ) ;
  assign n2196 = n2194 ^ n2193 ^ n2185 ;
  assign n2197 = ( ~n2179 & n2180 ) | ( ~n2179 & n2190 ) | ( n2180 & n2190 ) ;
  assign n2198 = n1654 ^ n56 ^ 1'b0 ;
  assign n2199 = n2190 ^ n2180 ^ n2179 ;
  assign n2200 = n2199 ^ n2178 ^ n1609 ;
  assign n2201 = ( ~n1609 & n2178 ) | ( ~n1609 & n2199 ) | ( n2178 & n2199 ) ;
  assign n2202 = n2198 ^ n1853 ^ n1852 ;
  assign n2203 = ( ~n2191 & n2196 ) | ( ~n2191 & n2197 ) | ( n2196 & n2197 ) ;
  assign n2204 = n1409 & ~n2202 ;
  assign n2205 = n2197 ^ n2196 ^ n2191 ;
  assign n2206 = n2204 ^ n2203 ^ n2195 ;
  assign n2207 = ( ~n632 & n2201 ) | ( ~n632 & n2205 ) | ( n2201 & n2205 ) ;
  assign n2208 = ( n1549 & n2206 ) | ( n1549 & n2207 ) | ( n2206 & n2207 ) ;
  assign n2209 = ~n1610 & n2208 ;
  assign n2210 = ~n480 & n2209 ;
  assign n2211 = n1616 & n2210 ;
  assign n2212 = ~n1584 & n2211 ;
  assign n2213 = n1586 & n2212 ;
  assign n2214 = n1636 ^ n52 ^ 1'b0 ;
  assign n2215 = n1409 | n1563 ;
  assign n2216 = n2212 ^ n1586 ^ 1'b0 ;
  assign n2217 = n2205 ^ n2201 ^ n632 ;
  assign n2218 = n1409 | n1590 ;
  assign n2219 = n2208 ^ n1610 ^ 1'b0 ;
  assign n2220 = n2209 ^ n480 ^ 1'b0 ;
  assign n2221 = n2210 ^ n1616 ^ 1'b0 ;
  assign n2222 = n2211 ^ n1584 ^ 1'b0 ;
  assign n2223 = n2207 ^ n2206 ^ n1549 ;
  assign n2224 = n2213 ^ n2212 ^ n1595 ;
  assign n2225 = ( ~x21 & x22 ) | ( ~x21 & n66 ) | ( x22 & n66 ) ;
  assign n2226 = n27 & ~n2042 ;
  assign n2227 = n26 & ~n2014 ;
  assign n2228 = ( n26 & n2018 ) | ( n26 & n2226 ) | ( n2018 & n2226 ) ;
  assign n2229 = n2014 & n2018 ;
  assign n2230 = ( x0 & x1 ) | ( x0 & x22 ) | ( x1 & x22 ) ;
  assign n2231 = n27 & n2018 ;
  assign n2232 = x1 & n2230 ;
  assign n2233 = n2232 ^ x2 ^ 1'b0 ;
  assign n2234 = n2226 | n2228 ;
  assign n2235 = x0 & ~n2233 ;
  assign n2236 = ( ~n2042 & n2231 ) | ( ~n2042 & n2235 ) | ( n2231 & n2235 ) ;
  assign n2237 = x0 & n2014 ;
  assign n2238 = n2018 ^ n2014 ^ 1'b0 ;
  assign n2239 = ( x0 & ~x22 ) | ( x0 & n27 ) | ( ~x22 & n27 ) ;
  assign n2240 = n2239 ^ x2 ^ 1'b0 ;
  assign n2241 = n27 & n2014 ;
  assign n2242 = ( n2018 & n2235 ) | ( n2018 & ~n2240 ) | ( n2235 & ~n2240 ) ;
  assign n2243 = n2240 & ~n2242 ;
  assign n2244 = ~n2241 & n2243 ;
  assign n2245 = n2231 | n2236 ;
  assign n2246 = ( n26 & ~n2227 ) | ( n26 & n2245 ) | ( ~n2227 & n2245 ) ;
  assign n2247 = n2169 & ~n2235 ;
  assign n2248 = n2229 ^ n2042 ^ n2018 ;
  assign n2249 = x0 & n2233 ;
  assign n2250 = n27 & n2135 ;
  assign n2251 = ( n26 & n2117 ) | ( n26 & n2250 ) | ( n2117 & n2250 ) ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = ( n2169 & ~n2247 ) | ( n2169 & n2252 ) | ( ~n2247 & n2252 ) ;
  assign n2254 = n2240 & n2249 ;
  assign n2255 = n2238 & n2254 ;
  assign n2256 = ~n2248 & n2254 ;
  assign n2257 = ( n2240 & n2246 ) | ( n2240 & n2256 ) | ( n2246 & n2256 ) ;
  assign n2258 = ( n2244 & n2255 ) | ( n2244 & ~n2256 ) | ( n2255 & ~n2256 ) ;
  assign n2259 = ~n2255 & n2258 ;
  assign n2260 = n27 & n2095 ;
  assign n2261 = ( ~n2237 & n2257 ) | ( ~n2237 & n2259 ) | ( n2257 & n2259 ) ;
  assign n2262 = n27 & n2117 ;
  assign n2263 = ( n26 & n2095 ) | ( n26 & n2262 ) | ( n2095 & n2262 ) ;
  assign n2264 = n2262 | n2263 ;
  assign n2265 = n75 ^ n56 ^ 1'b0 ;
  assign n2266 = ~n2257 & n2261 ;
  assign n2267 = n2135 & ~n2235 ;
  assign n2268 = ( n26 & ~n2042 ) | ( n26 & n2260 ) | ( ~n2042 & n2260 ) ;
  assign n2269 = n1776 ^ n75 ^ 1'b0 ;
  assign n2270 = n2260 | n2268 ;
  assign n2271 = ( n2135 & n2264 ) | ( n2135 & ~n2267 ) | ( n2264 & ~n2267 ) ;
  assign n2272 = n27 & n2169 ;
  assign n2273 = ( ~n2174 & n2235 ) | ( ~n2174 & n2272 ) | ( n2235 & n2272 ) ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = n2117 & ~n2235 ;
  assign n2276 = ( n2117 & n2270 ) | ( n2117 & ~n2275 ) | ( n2270 & ~n2275 ) ;
  assign n2277 = n26 & ~n2135 ;
  assign n2278 = ( n26 & n2274 ) | ( n26 & ~n2277 ) | ( n2274 & ~n2277 ) ;
  assign n2279 = n84 ^ n70 ^ 1'b0 ;
  assign n2280 = n1636 ^ n70 ^ 1'b0 ;
  assign n2281 = n2240 ^ n84 ^ 1'b0 ;
  assign n2282 = n2279 & ~n2281 ;
  assign n2283 = ~n2014 & n2282 ;
  assign n2284 = ~n2279 & n2280 ;
  assign n2285 = ~n2280 & n2281 ;
  assign n2286 = n2018 & n2285 ;
  assign n2287 = ( n2282 & ~n2283 ) | ( n2282 & n2286 ) | ( ~n2283 & n2286 ) ;
  assign n2288 = n2280 & n2281 ;
  assign n2289 = ( n2238 & n2286 ) | ( n2238 & n2288 ) | ( n2286 & n2288 ) ;
  assign n2290 = n2287 | n2289 ;
  assign n2291 = n2290 ^ n1635 ^ x5 ;
  assign n2292 = n2014 & n2281 ;
  assign n2293 = n1636 & ~n2292 ;
  assign n2294 = ~n2281 & n2284 ;
  assign n2295 = n2018 & ~n2042 ;
  assign n2296 = ( n2014 & n2018 ) | ( n2014 & n2295 ) | ( n2018 & n2295 ) ;
  assign n2297 = ( ~n2042 & n2095 ) | ( ~n2042 & n2296 ) | ( n2095 & n2296 ) ;
  assign n2298 = n2296 ^ n2095 ^ n2042 ;
  assign n2299 = n2095 & ~n2235 ;
  assign n2300 = ( n2095 & n2234 ) | ( n2095 & ~n2299 ) | ( n2234 & ~n2299 ) ;
  assign n2301 = n2249 & n2298 ;
  assign n2302 = ( n2249 & n2300 ) | ( n2249 & ~n2301 ) | ( n2300 & ~n2301 ) ;
  assign n2303 = n2302 ^ n2239 ^ x2 ;
  assign n2304 = n2291 & n2293 ;
  assign n2305 = ( n2266 & n2292 ) | ( n2266 & n2303 ) | ( n2292 & n2303 ) ;
  assign n2306 = n2297 ^ n2117 ^ n2095 ;
  assign n2307 = n2293 ^ n2291 ^ 1'b0 ;
  assign n2308 = n2254 & n2306 ;
  assign n2309 = n2305 & ~n2307 ;
  assign n2310 = n2305 | n2307 ;
  assign n2311 = ~n2308 & n2310 ;
  assign n2312 = ~n2249 & n2306 ;
  assign n2313 = ( n2276 & n2306 ) | ( n2276 & ~n2312 ) | ( n2306 & ~n2312 ) ;
  assign n2314 = ( n2240 & n2276 ) | ( n2240 & ~n2311 ) | ( n2276 & ~n2311 ) ;
  assign n2315 = ( n2240 & n2311 ) | ( n2240 & n2313 ) | ( n2311 & n2313 ) ;
  assign n2316 = ( n2095 & n2117 ) | ( n2095 & n2297 ) | ( n2117 & n2297 ) ;
  assign n2317 = x21 | n2225 ;
  assign n2318 = ( n2117 & n2135 ) | ( n2117 & n2316 ) | ( n2135 & n2316 ) ;
  assign n2319 = ~n2314 & n2315 ;
  assign n2320 = ~n2014 & n2294 ;
  assign n2321 = n2316 ^ n2135 ^ n2117 ;
  assign n2322 = ( n2305 & ~n2309 ) | ( n2305 & n2319 ) | ( ~n2309 & n2319 ) ;
  assign n2323 = n2018 & n2282 ;
  assign n2324 = ( n2294 & ~n2320 ) | ( n2294 & n2323 ) | ( ~n2320 & n2323 ) ;
  assign n2325 = ~n2249 & n2321 ;
  assign n2326 = ( n2271 & n2321 ) | ( n2271 & ~n2325 ) | ( n2321 & ~n2325 ) ;
  assign n2327 = n2326 ^ n2239 ^ x2 ;
  assign n2328 = ~n2042 & n2285 ;
  assign n2329 = ( ~n2248 & n2288 ) | ( ~n2248 & n2328 ) | ( n2288 & n2328 ) ;
  assign n2330 = ( n2324 & ~n2328 ) | ( n2324 & n2329 ) | ( ~n2328 & n2329 ) ;
  assign n2331 = n2328 | n2330 ;
  assign n2332 = n2331 ^ n1635 ^ x5 ;
  assign n2333 = n2304 & n2332 ;
  assign n2334 = n2332 ^ n2304 ^ 1'b0 ;
  assign n2335 = ( n2322 & n2327 ) | ( n2322 & n2334 ) | ( n2327 & n2334 ) ;
  assign n2336 = n2095 & n2285 ;
  assign n2337 = ( ~n2042 & n2282 ) | ( ~n2042 & n2336 ) | ( n2282 & n2336 ) ;
  assign n2338 = n2336 | n2337 ;
  assign n2339 = n2018 & ~n2294 ;
  assign n2340 = n2318 ^ n2169 ^ n2135 ;
  assign n2341 = n2254 & n2340 ;
  assign n2342 = ( n2018 & n2338 ) | ( n2018 & ~n2339 ) | ( n2338 & ~n2339 ) ;
  assign n2343 = ~n2249 & n2340 ;
  assign n2344 = n2014 & n2214 ;
  assign n2345 = n2288 & n2298 ;
  assign n2346 = ( n2288 & n2342 ) | ( n2288 & ~n2345 ) | ( n2342 & ~n2345 ) ;
  assign n2347 = n2346 ^ n1635 ^ x5 ;
  assign n2348 = ( n2333 & n2344 ) | ( n2333 & n2347 ) | ( n2344 & n2347 ) ;
  assign n2349 = n2347 ^ n2344 ^ n2333 ;
  assign n2350 = n2335 | n2349 ;
  assign n2351 = ~n2341 & n2350 ;
  assign n2352 = ( n2240 & n2253 ) | ( n2240 & ~n2351 ) | ( n2253 & ~n2351 ) ;
  assign n2353 = ( n2253 & n2340 ) | ( n2253 & ~n2343 ) | ( n2340 & ~n2343 ) ;
  assign n2354 = ( n2240 & n2351 ) | ( n2240 & n2353 ) | ( n2351 & n2353 ) ;
  assign n2355 = ~n2352 & n2354 ;
  assign n2356 = n2335 & ~n2349 ;
  assign n2357 = n2126 & n2214 ;
  assign n2358 = ( n2335 & n2355 ) | ( n2335 & ~n2356 ) | ( n2355 & ~n2356 ) ;
  assign n2359 = n2238 & n2357 ;
  assign n2360 = ~n2126 & n2214 ;
  assign n2361 = n2182 & ~n2214 ;
  assign n2362 = ( n2014 & n2359 ) | ( n2014 & n2361 ) | ( n2359 & n2361 ) ;
  assign n2363 = ( n2135 & n2169 ) | ( n2135 & n2318 ) | ( n2169 & n2318 ) ;
  assign n2364 = ( n2126 & ~n2182 ) | ( n2126 & n2214 ) | ( ~n2182 & n2214 ) ;
  assign n2365 = n1695 & ~n2344 ;
  assign n2366 = ~n2018 & n2360 ;
  assign n2367 = ( n2359 & n2360 ) | ( n2359 & ~n2366 ) | ( n2360 & ~n2366 ) ;
  assign n2368 = n2362 | n2367 ;
  assign n2369 = n2368 ^ n1678 ^ x8 ;
  assign n2370 = n2117 & n2285 ;
  assign n2371 = ( ~n2042 & n2294 ) | ( ~n2042 & n2370 ) | ( n2294 & n2370 ) ;
  assign n2372 = n2370 | n2371 ;
  assign n2373 = n2095 & ~n2282 ;
  assign n2374 = ( n2095 & n2372 ) | ( n2095 & ~n2373 ) | ( n2372 & ~n2373 ) ;
  assign n2375 = n2288 & ~n2306 ;
  assign n2376 = ( n2288 & n2374 ) | ( n2288 & ~n2375 ) | ( n2374 & ~n2375 ) ;
  assign n2377 = n2365 & n2369 ;
  assign n2378 = n2376 ^ n1635 ^ x5 ;
  assign n2379 = n2369 ^ n2365 ^ 1'b0 ;
  assign n2380 = n2379 ^ n2378 ^ n2348 ;
  assign n2381 = ( n2348 & n2378 ) | ( n2348 & n2379 ) | ( n2378 & n2379 ) ;
  assign n2382 = n2363 ^ n2174 ^ n2169 ;
  assign n2383 = n2249 & n2382 ;
  assign n2384 = ( n2249 & n2278 ) | ( n2249 & ~n2383 ) | ( n2278 & ~n2383 ) ;
  assign n2385 = n2169 & n2361 ;
  assign n2386 = ~n2214 & n2364 ;
  assign n2387 = n2384 ^ n2239 ^ x2 ;
  assign n2388 = ( n2358 & n2380 ) | ( n2358 & n2387 ) | ( n2380 & n2387 ) ;
  assign n2389 = ( ~n2174 & n2360 ) | ( ~n2174 & n2385 ) | ( n2360 & n2385 ) ;
  assign n2390 = n2385 | n2389 ;
  assign n2391 = n2135 & ~n2386 ;
  assign n2392 = ( n2135 & n2390 ) | ( n2135 & ~n2391 ) | ( n2390 & ~n2391 ) ;
  assign n2393 = ( n2360 & n2382 ) | ( n2360 & ~n2392 ) | ( n2382 & ~n2392 ) ;
  assign n2394 = ( n2214 & n2392 ) | ( n2214 & ~n2393 ) | ( n2392 & ~n2393 ) ;
  assign n2395 = n2394 ^ n1678 ^ x8 ;
  assign n2396 = n79 ^ n38 ^ 1'b0 ;
  assign n2397 = n1776 ^ n38 ^ 1'b0 ;
  assign n2398 = n1695 ^ n79 ^ 1'b0 ;
  assign n2399 = ~n2396 & n2397 ;
  assign n2400 = ~n2398 & n2399 ;
  assign n2401 = ~n2014 & n2400 ;
  assign n2402 = ~n2397 & n2398 ;
  assign n2403 = ~n2042 & n2402 ;
  assign n2404 = n2018 & n2361 ;
  assign n2405 = ~n2014 & n2386 ;
  assign n2406 = ~n2042 & n2360 ;
  assign n2407 = ( ~n2248 & n2357 ) | ( ~n2248 & n2406 ) | ( n2357 & n2406 ) ;
  assign n2408 = ( n2386 & n2404 ) | ( n2386 & ~n2405 ) | ( n2404 & ~n2405 ) ;
  assign n2409 = ( ~n2406 & n2407 ) | ( ~n2406 & n2408 ) | ( n2407 & n2408 ) ;
  assign n2410 = n2095 & n2360 ;
  assign n2411 = n2396 & ~n2398 ;
  assign n2412 = n2397 & n2398 ;
  assign n2413 = n2018 & n2411 ;
  assign n2414 = ( n2400 & ~n2401 ) | ( n2400 & n2413 ) | ( ~n2401 & n2413 ) ;
  assign n2415 = ( ~n2042 & n2361 ) | ( ~n2042 & n2410 ) | ( n2361 & n2410 ) ;
  assign n2416 = n2410 | n2415 ;
  assign n2417 = n2014 & n2398 ;
  assign n2418 = ( ~n2248 & n2403 ) | ( ~n2248 & n2412 ) | ( n2403 & n2412 ) ;
  assign n2419 = ( ~n2403 & n2414 ) | ( ~n2403 & n2418 ) | ( n2414 & n2418 ) ;
  assign n2420 = n2018 & ~n2386 ;
  assign n2421 = ( n2018 & n2416 ) | ( n2018 & ~n2420 ) | ( n2416 & ~n2420 ) ;
  assign n2422 = n2018 & n2402 ;
  assign n2423 = n2406 | n2409 ;
  assign n2424 = n2423 ^ n1678 ^ x8 ;
  assign n2425 = ~n2014 & n2411 ;
  assign n2426 = ( n2411 & n2422 ) | ( n2411 & ~n2425 ) | ( n2422 & ~n2425 ) ;
  assign n2427 = ( n2238 & n2412 ) | ( n2238 & n2422 ) | ( n2412 & n2422 ) ;
  assign n2428 = n2403 | n2419 ;
  assign n2429 = n2424 ^ n2377 ^ 1'b0 ;
  assign n2430 = n2426 | n2427 ;
  assign n2431 = n2377 & n2424 ;
  assign n2432 = n2298 & n2357 ;
  assign n2433 = n1776 & ~n2417 ;
  assign n2434 = ( n2357 & n2421 ) | ( n2357 & ~n2432 ) | ( n2421 & ~n2432 ) ;
  assign n2435 = n2430 ^ n40 ^ x11 ;
  assign n2436 = n2435 ^ n2433 ^ 1'b0 ;
  assign n2437 = n2433 & n2435 ;
  assign n2438 = n2434 ^ n1678 ^ x8 ;
  assign n2439 = n2438 ^ n2431 ^ n2417 ;
  assign n2440 = ( n2417 & n2431 ) | ( n2417 & n2438 ) | ( n2431 & n2438 ) ;
  assign n2441 = n2117 & n2360 ;
  assign n2442 = ( ~n2042 & n2386 ) | ( ~n2042 & n2441 ) | ( n2386 & n2441 ) ;
  assign n2443 = n2441 | n2442 ;
  assign n2444 = n2095 & ~n2361 ;
  assign n2445 = ( n2095 & n2443 ) | ( n2095 & ~n2444 ) | ( n2443 & ~n2444 ) ;
  assign n2446 = ~n2306 & n2357 ;
  assign n2447 = n2428 ^ n40 ^ x11 ;
  assign n2448 = ( n2357 & n2445 ) | ( n2357 & ~n2446 ) | ( n2445 & ~n2446 ) ;
  assign n2449 = n2448 ^ n1678 ^ x8 ;
  assign n2450 = ( n2436 & n2440 ) | ( n2436 & n2449 ) | ( n2440 & n2449 ) ;
  assign n2451 = n2449 ^ n2440 ^ n2436 ;
  assign n2452 = n2437 & n2447 ;
  assign n2453 = n2447 ^ n2437 ^ 1'b0 ;
  assign n2454 = n2095 & n2402 ;
  assign n2455 = n2265 & ~n2269 ;
  assign n2456 = ~n2014 & n2455 ;
  assign n2457 = ( n2198 & ~n2265 ) | ( n2198 & n2269 ) | ( ~n2265 & n2269 ) ;
  assign n2458 = ( ~n2042 & n2411 ) | ( ~n2042 & n2454 ) | ( n2411 & n2454 ) ;
  assign n2459 = n2454 | n2458 ;
  assign n2460 = ~n2198 & n2269 ;
  assign n2461 = n2198 & n2269 ;
  assign n2462 = n2018 & ~n2400 ;
  assign n2463 = ( n2018 & n2459 ) | ( n2018 & ~n2462 ) | ( n2459 & ~n2462 ) ;
  assign n2464 = n2018 & n2460 ;
  assign n2465 = ( n2238 & n2461 ) | ( n2238 & n2464 ) | ( n2461 & n2464 ) ;
  assign n2466 = ~n2269 & n2457 ;
  assign n2467 = ( n2455 & ~n2456 ) | ( n2455 & n2464 ) | ( ~n2456 & n2464 ) ;
  assign n2468 = n2465 | n2467 ;
  assign n2469 = n2018 & n2455 ;
  assign n2470 = n2298 & ~n2463 ;
  assign n2471 = ( n2412 & n2463 ) | ( n2412 & ~n2470 ) | ( n2463 & ~n2470 ) ;
  assign n2472 = n2471 ^ n40 ^ x11 ;
  assign n2473 = ~n2014 & n2466 ;
  assign n2474 = ( n2466 & n2469 ) | ( n2466 & ~n2473 ) | ( n2469 & ~n2473 ) ;
  assign n2475 = ~n2042 & n2460 ;
  assign n2476 = ( ~n2248 & n2461 ) | ( ~n2248 & n2475 ) | ( n2461 & n2475 ) ;
  assign n2477 = ( n2474 & ~n2475 ) | ( n2474 & n2476 ) | ( ~n2475 & n2476 ) ;
  assign n2478 = n2468 ^ n82 ^ x14 ;
  assign n2479 = n2475 | n2477 ;
  assign n2480 = n2095 & n2460 ;
  assign n2481 = n2298 & n2461 ;
  assign n2482 = ( ~n2042 & n2455 ) | ( ~n2042 & n2480 ) | ( n2455 & n2480 ) ;
  assign n2483 = n2480 | n2482 ;
  assign n2484 = n2018 & ~n2466 ;
  assign n2485 = ( n2018 & n2483 ) | ( n2018 & ~n2484 ) | ( n2483 & ~n2484 ) ;
  assign n2486 = n1654 & n2014 ;
  assign n2487 = n2014 & n2269 ;
  assign n2488 = n2487 ^ n2472 ^ n2452 ;
  assign n2489 = ( n2452 & n2472 ) | ( n2452 & n2487 ) | ( n2472 & n2487 ) ;
  assign n2490 = n1654 & ~n2487 ;
  assign n2491 = n2490 ^ n2478 ^ 1'b0 ;
  assign n2492 = n2478 & n2490 ;
  assign n2493 = ( n2461 & ~n2481 ) | ( n2461 & n2485 ) | ( ~n2481 & n2485 ) ;
  assign n2494 = n2479 ^ n82 ^ x14 ;
  assign n2495 = n2492 & n2494 ;
  assign n2496 = n2493 ^ n82 ^ x14 ;
  assign n2497 = ( n2486 & n2495 ) | ( n2486 & n2496 ) | ( n2495 & n2496 ) ;
  assign n2498 = n2496 ^ n2495 ^ n2486 ;
  assign n2499 = n2117 & n2402 ;
  assign n2500 = ( ~n2042 & n2400 ) | ( ~n2042 & n2499 ) | ( n2400 & n2499 ) ;
  assign n2501 = n2499 | n2500 ;
  assign n2502 = n2095 & ~n2411 ;
  assign n2503 = ( n2095 & n2501 ) | ( n2095 & ~n2502 ) | ( n2501 & ~n2502 ) ;
  assign n2504 = ~n2306 & n2461 ;
  assign n2505 = ~n2306 & n2412 ;
  assign n2506 = n1654 & n2018 ;
  assign n2507 = ( n2412 & n2503 ) | ( n2412 & ~n2505 ) | ( n2503 & ~n2505 ) ;
  assign n2508 = n2117 & n2460 ;
  assign n2509 = n2494 ^ n2492 ^ 1'b0 ;
  assign n2510 = ( ~n2042 & n2466 ) | ( ~n2042 & n2508 ) | ( n2466 & n2508 ) ;
  assign n2511 = n2508 | n2510 ;
  assign n2512 = n2095 & ~n2455 ;
  assign n2513 = ( n2095 & n2511 ) | ( n2095 & ~n2512 ) | ( n2511 & ~n2512 ) ;
  assign n2514 = ( n2461 & ~n2504 ) | ( n2461 & n2513 ) | ( ~n2504 & n2513 ) ;
  assign n2515 = n2514 ^ n82 ^ x14 ;
  assign n2516 = ( n2497 & n2506 ) | ( n2497 & n2515 ) | ( n2506 & n2515 ) ;
  assign n2517 = n2507 ^ n40 ^ x11 ;
  assign n2518 = n2517 ^ n2491 ^ n2489 ;
  assign n2519 = ( n2489 & n2491 ) | ( n2489 & n2517 ) | ( n2491 & n2517 ) ;
  assign n2520 = n2515 ^ n2506 ^ n2497 ;
  assign n2521 = n2135 & n2402 ;
  assign n2522 = ( n2095 & n2400 ) | ( n2095 & n2521 ) | ( n2400 & n2521 ) ;
  assign n2523 = n2521 | n2522 ;
  assign n2524 = n2117 & ~n2411 ;
  assign n2525 = ( n2117 & n2523 ) | ( n2117 & ~n2524 ) | ( n2523 & ~n2524 ) ;
  assign n2526 = ~n2321 & n2412 ;
  assign n2527 = ( n2412 & n2525 ) | ( n2412 & ~n2526 ) | ( n2525 & ~n2526 ) ;
  assign n2528 = n2527 ^ n40 ^ x11 ;
  assign n2529 = ( n2509 & n2519 ) | ( n2509 & n2528 ) | ( n2519 & n2528 ) ;
  assign n2530 = n2528 ^ n2519 ^ n2509 ;
  assign n2531 = n2135 & n2285 ;
  assign n2532 = ( n2095 & n2294 ) | ( n2095 & n2531 ) | ( n2294 & n2531 ) ;
  assign n2533 = n2531 | n2532 ;
  assign n2534 = n2117 & ~n2282 ;
  assign n2535 = ( n2117 & n2533 ) | ( n2117 & ~n2534 ) | ( n2533 & ~n2534 ) ;
  assign n2536 = n2288 & ~n2321 ;
  assign n2537 = ( n2288 & n2535 ) | ( n2288 & ~n2536 ) | ( n2535 & ~n2536 ) ;
  assign n2538 = n2537 ^ n1635 ^ x5 ;
  assign n2539 = n2538 ^ n2429 ^ n2381 ;
  assign n2540 = ( n2381 & n2429 ) | ( n2381 & n2538 ) | ( n2429 & n2538 ) ;
  assign n2541 = n2135 & n2360 ;
  assign n2542 = ( n2095 & n2386 ) | ( n2095 & n2541 ) | ( n2386 & n2541 ) ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = n2117 & ~n2361 ;
  assign n2545 = ( n2117 & n2543 ) | ( n2117 & ~n2544 ) | ( n2543 & ~n2544 ) ;
  assign n2546 = n2321 & ~n2357 ;
  assign n2547 = ( n2321 & n2545 ) | ( n2321 & ~n2546 ) | ( n2545 & ~n2546 ) ;
  assign n2548 = n2547 ^ n1678 ^ x8 ;
  assign n2549 = n2548 ^ n2453 ^ n2450 ;
  assign n2550 = ~n2321 & n2461 ;
  assign n2551 = ( n2450 & n2453 ) | ( n2450 & n2548 ) | ( n2453 & n2548 ) ;
  assign n2552 = n2135 & n2460 ;
  assign n2553 = ( n2095 & n2466 ) | ( n2095 & n2552 ) | ( n2466 & n2552 ) ;
  assign n2554 = n2552 | n2553 ;
  assign n2555 = n2117 & ~n2455 ;
  assign n2556 = ( n2117 & n2554 ) | ( n2117 & ~n2555 ) | ( n2554 & ~n2555 ) ;
  assign n2557 = ( n2461 & ~n2550 ) | ( n2461 & n2556 ) | ( ~n2550 & n2556 ) ;
  assign n2558 = n2169 & n2360 ;
  assign n2559 = ( n2117 & n2386 ) | ( n2117 & n2558 ) | ( n2386 & n2558 ) ;
  assign n2560 = n2558 | n2559 ;
  assign n2561 = n2135 & ~n2361 ;
  assign n2562 = ( n2135 & n2560 ) | ( n2135 & ~n2561 ) | ( n2560 & ~n2561 ) ;
  assign n2563 = n2340 & ~n2357 ;
  assign n2564 = ( n2340 & n2562 ) | ( n2340 & ~n2563 ) | ( n2562 & ~n2563 ) ;
  assign n2565 = n2564 ^ n1678 ^ x8 ;
  assign n2566 = ( n2488 & n2551 ) | ( n2488 & n2565 ) | ( n2551 & n2565 ) ;
  assign n2567 = n2565 ^ n2551 ^ n2488 ;
  assign n2568 = n2566 ^ n2518 ^ n2395 ;
  assign n2569 = ( n2395 & n2518 ) | ( n2395 & n2566 ) | ( n2518 & n2566 ) ;
  assign n2570 = n1654 & ~n2042 ;
  assign n2571 = n1654 & n2042 ;
  assign n2572 = n2571 ^ n2557 ^ n2516 ;
  assign n2573 = n2557 ^ n1654 ^ 1'b0 ;
  assign n2574 = ( n2516 & n2570 ) | ( n2516 & n2573 ) | ( n2570 & n2573 ) ;
  assign n2575 = n2169 & n2402 ;
  assign n2576 = ( n2117 & n2400 ) | ( n2117 & n2575 ) | ( n2400 & n2575 ) ;
  assign n2577 = n2575 | n2576 ;
  assign n2578 = n2135 & ~n2411 ;
  assign n2579 = ( n2135 & n2577 ) | ( n2135 & ~n2578 ) | ( n2577 & ~n2578 ) ;
  assign n2580 = ~n2340 & n2412 ;
  assign n2581 = ( n2412 & n2579 ) | ( n2412 & ~n2580 ) | ( n2579 & ~n2580 ) ;
  assign n2582 = n2581 ^ n40 ^ x11 ;
  assign n2583 = ( n2498 & n2529 ) | ( n2498 & n2582 ) | ( n2529 & n2582 ) ;
  assign n2584 = n2582 ^ n2529 ^ n2498 ;
  assign n2585 = n2169 & n2460 ;
  assign n2586 = ( n2117 & n2466 ) | ( n2117 & n2585 ) | ( n2466 & n2585 ) ;
  assign n2587 = n2585 | n2586 ;
  assign n2588 = n2135 & ~n2455 ;
  assign n2589 = ( n2135 & n2587 ) | ( n2135 & ~n2588 ) | ( n2587 & ~n2588 ) ;
  assign n2590 = ~n2340 & n2461 ;
  assign n2591 = ( n2461 & n2589 ) | ( n2461 & ~n2590 ) | ( n2589 & ~n2590 ) ;
  assign n2592 = n1654 & ~n2095 ;
  assign n2593 = n2592 ^ n2591 ^ n2574 ;
  assign n2594 = n2591 ^ n1654 ^ 1'b0 ;
  assign n2595 = n1654 & n2095 ;
  assign n2596 = ( n2574 & n2594 ) | ( n2574 & n2595 ) | ( n2594 & n2595 ) ;
  assign n2597 = n2169 & n2285 ;
  assign n2598 = ( n2117 & n2294 ) | ( n2117 & n2597 ) | ( n2294 & n2597 ) ;
  assign n2599 = n2597 | n2598 ;
  assign n2600 = n2288 & ~n2340 ;
  assign n2601 = n2135 & ~n2282 ;
  assign n2602 = ( n2135 & n2599 ) | ( n2135 & ~n2601 ) | ( n2599 & ~n2601 ) ;
  assign n2603 = ( n2288 & ~n2600 ) | ( n2288 & n2602 ) | ( ~n2600 & n2602 ) ;
  assign n2604 = n2603 ^ n1635 ^ x5 ;
  assign n2605 = n2169 & n2455 ;
  assign n2606 = ( ~n2174 & n2460 ) | ( ~n2174 & n2605 ) | ( n2460 & n2605 ) ;
  assign n2607 = n2605 | n2606 ;
  assign n2608 = n2135 & ~n2466 ;
  assign n2609 = ( n2135 & n2607 ) | ( n2135 & ~n2608 ) | ( n2607 & ~n2608 ) ;
  assign n2610 = n2604 ^ n2540 ^ n2439 ;
  assign n2611 = ( n2439 & n2540 ) | ( n2439 & n2604 ) | ( n2540 & n2604 ) ;
  assign n2612 = n2169 & n2411 ;
  assign n2613 = n2382 & n2461 ;
  assign n2614 = ( n2461 & n2609 ) | ( n2461 & ~n2613 ) | ( n2609 & ~n2613 ) ;
  assign n2615 = ( ~n2174 & n2402 ) | ( ~n2174 & n2612 ) | ( n2402 & n2612 ) ;
  assign n2616 = n2612 | n2615 ;
  assign n2617 = n2135 & ~n2400 ;
  assign n2618 = ( n2135 & n2616 ) | ( n2135 & ~n2617 ) | ( n2616 & ~n2617 ) ;
  assign n2619 = n2382 & n2412 ;
  assign n2620 = ( n2412 & n2618 ) | ( n2412 & ~n2619 ) | ( n2618 & ~n2619 ) ;
  assign n2621 = n1654 & n2117 ;
  assign n2622 = n1654 & ~n2117 ;
  assign n2623 = n2622 ^ n2614 ^ n2596 ;
  assign n2624 = n2620 ^ n40 ^ x11 ;
  assign n2625 = n2614 ^ n1654 ^ 1'b0 ;
  assign n2626 = ( n2596 & n2621 ) | ( n2596 & n2625 ) | ( n2621 & n2625 ) ;
  assign n2627 = n2169 & n2282 ;
  assign n2628 = ( ~n2174 & n2285 ) | ( ~n2174 & n2627 ) | ( n2285 & n2627 ) ;
  assign n2629 = n2627 | n2628 ;
  assign n2630 = n2135 & ~n2294 ;
  assign n2631 = ( n2135 & n2629 ) | ( n2135 & ~n2630 ) | ( n2629 & ~n2630 ) ;
  assign n2632 = n2288 & ~n2382 ;
  assign n2633 = n2631 | n2632 ;
  assign n2634 = n2633 ^ n1635 ^ x5 ;
  assign n2635 = n2634 ^ n2611 ^ n2451 ;
  assign n2636 = n2624 ^ n2583 ^ n2520 ;
  assign n2637 = ( n2451 & n2611 ) | ( n2451 & n2634 ) | ( n2611 & n2634 ) ;
  assign n2638 = ( n2520 & n2583 ) | ( n2520 & n2624 ) | ( n2583 & n2624 ) ;
  assign n2639 = ( n2169 & ~n2174 ) | ( n2169 & n2363 ) | ( ~n2174 & n2363 ) ;
  assign n2640 = n2169 & n2294 ;
  assign n2641 = ( ~n2174 & n2282 ) | ( ~n2174 & n2640 ) | ( n2282 & n2640 ) ;
  assign n2642 = n2169 & n2386 ;
  assign n2643 = n2640 | n2641 ;
  assign n2644 = n2181 & ~n2285 ;
  assign n2645 = ( n2181 & n2643 ) | ( n2181 & ~n2644 ) | ( n2643 & ~n2644 ) ;
  assign n2646 = ( ~n2174 & n2361 ) | ( ~n2174 & n2642 ) | ( n2361 & n2642 ) ;
  assign n2647 = n2642 | n2646 ;
  assign n2648 = n2639 ^ n2181 ^ n2174 ;
  assign n2649 = n2181 & ~n2360 ;
  assign n2650 = ( n2181 & n2647 ) | ( n2181 & ~n2649 ) | ( n2647 & ~n2649 ) ;
  assign n2651 = n2357 & n2648 ;
  assign n2652 = ( n2357 & n2650 ) | ( n2357 & ~n2651 ) | ( n2650 & ~n2651 ) ;
  assign n2653 = n2288 & ~n2648 ;
  assign n2654 = n2652 ^ n1678 ^ x8 ;
  assign n2655 = n2645 | n2653 ;
  assign n2656 = ( ~n2174 & n2181 ) | ( ~n2174 & n2639 ) | ( n2181 & n2639 ) ;
  assign n2657 = ( n2530 & n2569 ) | ( n2530 & n2654 ) | ( n2569 & n2654 ) ;
  assign n2658 = n2654 ^ n2569 ^ n2530 ;
  assign n2659 = n2388 & ~n2539 ;
  assign n2660 = n2655 ^ n1635 ^ x5 ;
  assign n2661 = n2254 & ~n2648 ;
  assign n2662 = ( n2388 & n2539 ) | ( n2388 & ~n2661 ) | ( n2539 & ~n2661 ) ;
  assign n2663 = ~n2661 & n2662 ;
  assign n2664 = n2660 ^ n2637 ^ n2549 ;
  assign n2665 = ( n2549 & n2637 ) | ( n2549 & n2660 ) | ( n2637 & n2660 ) ;
  assign n2666 = n26 & ~n2169 ;
  assign n2667 = n27 & ~n2174 ;
  assign n2668 = ( n26 & ~n2666 ) | ( n26 & n2667 ) | ( ~n2666 & n2667 ) ;
  assign n2669 = ( n2181 & n2235 ) | ( n2181 & n2667 ) | ( n2235 & n2667 ) ;
  assign n2670 = n2668 | n2669 ;
  assign n2671 = n2249 & ~n2648 ;
  assign n2672 = n2670 | n2671 ;
  assign n2673 = ( n2240 & ~n2663 ) | ( n2240 & n2670 ) | ( ~n2663 & n2670 ) ;
  assign n2674 = ( n2240 & n2663 ) | ( n2240 & n2672 ) | ( n2663 & n2672 ) ;
  assign n2675 = ~n2673 & n2674 ;
  assign n2676 = n27 & n2181 ;
  assign n2677 = n2656 ^ n2200 ^ n2181 ;
  assign n2678 = ( n2388 & ~n2659 ) | ( n2388 & n2675 ) | ( ~n2659 & n2675 ) ;
  assign n2679 = ~n2610 & n2678 ;
  assign n2680 = n2254 & n2677 ;
  assign n2681 = n2610 | n2678 ;
  assign n2682 = ~n2680 & n2681 ;
  assign n2683 = ( n2181 & n2200 ) | ( n2181 & n2656 ) | ( n2200 & n2656 ) ;
  assign n2684 = ( n26 & ~n2174 ) | ( n26 & n2676 ) | ( ~n2174 & n2676 ) ;
  assign n2685 = n2676 | n2684 ;
  assign n2686 = n2200 & ~n2235 ;
  assign n2687 = ( n2200 & n2685 ) | ( n2200 & ~n2686 ) | ( n2685 & ~n2686 ) ;
  assign n2688 = ~n2249 & n2677 ;
  assign n2689 = ( n2677 & n2687 ) | ( n2677 & ~n2688 ) | ( n2687 & ~n2688 ) ;
  assign n2690 = ( n2240 & ~n2682 ) | ( n2240 & n2687 ) | ( ~n2682 & n2687 ) ;
  assign n2691 = ( n2240 & n2682 ) | ( n2240 & n2689 ) | ( n2682 & n2689 ) ;
  assign n2692 = n2683 ^ n2217 ^ n2200 ;
  assign n2693 = n2254 & n2692 ;
  assign n2694 = ~n2690 & n2691 ;
  assign n2695 = n27 & n2200 ;
  assign n2696 = ( n2678 & ~n2679 ) | ( n2678 & n2694 ) | ( ~n2679 & n2694 ) ;
  assign n2697 = n26 & ~n2181 ;
  assign n2698 = ( n26 & n2695 ) | ( n26 & ~n2697 ) | ( n2695 & ~n2697 ) ;
  assign n2699 = ( n2217 & n2235 ) | ( n2217 & n2695 ) | ( n2235 & n2695 ) ;
  assign n2700 = n2635 | n2696 ;
  assign n2701 = ~n2635 & n2696 ;
  assign n2702 = n2698 | n2699 ;
  assign n2703 = ~n2693 & n2700 ;
  assign n2704 = ~n2249 & n2692 ;
  assign n2705 = ( n2692 & n2702 ) | ( n2692 & ~n2704 ) | ( n2702 & ~n2704 ) ;
  assign n2706 = ( n2240 & n2703 ) | ( n2240 & n2705 ) | ( n2703 & n2705 ) ;
  assign n2707 = ( n2240 & n2702 ) | ( n2240 & ~n2703 ) | ( n2702 & ~n2703 ) ;
  assign n2708 = n2706 & ~n2707 ;
  assign n2709 = ( n2696 & ~n2701 ) | ( n2696 & n2708 ) | ( ~n2701 & n2708 ) ;
  assign n2710 = n2169 & n2400 ;
  assign n2711 = ( ~n2174 & n2411 ) | ( ~n2174 & n2710 ) | ( n2411 & n2710 ) ;
  assign n2712 = n2710 | n2711 ;
  assign n2713 = n2181 & ~n2402 ;
  assign n2714 = ( n2181 & n2712 ) | ( n2181 & ~n2713 ) | ( n2712 & ~n2713 ) ;
  assign n2715 = n2412 & n2648 ;
  assign n2716 = ( n2412 & n2714 ) | ( n2412 & ~n2715 ) | ( n2714 & ~n2715 ) ;
  assign n2717 = n2716 ^ n40 ^ x11 ;
  assign n2718 = ( n2572 & n2638 ) | ( n2572 & n2717 ) | ( n2638 & n2717 ) ;
  assign n2719 = n2717 ^ n2638 ^ n2572 ;
  assign n2720 = n2181 & n2361 ;
  assign n2721 = ( ~n2174 & n2386 ) | ( ~n2174 & n2720 ) | ( n2386 & n2720 ) ;
  assign n2722 = n2720 | n2721 ;
  assign n2723 = n2200 & ~n2360 ;
  assign n2724 = ( n2200 & n2722 ) | ( n2200 & ~n2723 ) | ( n2722 & ~n2723 ) ;
  assign n2725 = n2461 & n2648 ;
  assign n2726 = n2357 & ~n2677 ;
  assign n2727 = ( n2357 & n2724 ) | ( n2357 & ~n2726 ) | ( n2724 & ~n2726 ) ;
  assign n2728 = n2727 ^ n1678 ^ x8 ;
  assign n2729 = ( n2584 & n2657 ) | ( n2584 & n2728 ) | ( n2657 & n2728 ) ;
  assign n2730 = n2728 ^ n2657 ^ n2584 ;
  assign n2731 = n2181 & n2386 ;
  assign n2732 = ( n2217 & n2360 ) | ( n2217 & n2731 ) | ( n2360 & n2731 ) ;
  assign n2733 = n2731 | n2732 ;
  assign n2734 = n2200 & ~n2361 ;
  assign n2735 = ( n2200 & n2733 ) | ( n2200 & ~n2734 ) | ( n2733 & ~n2734 ) ;
  assign n2736 = n2357 & ~n2692 ;
  assign n2737 = ( n2357 & n2735 ) | ( n2357 & ~n2736 ) | ( n2735 & ~n2736 ) ;
  assign n2738 = n2737 ^ n1678 ^ x8 ;
  assign n2739 = n2738 ^ n2729 ^ n2636 ;
  assign n2740 = ( n2636 & n2729 ) | ( n2636 & n2738 ) | ( n2729 & n2738 ) ;
  assign n2741 = n2169 & n2466 ;
  assign n2742 = ( ~n2174 & n2455 ) | ( ~n2174 & n2741 ) | ( n2455 & n2741 ) ;
  assign n2743 = n2741 | n2742 ;
  assign n2744 = n2181 & ~n2460 ;
  assign n2745 = ( n2181 & n2743 ) | ( n2181 & ~n2744 ) | ( n2743 & ~n2744 ) ;
  assign n2746 = n2181 & n2282 ;
  assign n2747 = ( n2461 & ~n2725 ) | ( n2461 & n2745 ) | ( ~n2725 & n2745 ) ;
  assign n2748 = ( ~n2174 & n2294 ) | ( ~n2174 & n2746 ) | ( n2294 & n2746 ) ;
  assign n2749 = n2746 | n2748 ;
  assign n2750 = n2200 & ~n2285 ;
  assign n2751 = ( n2200 & n2749 ) | ( n2200 & ~n2750 ) | ( n2749 & ~n2750 ) ;
  assign n2752 = ~n2288 & n2677 ;
  assign n2753 = ( n2677 & n2751 ) | ( n2677 & ~n2752 ) | ( n2751 & ~n2752 ) ;
  assign n2754 = n2753 ^ n1635 ^ x5 ;
  assign n2755 = n1654 & n2135 ;
  assign n2756 = n1654 & ~n2135 ;
  assign n2757 = n2756 ^ n2747 ^ n2626 ;
  assign n2758 = n2747 ^ n1654 ^ 1'b0 ;
  assign n2759 = ( n2626 & n2755 ) | ( n2626 & n2758 ) | ( n2755 & n2758 ) ;
  assign n2760 = n2181 & n2294 ;
  assign n2761 = ( n2217 & n2285 ) | ( n2217 & n2760 ) | ( n2285 & n2760 ) ;
  assign n2762 = n2760 | n2761 ;
  assign n2763 = n2754 ^ n2665 ^ n2567 ;
  assign n2764 = ( n2567 & n2665 ) | ( n2567 & n2754 ) | ( n2665 & n2754 ) ;
  assign n2765 = n2200 & ~n2282 ;
  assign n2766 = ( n2200 & n2762 ) | ( n2200 & ~n2765 ) | ( n2762 & ~n2765 ) ;
  assign n2767 = ~n2288 & n2692 ;
  assign n2768 = ( n2692 & n2766 ) | ( n2692 & ~n2767 ) | ( n2766 & ~n2767 ) ;
  assign n2769 = n2768 ^ n1635 ^ x5 ;
  assign n2770 = n2769 ^ n2764 ^ n2568 ;
  assign n2771 = ( n2568 & n2764 ) | ( n2568 & n2769 ) | ( n2764 & n2769 ) ;
  assign n2772 = n27 & n2217 ;
  assign n2773 = ( ~n2223 & n2235 ) | ( ~n2223 & n2772 ) | ( n2235 & n2772 ) ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = ( n2200 & n2217 ) | ( n2200 & n2683 ) | ( n2217 & n2683 ) ;
  assign n2776 = n2223 ^ n2217 ^ 1'b0 ;
  assign n2777 = n26 & ~n2200 ;
  assign n2778 = n2776 ^ n2775 ^ 1'b0 ;
  assign n2779 = ( n26 & n2774 ) | ( n26 & ~n2777 ) | ( n2774 & ~n2777 ) ;
  assign n2780 = n2249 & n2778 ;
  assign n2781 = ( n2249 & n2779 ) | ( n2249 & ~n2780 ) | ( n2779 & ~n2780 ) ;
  assign n2782 = n2181 & n2411 ;
  assign n2783 = n2781 ^ n2239 ^ x2 ;
  assign n2784 = ( n2664 & n2709 ) | ( n2664 & n2783 ) | ( n2709 & n2783 ) ;
  assign n2785 = ( ~n2174 & n2400 ) | ( ~n2174 & n2782 ) | ( n2400 & n2782 ) ;
  assign n2786 = n2782 | n2785 ;
  assign n2787 = n2200 & n2294 ;
  assign n2788 = ( ~n2223 & n2285 ) | ( ~n2223 & n2787 ) | ( n2285 & n2787 ) ;
  assign n2789 = n2787 | n2788 ;
  assign n2790 = n2217 & ~n2282 ;
  assign n2791 = ( n2217 & n2789 ) | ( n2217 & ~n2790 ) | ( n2789 & ~n2790 ) ;
  assign n2792 = n2778 & ~n2791 ;
  assign n2793 = ( n2288 & n2791 ) | ( n2288 & ~n2792 ) | ( n2791 & ~n2792 ) ;
  assign n2794 = n2200 & ~n2402 ;
  assign n2795 = ( n2200 & n2786 ) | ( n2200 & ~n2794 ) | ( n2786 & ~n2794 ) ;
  assign n2796 = n2412 & ~n2677 ;
  assign n2797 = ( n2412 & n2795 ) | ( n2412 & ~n2796 ) | ( n2795 & ~n2796 ) ;
  assign n2798 = n2797 ^ n40 ^ x11 ;
  assign n2799 = ( n2593 & n2718 ) | ( n2593 & n2798 ) | ( n2718 & n2798 ) ;
  assign n2800 = n2798 ^ n2718 ^ n2593 ;
  assign n2801 = n2217 & n2411 ;
  assign n2802 = n2223 & n2402 ;
  assign n2803 = ( n2402 & n2801 ) | ( n2402 & ~n2802 ) | ( n2801 & ~n2802 ) ;
  assign n2804 = ( n2200 & n2400 ) | ( n2200 & n2801 ) | ( n2400 & n2801 ) ;
  assign n2805 = n2803 | n2804 ;
  assign n2806 = n2412 & n2778 ;
  assign n2807 = ( n2412 & n2805 ) | ( n2412 & ~n2806 ) | ( n2805 & ~n2806 ) ;
  assign n2808 = n2793 ^ n1635 ^ x5 ;
  assign n2809 = ( n2658 & n2771 ) | ( n2658 & n2808 ) | ( n2771 & n2808 ) ;
  assign n2810 = n2808 ^ n2771 ^ n2658 ;
  assign n2811 = n2181 & n2400 ;
  assign n2812 = ( n2217 & n2402 ) | ( n2217 & n2811 ) | ( n2402 & n2811 ) ;
  assign n2813 = n2811 | n2812 ;
  assign n2814 = n2200 & ~n2411 ;
  assign n2815 = ( n2200 & n2813 ) | ( n2200 & ~n2814 ) | ( n2813 & ~n2814 ) ;
  assign n2816 = n2807 ^ n40 ^ x11 ;
  assign n2817 = n2412 & ~n2692 ;
  assign n2818 = ( n2217 & ~n2223 ) | ( n2217 & n2775 ) | ( ~n2223 & n2775 ) ;
  assign n2819 = ( n2412 & n2815 ) | ( n2412 & ~n2817 ) | ( n2815 & ~n2817 ) ;
  assign n2820 = n2819 ^ n40 ^ x11 ;
  assign n2821 = n2820 ^ n2799 ^ n2623 ;
  assign n2822 = ( n2623 & n2799 ) | ( n2623 & n2820 ) | ( n2799 & n2820 ) ;
  assign n2823 = n2822 ^ n2816 ^ n2757 ;
  assign n2824 = ( n2757 & n2816 ) | ( n2757 & n2822 ) | ( n2816 & n2822 ) ;
  assign n2825 = ~n2223 & n2282 ;
  assign n2826 = n2219 & ~n2285 ;
  assign n2827 = ( n2219 & n2825 ) | ( n2219 & ~n2826 ) | ( n2825 & ~n2826 ) ;
  assign n2828 = ( n2217 & n2294 ) | ( n2217 & n2825 ) | ( n2294 & n2825 ) ;
  assign n2829 = n2827 | n2828 ;
  assign n2830 = n2288 | n2829 ;
  assign n2831 = n2818 ^ n2223 ^ n2219 ;
  assign n2832 = ( n2829 & n2830 ) | ( n2829 & ~n2831 ) | ( n2830 & ~n2831 ) ;
  assign n2833 = n2832 ^ n1635 ^ x5 ;
  assign n2834 = n2833 ^ n2809 ^ n2730 ;
  assign n2835 = ( n2730 & n2809 ) | ( n2730 & n2833 ) | ( n2809 & n2833 ) ;
  assign n2836 = n26 & ~n2217 ;
  assign n2837 = n27 & ~n2223 ;
  assign n2838 = ( n26 & ~n2836 ) | ( n26 & n2837 ) | ( ~n2836 & n2837 ) ;
  assign n2839 = ( n2219 & n2235 ) | ( n2219 & n2837 ) | ( n2235 & n2837 ) ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = n2249 & n2831 ;
  assign n2842 = ( n2249 & n2840 ) | ( n2249 & ~n2841 ) | ( n2840 & ~n2841 ) ;
  assign n2843 = ( n2219 & ~n2223 ) | ( n2219 & n2818 ) | ( ~n2223 & n2818 ) ;
  assign n2844 = n2842 ^ n2239 ^ x2 ;
  assign n2845 = ( n2763 & n2784 ) | ( n2763 & n2844 ) | ( n2784 & n2844 ) ;
  assign n2846 = n27 & n2219 ;
  assign n2847 = ( n26 & ~n2223 ) | ( n26 & n2846 ) | ( ~n2223 & n2846 ) ;
  assign n2848 = n2846 | n2847 ;
  assign n2849 = n2220 & ~n2235 ;
  assign n2850 = n2843 ^ n2220 ^ n2219 ;
  assign n2851 = ( n2220 & n2848 ) | ( n2220 & ~n2849 ) | ( n2848 & ~n2849 ) ;
  assign n2852 = ~n2249 & n2850 ;
  assign n2853 = ( n2850 & n2851 ) | ( n2850 & ~n2852 ) | ( n2851 & ~n2852 ) ;
  assign n2854 = n2853 ^ n2239 ^ x2 ;
  assign n2855 = ( n2219 & n2220 ) | ( n2219 & n2843 ) | ( n2220 & n2843 ) ;
  assign n2856 = ( n2770 & n2845 ) | ( n2770 & n2854 ) | ( n2845 & n2854 ) ;
  assign n2857 = n27 & n2220 ;
  assign n2858 = n2855 ^ n2221 ^ n2220 ;
  assign n2859 = ( ~n2221 & n2235 ) | ( ~n2221 & n2857 ) | ( n2235 & n2857 ) ;
  assign n2860 = n2857 | n2859 ;
  assign n2861 = n26 & ~n2219 ;
  assign n2862 = ( n26 & n2860 ) | ( n26 & ~n2861 ) | ( n2860 & ~n2861 ) ;
  assign n2863 = n2858 & ~n2862 ;
  assign n2864 = ( n2249 & n2862 ) | ( n2249 & ~n2863 ) | ( n2862 & ~n2863 ) ;
  assign n2865 = n2864 ^ n2239 ^ x2 ;
  assign n2866 = n2865 ^ n2856 ^ n2810 ;
  assign n2867 = ( n2220 & ~n2221 ) | ( n2220 & n2855 ) | ( ~n2221 & n2855 ) ;
  assign n2868 = n1530 & n2866 ;
  assign n2869 = ~n2222 & n2235 ;
  assign n2870 = ( n2810 & n2856 ) | ( n2810 & n2865 ) | ( n2856 & n2865 ) ;
  assign n2871 = n27 & ~n2221 ;
  assign n2872 = ( n26 & n2220 ) | ( n26 & n2871 ) | ( n2220 & n2871 ) ;
  assign n2873 = n2871 | n2872 ;
  assign n2874 = ( n2235 & ~n2869 ) | ( n2235 & n2873 ) | ( ~n2869 & n2873 ) ;
  assign n2875 = n2867 ^ n2222 ^ n2221 ;
  assign n2876 = n2249 | n2874 ;
  assign n2877 = ( n2874 & ~n2875 ) | ( n2874 & n2876 ) | ( ~n2875 & n2876 ) ;
  assign n2878 = n2877 ^ n2239 ^ x2 ;
  assign n2879 = n2878 ^ n2870 ^ n2834 ;
  assign n2880 = ( n2834 & n2870 ) | ( n2834 & n2878 ) | ( n2870 & n2878 ) ;
  assign n2881 = ( n748 & n2868 ) | ( n748 & n2879 ) | ( n2868 & n2879 ) ;
  assign n2882 = n2219 & n2282 ;
  assign n2883 = ( ~n2223 & n2294 ) | ( ~n2223 & n2882 ) | ( n2294 & n2882 ) ;
  assign n2884 = ( ~n2221 & n2222 ) | ( ~n2221 & n2867 ) | ( n2222 & n2867 ) ;
  assign n2885 = n2288 & ~n2850 ;
  assign n2886 = n2882 | n2883 ;
  assign n2887 = n2220 & ~n2285 ;
  assign n2888 = ( n2220 & n2886 ) | ( n2220 & ~n2887 ) | ( n2886 & ~n2887 ) ;
  assign n2889 = ( n2288 & ~n2885 ) | ( n2288 & n2888 ) | ( ~n2885 & n2888 ) ;
  assign n2890 = n2889 ^ n1635 ^ x5 ;
  assign n2891 = n2890 ^ n2835 ^ n2739 ;
  assign n2892 = ( n2739 & n2835 ) | ( n2739 & n2890 ) | ( n2835 & n2890 ) ;
  assign n2893 = n2884 ^ n2222 ^ n2216 ;
  assign n2894 = n27 & n2222 ;
  assign n2895 = ( n26 & ~n2221 ) | ( n26 & n2894 ) | ( ~n2221 & n2894 ) ;
  assign n2896 = n2894 | n2895 ;
  assign n2897 = ~n2216 & n2235 ;
  assign n2898 = ( n2235 & n2896 ) | ( n2235 & ~n2897 ) | ( n2896 & ~n2897 ) ;
  assign n2899 = ~n2249 & n2893 ;
  assign n2900 = ( n2893 & n2898 ) | ( n2893 & ~n2899 ) | ( n2898 & ~n2899 ) ;
  assign n2901 = n2900 ^ n2239 ^ x2 ;
  assign n2902 = n2901 ^ n2891 ^ n2880 ;
  assign n2903 = ( n2880 & n2891 ) | ( n2880 & n2901 ) | ( n2891 & n2901 ) ;
  assign n2904 = ( n1421 & n2881 ) | ( n1421 & n2902 ) | ( n2881 & n2902 ) ;
  assign n2905 = n2357 & n2831 ;
  assign n2906 = n2902 ^ n2881 ^ n1421 ;
  assign n2907 = n2223 & n2360 ;
  assign n2908 = n2217 & n2361 ;
  assign n2909 = ( n2360 & ~n2907 ) | ( n2360 & n2908 ) | ( ~n2907 & n2908 ) ;
  assign n2910 = ( n2200 & n2386 ) | ( n2200 & n2908 ) | ( n2386 & n2908 ) ;
  assign n2911 = n2909 | n2910 ;
  assign n2912 = n2357 & n2778 ;
  assign n2913 = ( n2357 & n2911 ) | ( n2357 & ~n2912 ) | ( n2911 & ~n2912 ) ;
  assign n2914 = n2913 ^ n1678 ^ x8 ;
  assign n2915 = n2914 ^ n2740 ^ n2719 ;
  assign n2916 = ( n2719 & n2740 ) | ( n2719 & n2914 ) | ( n2740 & n2914 ) ;
  assign n2917 = ~n2223 & n2361 ;
  assign n2918 = n2219 & ~n2360 ;
  assign n2919 = ( n2219 & n2917 ) | ( n2219 & ~n2918 ) | ( n2917 & ~n2918 ) ;
  assign n2920 = ( n2217 & n2386 ) | ( n2217 & n2917 ) | ( n2386 & n2917 ) ;
  assign n2921 = n2919 | n2920 ;
  assign n2922 = ( n2357 & ~n2905 ) | ( n2357 & n2921 ) | ( ~n2905 & n2921 ) ;
  assign n2923 = n2922 ^ n1678 ^ x8 ;
  assign n2924 = ( n2800 & n2916 ) | ( n2800 & n2923 ) | ( n2916 & n2923 ) ;
  assign n2925 = n2923 ^ n2916 ^ n2800 ;
  assign n2926 = n2220 & n2282 ;
  assign n2927 = n2221 & n2285 ;
  assign n2928 = ( n2285 & n2926 ) | ( n2285 & ~n2927 ) | ( n2926 & ~n2927 ) ;
  assign n2929 = n2288 & n2858 ;
  assign n2930 = ( n2219 & n2294 ) | ( n2219 & n2926 ) | ( n2294 & n2926 ) ;
  assign n2931 = n2928 | n2930 ;
  assign n2932 = ( n2288 & ~n2929 ) | ( n2288 & n2931 ) | ( ~n2929 & n2931 ) ;
  assign n2933 = n2932 ^ n1635 ^ x5 ;
  assign n2934 = n2933 ^ n2915 ^ n2892 ;
  assign n2935 = ( n2892 & n2915 ) | ( n2892 & n2933 ) | ( n2915 & n2933 ) ;
  assign n2936 = n2357 & ~n2850 ;
  assign n2937 = n2219 & n2361 ;
  assign n2938 = ( ~n2223 & n2386 ) | ( ~n2223 & n2937 ) | ( n2386 & n2937 ) ;
  assign n2939 = n2937 | n2938 ;
  assign n2940 = n2220 & ~n2360 ;
  assign n2941 = ( n2220 & n2939 ) | ( n2220 & ~n2940 ) | ( n2939 & ~n2940 ) ;
  assign n2942 = ( n2357 & ~n2936 ) | ( n2357 & n2941 ) | ( ~n2936 & n2941 ) ;
  assign n2943 = n2942 ^ n1678 ^ x8 ;
  assign n2944 = n2943 ^ n2924 ^ n2821 ;
  assign n2945 = ( n2821 & n2924 ) | ( n2821 & n2943 ) | ( n2924 & n2943 ) ;
  assign n2946 = n26 & ~n2222 ;
  assign n2947 = n27 & n2216 ;
  assign n2948 = ( n2216 & n2222 ) | ( n2216 & n2884 ) | ( n2222 & n2884 ) ;
  assign n2949 = ( ~n2224 & n2235 ) | ( ~n2224 & n2947 ) | ( n2235 & n2947 ) ;
  assign n2950 = n2947 | n2949 ;
  assign n2951 = ( n26 & ~n2946 ) | ( n26 & n2950 ) | ( ~n2946 & n2950 ) ;
  assign n2952 = ~n2222 & n2285 ;
  assign n2953 = ~n2221 & n2282 ;
  assign n2954 = ( n2285 & ~n2952 ) | ( n2285 & n2953 ) | ( ~n2952 & n2953 ) ;
  assign n2955 = n2288 & ~n2875 ;
  assign n2956 = ( n2220 & n2294 ) | ( n2220 & n2953 ) | ( n2294 & n2953 ) ;
  assign n2957 = ( n2954 & ~n2955 ) | ( n2954 & n2956 ) | ( ~n2955 & n2956 ) ;
  assign n2958 = n2955 | n2957 ;
  assign n2959 = n2958 ^ n1635 ^ x5 ;
  assign n2960 = ( n2925 & n2935 ) | ( n2925 & n2959 ) | ( n2935 & n2959 ) ;
  assign n2961 = n2959 ^ n2935 ^ n2925 ;
  assign n2962 = n2224 ^ n2216 ^ 1'b0 ;
  assign n2963 = n2962 ^ n2948 ^ 1'b0 ;
  assign n2964 = ~n2951 & n2963 ;
  assign n2965 = ( n2249 & n2951 ) | ( n2249 & ~n2964 ) | ( n2951 & ~n2964 ) ;
  assign n2966 = n2965 ^ n2239 ^ x2 ;
  assign n2967 = n2966 ^ n2934 ^ n2903 ;
  assign n2968 = ( n2903 & n2934 ) | ( n2903 & n2966 ) | ( n2934 & n2966 ) ;
  assign n2969 = n2222 & n2282 ;
  assign n2970 = ( ~n2221 & n2294 ) | ( ~n2221 & n2969 ) | ( n2294 & n2969 ) ;
  assign n2971 = n2969 | n2970 ;
  assign n2972 = ~n2216 & n2285 ;
  assign n2973 = ( n2285 & n2971 ) | ( n2285 & ~n2972 ) | ( n2971 & ~n2972 ) ;
  assign n2974 = n2288 & ~n2893 ;
  assign n2975 = ( n2288 & n2973 ) | ( n2288 & ~n2974 ) | ( n2973 & ~n2974 ) ;
  assign n2976 = ( n1557 & n2904 ) | ( n1557 & n2967 ) | ( n2904 & n2967 ) ;
  assign n2977 = n2967 ^ n2904 ^ n1557 ;
  assign n2978 = n2975 ^ n1635 ^ x5 ;
  assign n2979 = ( n2216 & ~n2224 ) | ( n2216 & n2948 ) | ( ~n2224 & n2948 ) ;
  assign n2980 = n2978 ^ n2960 ^ n2944 ;
  assign n2981 = ( n2944 & n2960 ) | ( n2944 & n2978 ) | ( n2960 & n2978 ) ;
  assign n2982 = ~n1620 & n2235 ;
  assign n2983 = n27 & ~n2224 ;
  assign n2984 = ( n1620 & n2224 ) | ( n1620 & n2979 ) | ( n2224 & n2979 ) ;
  assign n2985 = n2982 | n2983 ;
  assign n2986 = ( n1620 & n2224 ) | ( n1620 & ~n2979 ) | ( n2224 & ~n2979 ) ;
  assign n2987 = n2986 ^ n2984 ^ n2979 ;
  assign n2988 = ( n26 & n2216 ) | ( n26 & n2983 ) | ( n2216 & n2983 ) ;
  assign n2989 = n2985 | n2988 ;
  assign n2990 = ~n2249 & n2987 ;
  assign n2991 = ( n2987 & n2989 ) | ( n2987 & ~n2990 ) | ( n2989 & ~n2990 ) ;
  assign n2992 = n2991 ^ n2239 ^ x2 ;
  assign n2993 = n2992 ^ n2968 ^ n2961 ;
  assign n2994 = ( n2961 & n2968 ) | ( n2961 & n2992 ) | ( n2968 & n2992 ) ;
  assign n2995 = ( n1617 & n2976 ) | ( n1617 & n2993 ) | ( n2976 & n2993 ) ;
  assign n2996 = n2993 ^ n2976 ^ n1617 ;
  assign n2997 = n2984 ^ n2224 ^ 1'b0 ;
  assign n2998 = ~n2249 & n2997 ;
  assign n2999 = n27 & ~n1620 ;
  assign n3000 = ( n26 & ~n2224 ) | ( n26 & n2999 ) | ( ~n2224 & n2999 ) ;
  assign n3001 = ( n2997 & ~n2998 ) | ( n2997 & n2999 ) | ( ~n2998 & n2999 ) ;
  assign n3002 = n3000 | n3001 ;
  assign n3003 = n3002 ^ n2239 ^ x2 ;
  assign n3004 = n3003 ^ n2994 ^ n2980 ;
  assign n3005 = n1620 | n2986 ;
  assign n3006 = ( n2980 & n2994 ) | ( n2980 & n3003 ) | ( n2994 & n3003 ) ;
  assign n3007 = ( n1625 & n2995 ) | ( n1625 & n3004 ) | ( n2995 & n3004 ) ;
  assign n3008 = n3004 ^ n2995 ^ n1625 ;
  assign n3009 = n2249 & ~n3005 ;
  assign n3010 = n2461 & n2778 ;
  assign n3011 = n2216 & n2282 ;
  assign n3012 = n26 & ~n1620 ;
  assign n3013 = n3009 | n3012 ;
  assign n3014 = ~n2224 & n2285 ;
  assign n3015 = n3011 | n3014 ;
  assign n3016 = ~n1620 & n2285 ;
  assign n3017 = ( n2222 & n2294 ) | ( n2222 & n3011 ) | ( n2294 & n3011 ) ;
  assign n3018 = n3013 ^ n2239 ^ x2 ;
  assign n3019 = n2461 & ~n2692 ;
  assign n3020 = ~n2224 & n2282 ;
  assign n3021 = n3016 | n3020 ;
  assign n3022 = ( n2216 & n2294 ) | ( n2216 & n3020 ) | ( n2294 & n3020 ) ;
  assign n3023 = n3021 | n3022 ;
  assign n3024 = n2288 & ~n2987 ;
  assign n3025 = ( n2288 & n3023 ) | ( n2288 & ~n3024 ) | ( n3023 & ~n3024 ) ;
  assign n3026 = n2288 & ~n2963 ;
  assign n3027 = ( n3015 & n3017 ) | ( n3015 & ~n3026 ) | ( n3017 & ~n3026 ) ;
  assign n3028 = n2288 & n2997 ;
  assign n3029 = ~n1620 & n2282 ;
  assign n3030 = n3028 | n3029 ;
  assign n3031 = ( ~n2224 & n2294 ) | ( ~n2224 & n3028 ) | ( n2294 & n3028 ) ;
  assign n3032 = n3030 | n3031 ;
  assign n3033 = n2220 & n2361 ;
  assign n3034 = n3026 | n3027 ;
  assign n3035 = n2221 & n2360 ;
  assign n3036 = ( n2360 & n3033 ) | ( n2360 & ~n3035 ) | ( n3033 & ~n3035 ) ;
  assign n3037 = ( n2219 & n2386 ) | ( n2219 & n3033 ) | ( n2386 & n3033 ) ;
  assign n3038 = n3036 | n3037 ;
  assign n3039 = n2357 & n2858 ;
  assign n3040 = ( n2357 & n3038 ) | ( n2357 & ~n3039 ) | ( n3038 & ~n3039 ) ;
  assign n3041 = n3040 ^ n1678 ^ x8 ;
  assign n3042 = ( n2823 & n2945 ) | ( n2823 & n3041 ) | ( n2945 & n3041 ) ;
  assign n3043 = n3025 ^ n1635 ^ x5 ;
  assign n3044 = n3034 ^ n1635 ^ x5 ;
  assign n3045 = ~n1620 & n2294 ;
  assign n3046 = n3032 ^ n1635 ^ x5 ;
  assign n3047 = n2288 & ~n3005 ;
  assign n3048 = n3045 | n3047 ;
  assign n3049 = n3048 ^ n1635 ^ x5 ;
  assign n3050 = n3041 ^ n2945 ^ n2823 ;
  assign n3051 = n3050 ^ n3044 ^ n3018 ;
  assign n3052 = n3051 ^ n3006 ^ n2981 ;
  assign n3053 = ( n530 & n3007 ) | ( n530 & n3052 ) | ( n3007 & n3052 ) ;
  assign n3054 = ( n2981 & n3006 ) | ( n2981 & n3051 ) | ( n3006 & n3051 ) ;
  assign n3055 = ( n3018 & n3044 ) | ( n3018 & n3050 ) | ( n3044 & n3050 ) ;
  assign n3056 = n3052 ^ n3007 ^ n530 ;
  assign n3057 = n2181 & n2455 ;
  assign n3058 = ( ~n2174 & n2466 ) | ( ~n2174 & n3057 ) | ( n2466 & n3057 ) ;
  assign n3059 = n3057 | n3058 ;
  assign n3060 = n2461 & ~n2677 ;
  assign n3061 = n2200 & ~n2460 ;
  assign n3062 = ( n2200 & n3059 ) | ( n2200 & ~n3061 ) | ( n3059 & ~n3061 ) ;
  assign n3063 = ( n2461 & ~n3060 ) | ( n2461 & n3062 ) | ( ~n3060 & n3062 ) ;
  assign n3064 = ~n2223 & n2411 ;
  assign n3065 = n2219 & ~n2402 ;
  assign n3066 = ( n2219 & n3064 ) | ( n2219 & ~n3065 ) | ( n3064 & ~n3065 ) ;
  assign n3067 = ( n2217 & n2400 ) | ( n2217 & n3064 ) | ( n2400 & n3064 ) ;
  assign n3068 = n3066 | n3067 ;
  assign n3069 = n2412 & n2831 ;
  assign n3070 = ( n2412 & n3068 ) | ( n2412 & ~n3069 ) | ( n3068 & ~n3069 ) ;
  assign n3071 = n1654 & n2169 ;
  assign n3072 = n3063 ^ n82 ^ x14 ;
  assign n3073 = n3072 ^ n3071 ^ n2240 ;
  assign n3074 = ( n2240 & n3071 ) | ( n2240 & n3072 ) | ( n3071 & n3072 ) ;
  assign n3075 = n1654 & ~n2174 ;
  assign n3076 = n3070 ^ n40 ^ x11 ;
  assign n3077 = n3076 ^ n3073 ^ n2759 ;
  assign n3078 = ( n2759 & n3073 ) | ( n2759 & n3076 ) | ( n3073 & n3076 ) ;
  assign n3079 = n1654 & n2181 ;
  assign n3080 = ( n2240 & n3074 ) | ( n2240 & n3075 ) | ( n3074 & n3075 ) ;
  assign n3081 = n3075 ^ n3074 ^ n2240 ;
  assign n3082 = n2217 & ~n2460 ;
  assign n3083 = n2181 & n2466 ;
  assign n3084 = ( n2217 & ~n3082 ) | ( n2217 & n3083 ) | ( ~n3082 & n3083 ) ;
  assign n3085 = ( n2200 & n2455 ) | ( n2200 & n3083 ) | ( n2455 & n3083 ) ;
  assign n3086 = n3084 | n3085 ;
  assign n3087 = ( n2461 & ~n3019 ) | ( n2461 & n3086 ) | ( ~n3019 & n3086 ) ;
  assign n3088 = ~n2223 & n2460 ;
  assign n3089 = n2217 & ~n2455 ;
  assign n3090 = ( n2217 & n3088 ) | ( n2217 & ~n3089 ) | ( n3088 & ~n3089 ) ;
  assign n3091 = ( n2200 & n2466 ) | ( n2200 & n3088 ) | ( n2466 & n3088 ) ;
  assign n3092 = n3090 | n3091 ;
  assign n3093 = ( n2461 & ~n3010 ) | ( n2461 & n3092 ) | ( ~n3010 & n3092 ) ;
  assign n3094 = n1654 & n2200 ;
  assign n3095 = ( n1636 & n2240 ) | ( n1636 & ~n3094 ) | ( n2240 & ~n3094 ) ;
  assign n3096 = n3080 ^ n3079 ^ n2240 ;
  assign n3097 = n3094 ^ n2240 ^ n1636 ;
  assign n3098 = ~n2221 & n2361 ;
  assign n3099 = ( n2240 & n3079 ) | ( n2240 & n3080 ) | ( n3079 & n3080 ) ;
  assign n3100 = ~n2222 & n2360 ;
  assign n3101 = ( n2360 & n3098 ) | ( n2360 & ~n3100 ) | ( n3098 & ~n3100 ) ;
  assign n3102 = n2357 & ~n2875 ;
  assign n3103 = ( n2220 & n2386 ) | ( n2220 & n3098 ) | ( n2386 & n3098 ) ;
  assign n3104 = ( n3101 & ~n3102 ) | ( n3101 & n3103 ) | ( ~n3102 & n3103 ) ;
  assign n3105 = n3102 | n3104 ;
  assign n3106 = n3105 ^ n1678 ^ x8 ;
  assign n3107 = n3106 ^ n3077 ^ n2824 ;
  assign n3108 = n3107 ^ n3043 ^ n3042 ;
  assign n3109 = ( n2824 & n3077 ) | ( n2824 & n3106 ) | ( n3077 & n3106 ) ;
  assign n3110 = ( n3042 & n3043 ) | ( n3042 & n3107 ) | ( n3043 & n3107 ) ;
  assign n3111 = n3108 ^ n3055 ^ n3054 ;
  assign n3112 = ( n1548 & n3053 ) | ( n1548 & n3111 ) | ( n3053 & n3111 ) ;
  assign n3113 = ( n3054 & n3055 ) | ( n3054 & n3108 ) | ( n3055 & n3108 ) ;
  assign n3114 = n3111 ^ n3053 ^ n1548 ;
  assign n3115 = n2219 & n2411 ;
  assign n3116 = ( ~n2223 & n2400 ) | ( ~n2223 & n3115 ) | ( n2400 & n3115 ) ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = n2220 & ~n2402 ;
  assign n3119 = ( n2220 & n3117 ) | ( n2220 & ~n3118 ) | ( n3117 & ~n3118 ) ;
  assign n3120 = n3087 ^ n82 ^ x14 ;
  assign n3121 = n2412 & ~n2850 ;
  assign n3122 = ( n2412 & n3119 ) | ( n2412 & ~n3121 ) | ( n3119 & ~n3121 ) ;
  assign n3123 = n3122 ^ n40 ^ x11 ;
  assign n3124 = n3123 ^ n3120 ^ n3081 ;
  assign n3125 = ( n3081 & n3120 ) | ( n3081 & n3123 ) | ( n3120 & n3123 ) ;
  assign n3126 = n2222 & n2361 ;
  assign n3127 = ( ~n2221 & n2386 ) | ( ~n2221 & n3126 ) | ( n2386 & n3126 ) ;
  assign n3128 = n3126 | n3127 ;
  assign n3129 = ~n2216 & n2360 ;
  assign n3130 = ( n2360 & n3128 ) | ( n2360 & ~n3129 ) | ( n3128 & ~n3129 ) ;
  assign n3131 = n2357 & ~n2893 ;
  assign n3132 = ( n2357 & n3130 ) | ( n2357 & ~n3131 ) | ( n3130 & ~n3131 ) ;
  assign n3133 = n3132 ^ n1678 ^ x8 ;
  assign n3134 = n3133 ^ n3124 ^ n3078 ;
  assign n3135 = ( n3078 & n3124 ) | ( n3078 & n3133 ) | ( n3124 & n3133 ) ;
  assign n3136 = n3134 ^ n3109 ^ n3046 ;
  assign n3137 = n3136 ^ n3113 ^ n3110 ;
  assign n3138 = ( n3110 & n3113 ) | ( n3110 & n3136 ) | ( n3113 & n3136 ) ;
  assign n3139 = n2221 & n2402 ;
  assign n3140 = n2220 & n2411 ;
  assign n3141 = ( n2402 & ~n3139 ) | ( n2402 & n3140 ) | ( ~n3139 & n3140 ) ;
  assign n3142 = ( n2219 & n2400 ) | ( n2219 & n3140 ) | ( n2400 & n3140 ) ;
  assign n3143 = n3141 | n3142 ;
  assign n3144 = n2412 & n2858 ;
  assign n3145 = ( n2412 & n3143 ) | ( n2412 & ~n3144 ) | ( n3143 & ~n3144 ) ;
  assign n3146 = ( n1626 & n3112 ) | ( n1626 & n3137 ) | ( n3112 & n3137 ) ;
  assign n3147 = n3145 ^ n40 ^ x11 ;
  assign n3148 = ( n3046 & n3109 ) | ( n3046 & n3134 ) | ( n3109 & n3134 ) ;
  assign n3149 = n3093 ^ n82 ^ x14 ;
  assign n3150 = ( n3096 & n3147 ) | ( n3096 & n3149 ) | ( n3147 & n3149 ) ;
  assign n3151 = ~n2224 & n2360 ;
  assign n3152 = ~n1620 & n2360 ;
  assign n3153 = n3137 ^ n3112 ^ n1626 ;
  assign n3154 = n3149 ^ n3147 ^ n3096 ;
  assign n3155 = n2357 & ~n2963 ;
  assign n3156 = n2216 & n2361 ;
  assign n3157 = n3151 | n3156 ;
  assign n3158 = ( n2222 & n2386 ) | ( n2222 & n3156 ) | ( n2386 & n3156 ) ;
  assign n3159 = ( ~n3155 & n3157 ) | ( ~n3155 & n3158 ) | ( n3157 & n3158 ) ;
  assign n3160 = n3155 | n3159 ;
  assign n3161 = n3160 ^ n1678 ^ x8 ;
  assign n3162 = ( n3125 & n3154 ) | ( n3125 & n3161 ) | ( n3154 & n3161 ) ;
  assign n3163 = n3161 ^ n3154 ^ n3125 ;
  assign n3164 = n3163 ^ n3135 ^ n3049 ;
  assign n3165 = n3164 ^ n3148 ^ n3138 ;
  assign n3166 = ( n3138 & n3148 ) | ( n3138 & n3164 ) | ( n3148 & n3164 ) ;
  assign n3167 = ( n3049 & n3135 ) | ( n3049 & n3163 ) | ( n3135 & n3163 ) ;
  assign n3168 = ~n1620 & n2361 ;
  assign n3169 = ~n2224 & n2361 ;
  assign n3170 = n3152 | n3169 ;
  assign n3171 = ( n2216 & n2386 ) | ( n2216 & n3169 ) | ( n2386 & n3169 ) ;
  assign n3172 = n3170 | n3171 ;
  assign n3173 = n2357 & ~n2987 ;
  assign n3174 = ( n2357 & n3172 ) | ( n2357 & ~n3173 ) | ( n3172 & ~n3173 ) ;
  assign n3175 = n2357 & n2997 ;
  assign n3176 = n3168 | n3175 ;
  assign n3177 = ( ~n2224 & n2386 ) | ( ~n2224 & n3175 ) | ( n2386 & n3175 ) ;
  assign n3178 = n3176 | n3177 ;
  assign n3179 = n2223 & n2455 ;
  assign n3180 = n2461 & n2831 ;
  assign n3181 = ~n1620 & n2386 ;
  assign n3182 = n3178 ^ n1678 ^ x8 ;
  assign n3183 = n2357 & ~n3005 ;
  assign n3184 = n3181 | n3183 ;
  assign n3185 = ( n1554 & n3146 ) | ( n1554 & n3165 ) | ( n3146 & n3165 ) ;
  assign n3186 = n3174 ^ n1678 ^ x8 ;
  assign n3187 = n3184 ^ n1678 ^ x8 ;
  assign n3188 = n2220 & n2400 ;
  assign n3189 = n3165 ^ n3146 ^ n1554 ;
  assign n3190 = n2412 & ~n2875 ;
  assign n3191 = n2221 & n2411 ;
  assign n3192 = ( n2411 & n3188 ) | ( n2411 & ~n3191 ) | ( n3188 & ~n3191 ) ;
  assign n3193 = ( n2222 & n2402 ) | ( n2222 & n3188 ) | ( n2402 & n3188 ) ;
  assign n3194 = ( ~n3190 & n3192 ) | ( ~n3190 & n3193 ) | ( n3192 & n3193 ) ;
  assign n3195 = n3190 | n3194 ;
  assign n3196 = n3195 ^ n40 ^ x11 ;
  assign n3197 = n2219 & n2460 ;
  assign n3198 = ( n2455 & ~n3179 ) | ( n2455 & n3197 ) | ( ~n3179 & n3197 ) ;
  assign n3199 = ( n2217 & n2466 ) | ( n2217 & n3197 ) | ( n2466 & n3197 ) ;
  assign n3200 = n3198 | n3199 ;
  assign n3201 = ( n2461 & ~n3180 ) | ( n2461 & n3200 ) | ( ~n3180 & n3200 ) ;
  assign n3202 = n3201 ^ n82 ^ x14 ;
  assign n3203 = n3202 ^ n3099 ^ n3097 ;
  assign n3204 = ( n3097 & n3099 ) | ( n3097 & n3202 ) | ( n3099 & n3202 ) ;
  assign n3205 = n3203 ^ n3196 ^ n3150 ;
  assign n3206 = ( n3150 & n3196 ) | ( n3150 & n3203 ) | ( n3196 & n3203 ) ;
  assign n3207 = ( n3162 & n3186 ) | ( n3162 & n3205 ) | ( n3186 & n3205 ) ;
  assign n3208 = n3205 ^ n3186 ^ n3162 ;
  assign n3209 = ( n3166 & n3167 ) | ( n3166 & n3208 ) | ( n3167 & n3208 ) ;
  assign n3210 = n3208 ^ n3167 ^ n3166 ;
  assign n3211 = ( n1627 & n3185 ) | ( n1627 & n3210 ) | ( n3185 & n3210 ) ;
  assign n3212 = n3210 ^ n3185 ^ n1627 ;
  assign n3213 = ~n2221 & n2460 ;
  assign n3214 = n2220 & ~n2455 ;
  assign n3215 = ( n2220 & n3213 ) | ( n2220 & ~n3214 ) | ( n3213 & ~n3214 ) ;
  assign n3216 = ( n2219 & n2466 ) | ( n2219 & n3213 ) | ( n2466 & n3213 ) ;
  assign n3217 = n3215 | n3216 ;
  assign n3218 = n2461 & n2858 ;
  assign n3219 = ( n2461 & n3217 ) | ( n2461 & ~n3218 ) | ( n3217 & ~n3218 ) ;
  assign n3220 = n2220 & n2460 ;
  assign n3221 = ( ~n2223 & n2466 ) | ( ~n2223 & n3220 ) | ( n2466 & n3220 ) ;
  assign n3222 = n3220 | n3221 ;
  assign n3223 = n2219 & ~n2455 ;
  assign n3224 = ( n2219 & n3222 ) | ( n2219 & ~n3223 ) | ( n3222 & ~n3223 ) ;
  assign n3225 = n2461 & ~n2850 ;
  assign n3226 = ( n2217 & ~n2223 ) | ( n2217 & n3219 ) | ( ~n2223 & n3219 ) ;
  assign n3227 = n3219 ^ n1654 ^ 1'b0 ;
  assign n3228 = ( ~n2217 & n3226 ) | ( ~n2217 & n3227 ) | ( n3226 & n3227 ) ;
  assign n3229 = n1654 & n2219 ;
  assign n3230 = n1654 & n2217 ;
  assign n3231 = ( n2461 & n3224 ) | ( n2461 & ~n3225 ) | ( n3224 & ~n3225 ) ;
  assign n3232 = n1654 & n2776 ;
  assign n3233 = n3232 ^ n3219 ^ 1'b0 ;
  assign n3234 = n3230 ^ n3229 ^ n1695 ;
  assign n3235 = n2216 & n2411 ;
  assign n3236 = ( ~n1695 & n3229 ) | ( ~n1695 & n3230 ) | ( n3229 & n3230 ) ;
  assign n3237 = ( n2222 & n2400 ) | ( n2222 & n3235 ) | ( n2400 & n3235 ) ;
  assign n3238 = n3231 ^ n82 ^ x14 ;
  assign n3239 = n3238 ^ n3230 ^ n3095 ;
  assign n3240 = ( n3095 & n3230 ) | ( n3095 & ~n3238 ) | ( n3230 & ~n3238 ) ;
  assign n3241 = n2222 & n2411 ;
  assign n3242 = ( ~n2221 & n2400 ) | ( ~n2221 & n3241 ) | ( n2400 & n3241 ) ;
  assign n3243 = n3241 | n3242 ;
  assign n3244 = ~n2216 & n2402 ;
  assign n3245 = ( n2402 & n3243 ) | ( n2402 & ~n3244 ) | ( n3243 & ~n3244 ) ;
  assign n3246 = ~n2224 & n2402 ;
  assign n3247 = n3235 | n3246 ;
  assign n3248 = n2412 & ~n2893 ;
  assign n3249 = ( n2412 & n3245 ) | ( n2412 & ~n3248 ) | ( n3245 & ~n3248 ) ;
  assign n3250 = n2412 & ~n2963 ;
  assign n3251 = ( n3237 & n3247 ) | ( n3237 & ~n3250 ) | ( n3247 & ~n3250 ) ;
  assign n3252 = n3250 | n3251 ;
  assign n3253 = n3252 ^ n40 ^ x11 ;
  assign n3254 = n3249 ^ n40 ^ x11 ;
  assign n3255 = n3253 ^ n3240 ^ n3233 ;
  assign n3256 = n3254 ^ n3239 ^ n3204 ;
  assign n3257 = ( n3204 & n3239 ) | ( n3204 & n3254 ) | ( n3239 & n3254 ) ;
  assign n3258 = n3256 ^ n3206 ^ n3182 ;
  assign n3259 = ( n3207 & n3209 ) | ( n3207 & n3258 ) | ( n3209 & n3258 ) ;
  assign n3260 = n3258 ^ n3209 ^ n3207 ;
  assign n3261 = ( n3187 & n3255 ) | ( n3187 & n3257 ) | ( n3255 & n3257 ) ;
  assign n3262 = ( n3182 & n3206 ) | ( n3182 & n3256 ) | ( n3206 & n3256 ) ;
  assign n3263 = ( n3233 & n3240 ) | ( n3233 & ~n3253 ) | ( n3240 & ~n3253 ) ;
  assign n3264 = n3260 ^ n3211 ^ n1587 ;
  assign n3265 = n3257 ^ n3255 ^ n3187 ;
  assign n3266 = n3265 ^ n3262 ^ n3259 ;
  assign n3267 = ( n3259 & n3262 ) | ( n3259 & n3265 ) | ( n3262 & n3265 ) ;
  assign n3268 = ( n1587 & n3211 ) | ( n1587 & n3260 ) | ( n3211 & n3260 ) ;
  assign n3269 = n3268 ^ n3266 ^ n1502 ;
  assign n3270 = ( n1502 & n3266 ) | ( n1502 & n3268 ) | ( n3266 & n3268 ) ;
  assign n3271 = ~n2224 & n2411 ;
  assign n3272 = ~n1620 & n2402 ;
  assign n3273 = n3271 | n3272 ;
  assign n3274 = ( n2216 & n2400 ) | ( n2216 & n3271 ) | ( n2400 & n3271 ) ;
  assign n3275 = n3273 | n3274 ;
  assign n3276 = ~n1620 & n2411 ;
  assign n3277 = n2412 & n2997 ;
  assign n3278 = n3276 | n3277 ;
  assign n3279 = ( ~n2224 & n2400 ) | ( ~n2224 & n3277 ) | ( n2400 & n3277 ) ;
  assign n3280 = n3278 | n3279 ;
  assign n3281 = n3280 ^ n40 ^ x11 ;
  assign n3282 = n2412 & ~n3005 ;
  assign n3283 = ~n1620 & n2400 ;
  assign n3284 = n3282 | n3283 ;
  assign n3285 = n3284 ^ n40 ^ x11 ;
  assign n3286 = n2461 & ~n2893 ;
  assign n3287 = n2461 & ~n2875 ;
  assign n3288 = n2412 & ~n2987 ;
  assign n3289 = ( n2412 & n3275 ) | ( n2412 & ~n3288 ) | ( n3275 & ~n3288 ) ;
  assign n3290 = n1654 & n2220 ;
  assign n3291 = n3289 ^ n40 ^ x11 ;
  assign n3292 = n2220 & n2466 ;
  assign n3293 = n2216 & n2460 ;
  assign n3294 = ( ~n2221 & n2466 ) | ( ~n2221 & n3293 ) | ( n2466 & n3293 ) ;
  assign n3295 = n3293 | n3294 ;
  assign n3296 = ~n2222 & n2455 ;
  assign n3297 = ( n2455 & n3295 ) | ( n2455 & ~n3296 ) | ( n3295 & ~n3296 ) ;
  assign n3298 = n2221 & n2455 ;
  assign n3299 = ( n2455 & n3292 ) | ( n2455 & ~n3298 ) | ( n3292 & ~n3298 ) ;
  assign n3300 = ( n2222 & n2460 ) | ( n2222 & n3292 ) | ( n2460 & n3292 ) ;
  assign n3301 = ( ~n3287 & n3299 ) | ( ~n3287 & n3300 ) | ( n3299 & n3300 ) ;
  assign n3302 = ( n2461 & ~n3286 ) | ( n2461 & n3297 ) | ( ~n3286 & n3297 ) ;
  assign n3303 = n3287 | n3301 ;
  assign n3304 = n3302 ^ n82 ^ x14 ;
  assign n3305 = n3303 ^ n82 ^ x14 ;
  assign n3306 = ( n3228 & ~n3234 ) | ( n3228 & n3305 ) | ( ~n3234 & n3305 ) ;
  assign n3307 = ( n3236 & ~n3290 ) | ( n3236 & n3304 ) | ( ~n3290 & n3304 ) ;
  assign n3308 = n3305 ^ n3234 ^ n3228 ;
  assign n3309 = n3308 ^ n3291 ^ n3263 ;
  assign n3310 = n3309 ^ n3267 ^ n3261 ;
  assign n3311 = ( n3261 & n3267 ) | ( n3261 & n3309 ) | ( n3267 & n3309 ) ;
  assign n3312 = n3310 ^ n3270 ^ n1540 ;
  assign n3313 = ( n1540 & n3270 ) | ( n1540 & n3310 ) | ( n3270 & n3310 ) ;
  assign n3314 = ( n3263 & ~n3291 ) | ( n3263 & n3308 ) | ( ~n3291 & n3308 ) ;
  assign n3315 = n3304 ^ n3290 ^ n3236 ;
  assign n3316 = ( n3281 & n3306 ) | ( n3281 & ~n3315 ) | ( n3306 & ~n3315 ) ;
  assign n3317 = n3315 ^ n3306 ^ n3281 ;
  assign n3318 = ( ~n3311 & n3314 ) | ( ~n3311 & n3317 ) | ( n3314 & n3317 ) ;
  assign n3319 = n3317 ^ n3314 ^ n3311 ;
  assign n3320 = ( n1628 & n3313 ) | ( n1628 & n3319 ) | ( n3313 & n3319 ) ;
  assign n3321 = n3319 ^ n3313 ^ n1628 ;
  assign n3322 = n1654 & ~n2221 ;
  assign n3323 = ~n1620 & n2455 ;
  assign n3324 = ~n2224 & n2460 ;
  assign n3325 = n2461 & n2997 ;
  assign n3326 = n3323 | n3325 ;
  assign n3327 = ( ~n2224 & n2466 ) | ( ~n2224 & n3325 ) | ( n2466 & n3325 ) ;
  assign n3328 = ~n1620 & n2460 ;
  assign n3329 = n3326 | n3327 ;
  assign n3330 = n2461 & ~n2963 ;
  assign n3331 = n2216 & n2455 ;
  assign n3332 = n3329 ^ n82 ^ x14 ;
  assign n3333 = ~n2224 & n2455 ;
  assign n3334 = n3328 | n3333 ;
  assign n3335 = ( n2216 & n2466 ) | ( n2216 & n3328 ) | ( n2466 & n3328 ) ;
  assign n3336 = n2461 & ~n2987 ;
  assign n3337 = n3334 | n3335 ;
  assign n3338 = n3324 | n3331 ;
  assign n3339 = ( n2461 & ~n3336 ) | ( n2461 & n3337 ) | ( ~n3336 & n3337 ) ;
  assign n3340 = n3322 ^ n3307 ^ n3290 ;
  assign n3341 = ( n2222 & n2466 ) | ( n2222 & n3331 ) | ( n2466 & n3331 ) ;
  assign n3342 = ( ~n3330 & n3338 ) | ( ~n3330 & n3341 ) | ( n3338 & n3341 ) ;
  assign n3343 = n3330 | n3342 ;
  assign n3344 = n3343 ^ n82 ^ x14 ;
  assign n3345 = n3344 ^ n3340 ^ n3285 ;
  assign n3346 = ( n3290 & n3307 ) | ( n3290 & ~n3322 ) | ( n3307 & ~n3322 ) ;
  assign n3347 = n1654 & n2222 ;
  assign n3348 = n3347 ^ n3322 ^ n1776 ;
  assign n3349 = n3339 ^ n82 ^ x14 ;
  assign n3350 = n3345 ^ n3318 ^ n3316 ;
  assign n3351 = ( n3285 & ~n3340 ) | ( n3285 & n3344 ) | ( ~n3340 & n3344 ) ;
  assign n3352 = ( ~n1776 & n3322 ) | ( ~n1776 & n3347 ) | ( n3322 & n3347 ) ;
  assign n3353 = ( n3346 & ~n3348 ) | ( n3346 & n3349 ) | ( ~n3348 & n3349 ) ;
  assign n3354 = ( ~n3316 & n3318 ) | ( ~n3316 & n3345 ) | ( n3318 & n3345 ) ;
  assign n3355 = n2461 & ~n3005 ;
  assign n3356 = n3349 ^ n3348 ^ n3346 ;
  assign n3357 = n3356 ^ n3354 ^ n3351 ;
  assign n3358 = n1654 & n2962 ;
  assign n3359 = n1654 & n2216 ;
  assign n3360 = n3359 ^ n3352 ^ n3332 ;
  assign n3361 = ( n3332 & n3352 ) | ( n3332 & ~n3359 ) | ( n3352 & ~n3359 ) ;
  assign n3362 = ( n1552 & n3320 ) | ( n1552 & n3350 ) | ( n3320 & n3350 ) ;
  assign n3363 = n3350 ^ n3320 ^ n1552 ;
  assign n3364 = ( n1297 & n3357 ) | ( n1297 & n3362 ) | ( n3357 & n3362 ) ;
  assign n3365 = ( ~n3351 & n3354 ) | ( ~n3351 & n3356 ) | ( n3354 & n3356 ) ;
  assign n3366 = n3365 ^ n3360 ^ n3353 ;
  assign n3367 = ( n1630 & n3364 ) | ( n1630 & n3366 ) | ( n3364 & n3366 ) ;
  assign n3368 = ( ~n3353 & n3360 ) | ( ~n3353 & n3365 ) | ( n3360 & n3365 ) ;
  assign n3369 = n3366 ^ n3364 ^ n1630 ;
  assign n3370 = n3362 ^ n3357 ^ n1297 ;
  assign n3371 = ~n1620 & n2466 ;
  assign n3372 = n3355 | n3371 ;
  assign n3373 = n3372 ^ n3358 ^ 1'b0 ;
  assign n3374 = n3373 ^ n3368 ^ n3361 ;
  assign n3375 = ( ~n3361 & n3368 ) | ( ~n3361 & n3373 ) | ( n3368 & n3373 ) ;
  assign n3376 = ( n2216 & ~n2224 ) | ( n2216 & n3372 ) | ( ~n2224 & n3372 ) ;
  assign n3377 = x23 ^ x22 ^ 1'b0 ;
  assign n3378 = n3372 ^ n1654 ^ 1'b0 ;
  assign n3379 = n3374 ^ n3367 ^ n1631 ;
  assign n3380 = ( ~n2216 & n3376 ) | ( ~n2216 & n3378 ) | ( n3376 & n3378 ) ;
  assign n3381 = ( ~n2906 & n2977 ) | ( ~n2906 & n2996 ) | ( n2977 & n2996 ) ;
  assign n3382 = ( n1631 & n3367 ) | ( n1631 & n3374 ) | ( n3367 & n3374 ) ;
  assign n3383 = n2977 ^ n2906 ^ 1'b0 ;
  assign n3384 = n2906 & n3381 ;
  assign n3385 = n3381 ^ n2906 ^ 1'b0 ;
  assign n3386 = ( n2906 & n2977 ) | ( n2906 & n3377 ) | ( n2977 & n3377 ) ;
  assign n3387 = n3385 ^ n3384 ^ n3008 ;
  assign n3388 = n3385 | n3387 ;
  assign n3389 = n3377 & n3385 ;
  assign n3390 = n3389 ^ n3384 ^ n3008 ;
  assign n3391 = n3386 ^ n2996 ^ 1'b0 ;
  assign n3392 = n3008 & n3384 ;
  assign n3393 = n3377 & n3388 ;
  assign n3394 = n2216 ^ n1620 ^ 1'b0 ;
  assign n3395 = n3056 & n3392 ;
  assign n3396 = n3114 & n3395 ;
  assign n3397 = n3393 ^ n3392 ^ n3056 ;
  assign n3398 = n3392 ^ n3388 ^ n3056 ;
  assign n3399 = n1654 & n3394 ;
  assign n3400 = n3399 ^ n3380 ^ n3375 ;
  assign n3401 = n3388 | n3398 ;
  assign n3402 = n3400 ^ n3382 ^ n1446 ;
  assign n3403 = n3377 & n3401 ;
  assign n3404 = ( n1446 & n3382 ) | ( n1446 & n3400 ) | ( n3382 & n3400 ) ;
  assign n3405 = n1632 & n3404 ;
  assign n3406 = n3401 ^ n3395 ^ n3114 ;
  assign n3407 = n744 | n3405 ;
  assign n3408 = n3401 | n3406 ;
  assign n3409 = n3403 ^ n3395 ^ n3114 ;
  assign n3410 = n744 & n3405 ;
  assign n3411 = n3404 ^ n1632 ^ 1'b0 ;
  assign n3412 = n3408 ^ n3396 ^ n3153 ;
  assign n3413 = n3408 | n3412 ;
  assign n3414 = n3377 & n3408 ;
  assign n3415 = n3414 ^ n3396 ^ n3153 ;
  assign n3416 = n3153 & n3396 ;
  assign n3417 = n3416 ^ n3413 ^ n3189 ;
  assign n3418 = n3413 | n3417 ;
  assign n3419 = n3377 & n3413 ;
  assign n3420 = n3419 ^ n3416 ^ n3189 ;
  assign n3421 = n3189 & n3416 ;
  assign n3422 = n3421 ^ n3418 ^ n3212 ;
  assign n3423 = n3418 | n3422 ;
  assign n3424 = n3377 & n3418 ;
  assign n3425 = n3424 ^ n3421 ^ n3212 ;
  assign n3426 = n3212 & n3421 ;
  assign n3427 = n3426 ^ n3423 ^ n3264 ;
  assign n3428 = n3423 | n3427 ;
  assign n3429 = n3377 & n3423 ;
  assign n3430 = n3429 ^ n3426 ^ n3264 ;
  assign n3431 = n3264 & n3426 ;
  assign n3432 = n3431 ^ n3428 ^ n3269 ;
  assign n3433 = n3428 | n3432 ;
  assign n3434 = n3377 & n3428 ;
  assign n3435 = n3434 ^ n3431 ^ n3269 ;
  assign n3436 = n3269 & n3431 ;
  assign n3437 = n3436 ^ n3433 ^ n3312 ;
  assign n3438 = n3433 | n3437 ;
  assign n3439 = n3377 & n3433 ;
  assign n3440 = n3439 ^ n3436 ^ n3312 ;
  assign n3441 = n3312 & n3436 ;
  assign n3442 = n3441 ^ n3438 ^ n3321 ;
  assign n3443 = n3438 | n3442 ;
  assign n3444 = n3377 & n3438 ;
  assign n3445 = n3444 ^ n3441 ^ n3321 ;
  assign n3446 = n3321 & n3441 ;
  assign n3447 = n3446 ^ n3443 ^ n3363 ;
  assign n3448 = n3443 | n3447 ;
  assign n3449 = n3377 & n3443 ;
  assign n3450 = n3449 ^ n3446 ^ n3363 ;
  assign n3451 = n3363 & n3446 ;
  assign n3452 = n3451 ^ n3448 ^ n3370 ;
  assign n3453 = n3448 | n3452 ;
  assign n3454 = n3377 & n3448 ;
  assign n3455 = n3454 ^ n3451 ^ n3370 ;
  assign n3456 = n3370 & n3451 ;
  assign n3457 = n3456 ^ n3453 ^ n3369 ;
  assign n3458 = n3453 | n3457 ;
  assign n3459 = n3377 & n3453 ;
  assign n3460 = n3459 ^ n3456 ^ n3369 ;
  assign n3461 = n3369 & n3456 ;
  assign n3462 = n3461 ^ n3458 ^ n3379 ;
  assign n3463 = n3458 | n3462 ;
  assign n3464 = n3377 & n3458 ;
  assign n3465 = n3464 ^ n3461 ^ n3379 ;
  assign n3466 = n3379 & n3461 ;
  assign n3467 = n3466 ^ n3463 ^ n3402 ;
  assign n3468 = n3463 | n3467 ;
  assign n3469 = n3377 & n3463 ;
  assign n3470 = n3469 ^ n3466 ^ n3402 ;
  assign n3471 = n3402 & n3466 ;
  assign n3472 = n3471 ^ n3468 ^ n3411 ;
  assign n3473 = n3468 | n3472 ;
  assign n3474 = n3377 & n3468 ;
  assign n3475 = n3474 ^ n3471 ^ n3411 ;
  assign n3476 = n3411 & n3471 ;
  assign n3477 = n3410 ^ n1526 ^ 1'b0 ;
  assign n3478 = n1526 & n3410 ;
  assign n3479 = n3476 ^ n3410 ^ n3407 ;
  assign n3480 = n3407 & n3476 ;
  assign n3481 = n3377 & n3473 ;
  assign n3482 = n3481 ^ n3479 ^ 1'b0 ;
  assign n3483 = n3473 | n3479 ;
  assign n3484 = n1634 & n3478 ;
  assign n3485 = n1634 | n3478 ;
  assign n3486 = n3483 ^ n3480 ^ n3477 ;
  assign n3487 = n3377 & n3483 ;
  assign n3488 = ( n3377 & n3486 ) | ( n3377 & n3487 ) | ( n3486 & n3487 ) ;
  assign n3489 = n3487 ^ n3480 ^ n3477 ;
  assign n3490 = n3477 & n3480 ;
  assign n3491 = n3490 ^ n3485 ^ n3484 ;
  assign n3492 = n3485 & n3490 ;
  assign n3493 = ( n2218 & n3484 ) | ( n2218 & n3492 ) | ( n3484 & n3492 ) ;
  assign n3494 = n3492 ^ n3484 ^ n2218 ;
  assign n3495 = ( n3377 & n3488 ) | ( n3377 & n3491 ) | ( n3488 & n3491 ) ;
  assign n3496 = ( n3377 & n3494 ) | ( n3377 & n3495 ) | ( n3494 & n3495 ) ;
  assign n3497 = n3495 ^ n3494 ^ 1'b0 ;
  assign n3498 = n2215 & n3493 ;
  assign n3499 = n3493 ^ n2215 ^ 1'b0 ;
  assign n3500 = n2317 & ~n3498 ;
  assign n3501 = n3491 ^ n3488 ^ 1'b0 ;
  assign n3502 = ( n3377 & n3496 ) | ( n3377 & n3499 ) | ( n3496 & n3499 ) ;
  assign n3503 = n3502 ^ n3498 ^ 1'b0 ;
  assign n3504 = n2317 & ~n3503 ;
  assign n3505 = ( n3377 & ~n3500 ) | ( n3377 & n3502 ) | ( ~n3500 & n3502 ) ;
  assign n3506 = n3499 ^ n3496 ^ 1'b0 ;
  assign y0 = n3383 ;
  assign y1 = n3391 ;
  assign y2 = n3390 ;
  assign y3 = n3397 ;
  assign y4 = n3409 ;
  assign y5 = n3415 ;
  assign y6 = n3420 ;
  assign y7 = n3425 ;
  assign y8 = n3430 ;
  assign y9 = n3435 ;
  assign y10 = n3440 ;
  assign y11 = n3445 ;
  assign y12 = n3450 ;
  assign y13 = n3455 ;
  assign y14 = n3460 ;
  assign y15 = n3465 ;
  assign y16 = n3470 ;
  assign y17 = n3475 ;
  assign y18 = n3482 ;
  assign y19 = n3489 ;
  assign y20 = n3501 ;
  assign y21 = n3497 ;
  assign y22 = n3506 ;
  assign y23 = ~n3504 ;
  assign y24 = n3505 ;
endmodule
