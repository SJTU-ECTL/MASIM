module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 ;
  assign n11 = x3 | x8 ;
  assign n12 = ~x3 & x9 ;
  assign n13 = x1 & n12 ;
  assign n14 = ~x5 & x6 ;
  assign n15 = ~x8 & n14 ;
  assign n16 = ~x8 & x9 ;
  assign n17 = x1 | x3 ;
  assign n18 = n15 & ~n17 ;
  assign n19 = x5 & x8 ;
  assign n20 = ~x6 & x8 ;
  assign n21 = x2 | x8 ;
  assign n22 = x3 | x5 ;
  assign n23 = ~x5 & x8 ;
  assign n24 = x0 | n21 ;
  assign n25 = ~x1 & n16 ;
  assign n26 = x2 & ~n25 ;
  assign n27 = ~x2 & x8 ;
  assign n28 = x2 | x3 ;
  assign n29 = x5 & ~n21 ;
  assign n30 = ( x2 & n21 ) | ( x2 & n28 ) | ( n21 & n28 ) ;
  assign n31 = x6 & ~x8 ;
  assign n32 = x2 & ~n20 ;
  assign n33 = ( ~x1 & x6 ) | ( ~x1 & n31 ) | ( x6 & n31 ) ;
  assign n34 = ( ~x2 & x9 ) | ( ~x2 & n33 ) | ( x9 & n33 ) ;
  assign n35 = ( n25 & ~n26 ) | ( n25 & n34 ) | ( ~n26 & n34 ) ;
  assign n36 = x5 & n32 ;
  assign n37 = n11 & ~n23 ;
  assign n38 = ( x2 & x9 ) | ( x2 & n37 ) | ( x9 & n37 ) ;
  assign n39 = ~x0 & n37 ;
  assign n40 = x0 & n27 ;
  assign n41 = ( n29 & n37 ) | ( n29 & ~n39 ) | ( n37 & ~n39 ) ;
  assign n42 = ( x5 & n30 ) | ( x5 & n36 ) | ( n30 & n36 ) ;
  assign n43 = ( ~x1 & n36 ) | ( ~x1 & n42 ) | ( n36 & n42 ) ;
  assign n44 = ( x3 & n35 ) | ( x3 & n43 ) | ( n35 & n43 ) ;
  assign n45 = n40 ^ x5 ^ x0 ;
  assign n46 = n40 | n45 ;
  assign n47 = n13 & n31 ;
  assign n48 = ( ~n43 & n44 ) | ( ~n43 & n47 ) | ( n44 & n47 ) ;
  assign n49 = ( ~x3 & n16 ) | ( ~x3 & n17 ) | ( n16 & n17 ) ;
  assign n50 = n43 | n48 ;
  assign n51 = ( ~x6 & n12 ) | ( ~x6 & n49 ) | ( n12 & n49 ) ;
  assign n52 = x3 & ~n27 ;
  assign n53 = n52 ^ n23 ^ n22 ;
  assign n54 = x1 & n53 ;
  assign n55 = n18 | n54 ;
  assign n56 = ~n12 & n51 ;
  assign n57 = ~x0 & n30 ;
  assign n58 = ( x1 & n46 ) | ( x1 & n57 ) | ( n46 & n57 ) ;
  assign n59 = ( ~x1 & n41 ) | ( ~x1 & n57 ) | ( n41 & n57 ) ;
  assign n60 = x9 & n55 ;
  assign n61 = ( n55 & n56 ) | ( n55 & ~n60 ) | ( n56 & ~n60 ) ;
  assign n62 = n50 | n61 ;
  assign n63 = x3 & ~x8 ;
  assign n64 = x6 | n63 ;
  assign n65 = ( x3 & n16 ) | ( x3 & n22 ) | ( n16 & n22 ) ;
  assign n66 = ~x2 & n65 ;
  assign n67 = ( x5 & ~n22 ) | ( x5 & n64 ) | ( ~n22 & n64 ) ;
  assign n68 = n58 | n59 ;
  assign n69 = ( x2 & ~x9 ) | ( x2 & n19 ) | ( ~x9 & n19 ) ;
  assign n70 = ~n38 & n69 ;
  assign n71 = x3 | x6 ;
  assign n72 = ( n66 & ~n67 ) | ( n66 & n70 ) | ( ~n67 & n70 ) ;
  assign n73 = ( n15 & ~n67 ) | ( n15 & n71 ) | ( ~n67 & n71 ) ;
  assign n74 = n67 & ~n72 ;
  assign n75 = ( x1 & n72 ) | ( x1 & n74 ) | ( n72 & n74 ) ;
  assign n76 = x1 | x6 ;
  assign n77 = n29 & ~n76 ;
  assign n78 = ~x9 & n77 ;
  assign n79 = ~x3 & n14 ;
  assign n80 = ( ~x9 & n78 ) | ( ~x9 & n79 ) | ( n78 & n79 ) ;
  assign n81 = n75 | n80 ;
  assign n82 = x0 & n81 ;
  assign n83 = x1 & x2 ;
  assign n84 = x1 | x8 ;
  assign n85 = x1 & x5 ;
  assign n86 = ~x2 & x5 ;
  assign n87 = ( x2 & ~x6 ) | ( x2 & n83 ) | ( ~x6 & n83 ) ;
  assign n88 = ( x3 & ~n84 ) | ( x3 & n87 ) | ( ~n84 & n87 ) ;
  assign n89 = x0 & ~x5 ;
  assign n90 = x3 & ~n88 ;
  assign n91 = x6 & n68 ;
  assign n92 = ~x0 & x8 ;
  assign n93 = x2 | n92 ;
  assign n94 = x5 | n92 ;
  assign n95 = x0 & x1 ;
  assign n96 = n76 & ~n95 ;
  assign n97 = ~n93 & n96 ;
  assign n98 = n90 | n97 ;
  assign n99 = ~x5 & n98 ;
  assign n100 = ~x1 & x3 ;
  assign n101 = ( n68 & ~n91 ) | ( n68 & n99 ) | ( ~n91 & n99 ) ;
  assign n102 = x3 & x5 ;
  assign n103 = x0 | x3 ;
  assign n104 = ~x0 & x5 ;
  assign n105 = ~x2 & n103 ;
  assign n106 = n100 & ~n104 ;
  assign n107 = ~n27 & n106 ;
  assign n108 = n16 & n104 ;
  assign n109 = ( x8 & n17 ) | ( x8 & ~n89 ) | ( n17 & ~n89 ) ;
  assign n110 = x8 & ~n109 ;
  assign n111 = n102 ^ n85 ^ x3 ;
  assign n112 = ( ~n22 & n30 ) | ( ~n22 & n86 ) | ( n30 & n86 ) ;
  assign n113 = x1 & n112 ;
  assign n114 = ( x8 & n110 ) | ( x8 & ~n111 ) | ( n110 & ~n111 ) ;
  assign n115 = ( n105 & n110 ) | ( n105 & n114 ) | ( n110 & n114 ) ;
  assign n116 = x1 | x2 ;
  assign n117 = x1 | x9 ;
  assign n118 = ( n106 & ~n107 ) | ( n106 & n113 ) | ( ~n107 & n113 ) ;
  assign n119 = n83 & ~n102 ;
  assign n120 = ~n94 & n119 ;
  assign n121 = ( n115 & n119 ) | ( n115 & ~n120 ) | ( n119 & ~n120 ) ;
  assign n122 = ~x2 & n117 ;
  assign n123 = ( ~n12 & n111 ) | ( ~n12 & n122 ) | ( n111 & n122 ) ;
  assign n124 = x9 ^ x1 ^ 1'b0 ;
  assign n125 = x1 | x5 ;
  assign n126 = ~n111 & n123 ;
  assign n127 = x0 & n85 ;
  assign n128 = ( x0 & n63 ) | ( x0 & n127 ) | ( n63 & n127 ) ;
  assign n129 = ( ~n116 & n127 ) | ( ~n116 & n128 ) | ( n127 & n128 ) ;
  assign n130 = n124 & n125 ;
  assign n131 = x2 & ~x3 ;
  assign n132 = ~n126 & n130 ;
  assign n133 = ( n126 & n131 ) | ( n126 & ~n132 ) | ( n131 & ~n132 ) ;
  assign n134 = n118 ^ x9 ^ 1'b0 ;
  assign n135 = ( n118 & n121 ) | ( n118 & ~n134 ) | ( n121 & ~n134 ) ;
  assign n136 = ~x0 & n13 ;
  assign n137 = x2 & n125 ;
  assign n138 = ( x3 & x5 ) | ( x3 & n137 ) | ( x5 & n137 ) ;
  assign n139 = n129 | n138 ;
  assign n140 = x5 & ~x9 ;
  assign n141 = ( n13 & ~n116 ) | ( n13 & n140 ) | ( ~n116 & n140 ) ;
  assign n142 = ( ~x0 & n136 ) | ( ~x0 & n141 ) | ( n136 & n141 ) ;
  assign n143 = x5 & ~x8 ;
  assign n144 = n133 | n142 ;
  assign n145 = x6 | x8 ;
  assign n146 = n144 & ~n145 ;
  assign n147 = ( ~x6 & n135 ) | ( ~x6 & n146 ) | ( n135 & n146 ) ;
  assign n148 = x3 & n83 ;
  assign n149 = ~n143 & n148 ;
  assign n150 = x6 & n139 ;
  assign n151 = ( n148 & ~n149 ) | ( n148 & n150 ) | ( ~n149 & n150 ) ;
  assign n152 = x2 & ~x9 ;
  assign n153 = ( ~x0 & n102 ) | ( ~x0 & n152 ) | ( n102 & n152 ) ;
  assign n154 = n20 & n152 ;
  assign n155 = ( x0 & n92 ) | ( x0 & n94 ) | ( n92 & n94 ) ;
  assign n156 = n151 ^ x9 ^ 1'b0 ;
  assign n157 = ( n101 & n151 ) | ( n101 & ~n156 ) | ( n151 & ~n156 ) ;
  assign n158 = x3 & n86 ;
  assign n159 = x0 & ~n158 ;
  assign n160 = ( n153 & n158 ) | ( n153 & ~n159 ) | ( n158 & ~n159 ) ;
  assign n161 = x3 & ~x6 ;
  assign n162 = x6 & x8 ;
  assign n163 = n92 & ~n161 ;
  assign n164 = ~x3 & x8 ;
  assign n165 = n162 ^ x9 ^ 1'b0 ;
  assign n166 = ( n31 & n92 ) | ( n31 & ~n163 ) | ( n92 & ~n163 ) ;
  assign n167 = ( n162 & n165 ) | ( n162 & n166 ) | ( n165 & n166 ) ;
  assign n168 = x8 & x9 ;
  assign n169 = ( x0 & n164 ) | ( x0 & n168 ) | ( n164 & n168 ) ;
  assign n170 = x6 & x9 ;
  assign n171 = n168 ^ x3 ^ 1'b0 ;
  assign n172 = ( x0 & ~n164 ) | ( x0 & n170 ) | ( ~n164 & n170 ) ;
  assign n173 = ( ~x6 & n169 ) | ( ~x6 & n171 ) | ( n169 & n171 ) ;
  assign n174 = x8 | x9 ;
  assign n175 = n71 | n174 ;
  assign n176 = ~n170 & n172 ;
  assign n177 = x5 | x9 ;
  assign n178 = ( x2 & n173 ) | ( x2 & ~n175 ) | ( n173 & ~n175 ) ;
  assign n179 = n145 & ~n177 ;
  assign n180 = x5 | n168 ;
  assign n181 = ( x2 & n145 ) | ( x2 & ~n179 ) | ( n145 & ~n179 ) ;
  assign n182 = ( x0 & n167 ) | ( x0 & ~n176 ) | ( n167 & ~n176 ) ;
  assign n183 = x1 & x9 ;
  assign n184 = ( n19 & n181 ) | ( n19 & n183 ) | ( n181 & n183 ) ;
  assign n185 = ( x2 & n175 ) | ( x2 & ~n182 ) | ( n175 & ~n182 ) ;
  assign n186 = x5 & x9 ;
  assign n187 = ~n178 & n185 ;
  assign n188 = ~x6 & n181 ;
  assign n189 = ( n184 & n186 ) | ( n184 & ~n188 ) | ( n186 & ~n188 ) ;
  assign n190 = n184 & ~n189 ;
  assign n191 = ~x6 & n11 ;
  assign n192 = x8 & n186 ;
  assign n193 = ( x3 & ~n181 ) | ( x3 & n190 ) | ( ~n181 & n190 ) ;
  assign n194 = x8 & ~x9 ;
  assign n195 = n145 & ~n194 ;
  assign n196 = ( x1 & n162 ) | ( x1 & n194 ) | ( n162 & n194 ) ;
  assign n197 = ~x2 & n196 ;
  assign n198 = ( x2 & n11 ) | ( x2 & ~n197 ) | ( n11 & ~n197 ) ;
  assign n199 = ( n124 & ~n197 ) | ( n124 & n198 ) | ( ~n197 & n198 ) ;
  assign n200 = n84 & n124 ;
  assign n201 = x6 | n192 ;
  assign n202 = x2 & n161 ;
  assign n203 = ( ~x3 & n170 ) | ( ~x3 & n177 ) | ( n170 & n177 ) ;
  assign n204 = ( ~x3 & n92 ) | ( ~x3 & n203 ) | ( n92 & n203 ) ;
  assign n205 = ~n180 & n202 ;
  assign n206 = ~x3 & n201 ;
  assign n207 = x8 | n177 ;
  assign n208 = ~x2 & n204 ;
  assign n209 = ( n205 & n206 ) | ( n205 & ~n208 ) | ( n206 & ~n208 ) ;
  assign n210 = n208 | n209 ;
  assign n211 = ~x1 & x9 ;
  assign n212 = n207 ^ n201 ^ x6 ;
  assign n213 = x2 & ~n212 ;
  assign n214 = ( n92 & n170 ) | ( n92 & n201 ) | ( n170 & n201 ) ;
  assign n215 = ~x9 & n14 ;
  assign n216 = n73 | n213 ;
  assign n217 = x1 & n216 ;
  assign n218 = ( ~n84 & n161 ) | ( ~n84 & n215 ) | ( n161 & n215 ) ;
  assign n219 = ( x7 & n89 ) | ( x7 & n202 ) | ( n89 & n202 ) ;
  assign n220 = x2 & n14 ;
  assign n221 = n217 | n220 ;
  assign n222 = x9 & n28 ;
  assign n223 = ( n14 & n202 ) | ( n14 & n222 ) | ( n202 & n222 ) ;
  assign n224 = x6 & ~n211 ;
  assign n225 = ( ~x1 & n218 ) | ( ~x1 & n223 ) | ( n218 & n223 ) ;
  assign n226 = ( n31 & n200 ) | ( n31 & n224 ) | ( n200 & n224 ) ;
  assign n227 = ( n32 & n76 ) | ( n32 & n226 ) | ( n76 & n226 ) ;
  assign n228 = ( n23 & n192 ) | ( n23 & n226 ) | ( n192 & n226 ) ;
  assign n229 = ( n193 & ~n225 ) | ( n193 & n228 ) | ( ~n225 & n228 ) ;
  assign n230 = n225 | n229 ;
  assign n231 = x2 & x3 ;
  assign n232 = x0 | n227 ;
  assign n233 = n192 & n231 ;
  assign n234 = ( x3 & n161 ) | ( x3 & n231 ) | ( n161 & n231 ) ;
  assign n235 = ~x1 & n174 ;
  assign n236 = n117 | n234 ;
  assign n237 = n82 | n230 ;
  assign n238 = x7 & ~n235 ;
  assign n239 = ( n219 & ~n235 ) | ( n219 & n238 ) | ( ~n235 & n238 ) ;
  assign n240 = x2 & ~n235 ;
  assign n241 = ( x0 & n224 ) | ( x0 & n240 ) | ( n224 & n240 ) ;
  assign n242 = ( n227 & n232 ) | ( n227 & n241 ) | ( n232 & n241 ) ;
  assign n243 = ( x3 & x5 ) | ( x3 & ~n242 ) | ( x5 & ~n242 ) ;
  assign n244 = ~n147 & n243 ;
  assign n245 = ( x3 & n147 ) | ( x3 & ~n244 ) | ( n147 & ~n244 ) ;
  assign n246 = x0 & x3 ;
  assign n247 = x9 ^ x8 ^ 1'b0 ;
  assign n248 = ( x2 & x3 ) | ( x2 & ~n247 ) | ( x3 & ~n247 ) ;
  assign n249 = x5 & n248 ;
  assign n250 = x2 & x9 ;
  assign n251 = ( x0 & x8 ) | ( x0 & n140 ) | ( x8 & n140 ) ;
  assign n252 = n143 & n250 ;
  assign n253 = n251 | n252 ;
  assign n254 = x9 ^ x2 ^ 1'b0 ;
  assign n255 = ( ~x0 & x8 ) | ( ~x0 & n254 ) | ( x8 & n254 ) ;
  assign n256 = ( n252 & n253 ) | ( n252 & n255 ) | ( n253 & n255 ) ;
  assign n257 = ~x3 & n256 ;
  assign n258 = x8 & ~n257 ;
  assign n259 = ( n160 & n257 ) | ( n160 & ~n258 ) | ( n257 & ~n258 ) ;
  assign n260 = x2 & ~n174 ;
  assign n261 = x0 & ~x2 ;
  assign n262 = ( x2 & n249 ) | ( x2 & n261 ) | ( n249 & n261 ) ;
  assign n263 = ~n246 & n260 ;
  assign n264 = ( n260 & n262 ) | ( n260 & ~n263 ) | ( n262 & ~n263 ) ;
  assign n265 = ( x2 & x3 ) | ( x2 & x6 ) | ( x3 & x6 ) ;
  assign n266 = x6 & ~n247 ;
  assign n267 = ( n31 & n207 ) | ( n31 & ~n266 ) | ( n207 & ~n266 ) ;
  assign n268 = ~x2 & x3 ;
  assign n269 = ( ~x1 & n233 ) | ( ~x1 & n264 ) | ( n233 & n264 ) ;
  assign n270 = ~n254 & n266 ;
  assign n271 = ~n140 & n268 ;
  assign n272 = ( n259 & n268 ) | ( n259 & ~n271 ) | ( n268 & ~n271 ) ;
  assign n273 = ( x3 & n246 ) | ( x3 & ~n266 ) | ( n246 & ~n266 ) ;
  assign n274 = x0 | x9 ;
  assign n275 = ( x1 & n233 ) | ( x1 & n272 ) | ( n233 & n272 ) ;
  assign n276 = n269 | n275 ;
  assign n277 = x0 & n162 ;
  assign n278 = ( x9 & n24 ) | ( x9 & ~n277 ) | ( n24 & ~n277 ) ;
  assign n279 = ~n16 & n274 ;
  assign n280 = ( x3 & n265 ) | ( x3 & n279 ) | ( n265 & n279 ) ;
  assign n281 = x2 & n174 ;
  assign n282 = n273 & n280 ;
  assign n283 = n278 & ~n281 ;
  assign n284 = ( n191 & n278 ) | ( n191 & n283 ) | ( n278 & n283 ) ;
  assign n285 = ~x9 & n31 ;
  assign n286 = n268 & n285 ;
  assign n287 = ( ~x3 & n282 ) | ( ~x3 & n284 ) | ( n282 & n284 ) ;
  assign n288 = ( x1 & ~n286 ) | ( x1 & n287 ) | ( ~n286 & n287 ) ;
  assign n289 = x5 | x7 ;
  assign n290 = ~x6 & n276 ;
  assign n291 = ( x1 & ~n187 ) | ( x1 & n286 ) | ( ~n187 & n286 ) ;
  assign n292 = n288 & n291 ;
  assign n293 = ( n288 & n289 ) | ( n288 & ~n292 ) | ( n289 & ~n292 ) ;
  assign n294 = ( x7 & ~n290 ) | ( x7 & n293 ) | ( ~n290 & n293 ) ;
  assign n295 = x1 & ~x8 ;
  assign n296 = ( n131 & n211 ) | ( n131 & n295 ) | ( n211 & n295 ) ;
  assign n297 = ( x8 & n236 ) | ( x8 & ~n250 ) | ( n236 & ~n250 ) ;
  assign n298 = ~x0 & n297 ;
  assign n299 = ( n22 & ~n24 ) | ( n22 & n183 ) | ( ~n24 & n183 ) ;
  assign n300 = ( ~n93 & n162 ) | ( ~n93 & n295 ) | ( n162 & n295 ) ;
  assign n301 = n295 & n298 ;
  assign n302 = ( n296 & n298 ) | ( n296 & n301 ) | ( n298 & n301 ) ;
  assign n303 = x5 & x6 ;
  assign n304 = ( x6 & n131 ) | ( x6 & n303 ) | ( n131 & n303 ) ;
  assign n305 = ( x5 & n297 ) | ( x5 & ~n302 ) | ( n297 & ~n302 ) ;
  assign n306 = ( x5 & x8 ) | ( x5 & x9 ) | ( x8 & x9 ) ;
  assign n307 = ( n279 & n285 ) | ( n279 & ~n306 ) | ( n285 & ~n306 ) ;
  assign n308 = n23 | n170 ;
  assign n309 = ~n162 & n308 ;
  assign n310 = ( n180 & n303 ) | ( n180 & n309 ) | ( n303 & n309 ) ;
  assign n311 = n261 & n309 ;
  assign n312 = ~x3 & n306 ;
  assign n313 = ( ~x2 & n108 ) | ( ~x2 & n311 ) | ( n108 & n311 ) ;
  assign n314 = x0 | x6 ;
  assign n315 = ~x0 & n131 ;
  assign n316 = ~x0 & n308 ;
  assign n317 = ( x2 & ~n267 ) | ( x2 & n316 ) | ( ~n267 & n316 ) ;
  assign n318 = ~x0 & x2 ;
  assign n319 = ( ~n261 & n314 ) | ( ~n261 & n318 ) | ( n314 & n318 ) ;
  assign n320 = n23 & n319 ;
  assign n321 = ( x8 & n31 ) | ( x8 & ~n320 ) | ( n31 & ~n320 ) ;
  assign n322 = ( x1 & n210 ) | ( x1 & n304 ) | ( n210 & n304 ) ;
  assign n323 = n312 ^ x2 ^ 1'b0 ;
  assign n324 = x9 & ~n321 ;
  assign n325 = ( ~n313 & n321 ) | ( ~n313 & n324 ) | ( n321 & n324 ) ;
  assign n326 = x1 & ~n325 ;
  assign n327 = x5 | x6 ;
  assign n328 = n154 | n326 ;
  assign n329 = x4 & n327 ;
  assign n330 = n329 ^ x3 ^ 1'b0 ;
  assign n331 = ( ~n214 & n329 ) | ( ~n214 & n330 ) | ( n329 & n330 ) ;
  assign n332 = ( ~n312 & n323 ) | ( ~n312 & n331 ) | ( n323 & n331 ) ;
  assign n333 = x2 | n17 ;
  assign n334 = x0 & ~n333 ;
  assign n335 = ( x1 & ~n304 ) | ( x1 & n332 ) | ( ~n304 & n332 ) ;
  assign n336 = ( x7 & ~n315 ) | ( x7 & n334 ) | ( ~n315 & n334 ) ;
  assign n337 = ( ~n239 & n335 ) | ( ~n239 & n336 ) | ( n335 & n336 ) ;
  assign n338 = ( ~n322 & n336 ) | ( ~n322 & n337 ) | ( n336 & n337 ) ;
  assign n339 = ~n336 & n338 ;
  assign n340 = x4 & ~n333 ;
  assign n341 = x5 & n183 ;
  assign n342 = ( ~x4 & n339 ) | ( ~x4 & n340 ) | ( n339 & n340 ) ;
  assign n343 = ( x6 & x9 ) | ( x6 & ~n341 ) | ( x9 & ~n341 ) ;
  assign n344 = n137 & ~n341 ;
  assign n345 = ( ~n341 & n343 ) | ( ~n341 & n344 ) | ( n343 & n344 ) ;
  assign n346 = ( x0 & x2 ) | ( x0 & ~x8 ) | ( x2 & ~x8 ) ;
  assign n347 = x4 & x8 ;
  assign n348 = ( ~x6 & n143 ) | ( ~x6 & n347 ) | ( n143 & n347 ) ;
  assign n349 = ( ~x0 & x9 ) | ( ~x0 & n27 ) | ( x9 & n27 ) ;
  assign n350 = n349 ^ n346 ^ 1'b0 ;
  assign n351 = n76 | n350 ;
  assign n352 = ( x6 & ~n299 ) | ( x6 & n351 ) | ( ~n299 & n351 ) ;
  assign n353 = n22 | n352 ;
  assign n354 = ( x7 & n245 ) | ( x7 & ~n353 ) | ( n245 & ~n353 ) ;
  assign n355 = n245 & ~n354 ;
  assign n356 = x4 & x9 ;
  assign n357 = n356 ^ n170 ^ x6 ;
  assign n358 = ( x5 & ~x6 ) | ( x5 & n347 ) | ( ~x6 & n347 ) ;
  assign n359 = ( x4 & n353 ) | ( x4 & ~n355 ) | ( n353 & ~n355 ) ;
  assign n360 = ( x5 & x6 ) | ( x5 & ~n174 ) | ( x6 & ~n174 ) ;
  assign n361 = n358 & n360 ;
  assign n362 = ~x8 & n303 ;
  assign n363 = ( ~x8 & n357 ) | ( ~x8 & n362 ) | ( n357 & n362 ) ;
  assign n364 = ( n361 & ~n362 ) | ( n361 & n363 ) | ( ~n362 & n363 ) ;
  assign n365 = x0 & x9 ;
  assign n366 = x0 | x2 ;
  assign n367 = ( ~x0 & x7 ) | ( ~x0 & n364 ) | ( x7 & n364 ) ;
  assign n368 = ~n333 & n367 ;
  assign n369 = x8 & n365 ;
  assign n370 = ( n348 & n356 ) | ( n348 & ~n366 ) | ( n356 & ~n366 ) ;
  assign n371 = ( n349 & n366 ) | ( n349 & ~n369 ) | ( n366 & ~n369 ) ;
  assign n372 = ~x2 & n317 ;
  assign n373 = x5 & ~n371 ;
  assign n374 = ( n317 & ~n372 ) | ( n317 & n373 ) | ( ~n372 & n373 ) ;
  assign n375 = n281 | n369 ;
  assign n376 = n174 & ~n369 ;
  assign n377 = ( n174 & n235 ) | ( n174 & n376 ) | ( n235 & n376 ) ;
  assign n378 = n222 | n246 ;
  assign n379 = x2 | x5 ;
  assign n380 = ( x2 & ~n100 ) | ( x2 & n379 ) | ( ~n100 & n379 ) ;
  assign n381 = n174 | n380 ;
  assign n382 = ~x1 & x8 ;
  assign n383 = ( ~x1 & x5 ) | ( ~x1 & n376 ) | ( x5 & n376 ) ;
  assign n384 = ( n222 & ~n381 ) | ( n222 & n382 ) | ( ~n381 & n382 ) ;
  assign n385 = n381 & ~n384 ;
  assign n386 = x4 & n374 ;
  assign n387 = ( n84 & n250 ) | ( n84 & n382 ) | ( n250 & n382 ) ;
  assign n388 = ( x1 & x5 ) | ( x1 & n250 ) | ( x5 & n250 ) ;
  assign n389 = ~n383 & n388 ;
  assign n390 = ~x6 & x9 ;
  assign n391 = n370 & ~n390 ;
  assign n392 = ~x4 & n157 ;
  assign n393 = x0 & ~n385 ;
  assign n394 = ~n366 & n391 ;
  assign n395 = ~x4 & n328 ;
  assign n396 = ( n374 & ~n386 ) | ( n374 & n394 ) | ( ~n386 & n394 ) ;
  assign n397 = ~x1 & x2 ;
  assign n398 = ~n17 & n396 ;
  assign n399 = n152 ^ x8 ^ 1'b0 ;
  assign n400 = ( n240 & n397 ) | ( n240 & ~n399 ) | ( n397 & ~n399 ) ;
  assign n401 = n389 | n400 ;
  assign n402 = ~x3 & n401 ;
  assign n403 = x6 | n399 ;
  assign n404 = ( ~x3 & n395 ) | ( ~x3 & n398 ) | ( n395 & n398 ) ;
  assign n405 = ( n387 & n399 ) | ( n387 & n403 ) | ( n399 & n403 ) ;
  assign n406 = ( x3 & ~n199 ) | ( x3 & n405 ) | ( ~n199 & n405 ) ;
  assign n407 = n199 & ~n406 ;
  assign n408 = ( x0 & x5 ) | ( x0 & ~n407 ) | ( x5 & ~n407 ) ;
  assign n409 = ~x5 & n408 ;
  assign n410 = n392 | n404 ;
  assign n411 = n393 | n402 ;
  assign n412 = ~x6 & n411 ;
  assign n413 = n409 | n412 ;
  assign n414 = x9 & n300 ;
  assign n415 = x1 & ~x9 ;
  assign n416 = ( x9 & n95 ) | ( x9 & n414 ) | ( n95 & n414 ) ;
  assign n417 = ( ~x8 & n414 ) | ( ~x8 & n416 ) | ( n414 & n416 ) ;
  assign n418 = n155 & ~n415 ;
  assign n419 = ( n155 & n417 ) | ( n155 & ~n418 ) | ( n417 & ~n418 ) ;
  assign n420 = x7 & x8 ;
  assign n421 = ~x9 & n420 ;
  assign n422 = ( n318 & ~n350 ) | ( n318 & n421 ) | ( ~n350 & n421 ) ;
  assign n423 = x2 & n415 ;
  assign n424 = ( n200 & ~n314 ) | ( n200 & n423 ) | ( ~n314 & n423 ) ;
  assign n425 = ~n22 & n294 ;
  assign n426 = ( ~n274 & n379 ) | ( ~n274 & n423 ) | ( n379 & n423 ) ;
  assign n427 = ( n76 & n422 ) | ( n76 & ~n425 ) | ( n422 & ~n425 ) ;
  assign n428 = n422 & ~n427 ;
  assign n429 = ~x2 & n415 ;
  assign n430 = ( x6 & n250 ) | ( x6 & n429 ) | ( n250 & n429 ) ;
  assign n431 = ( x4 & n294 ) | ( x4 & ~n428 ) | ( n294 & ~n428 ) ;
  assign n432 = x3 ^ x1 ^ 1'b0 ;
  assign n433 = ( ~x3 & n378 ) | ( ~x3 & n432 ) | ( n378 & n432 ) ;
  assign n434 = ~x0 & n429 ;
  assign n435 = n426 | n433 ;
  assign n436 = ( x0 & x8 ) | ( x0 & ~n421 ) | ( x8 & ~n421 ) ;
  assign n437 = ( x8 & n397 ) | ( x8 & ~n421 ) | ( n397 & ~n421 ) ;
  assign n438 = ( n434 & ~n436 ) | ( n434 & n437 ) | ( ~n436 & n437 ) ;
  assign n439 = x2 & x7 ;
  assign n440 = ( x7 & n438 ) | ( x7 & ~n439 ) | ( n438 & ~n439 ) ;
  assign n441 = ( ~n377 & n438 ) | ( ~n377 & n440 ) | ( n438 & n440 ) ;
  assign n442 = ( x0 & x1 ) | ( x0 & ~x8 ) | ( x1 & ~x8 ) ;
  assign n443 = ( x1 & ~x9 ) | ( x1 & n442 ) | ( ~x9 & n442 ) ;
  assign n444 = x0 & ~x9 ;
  assign n445 = ~n84 & n444 ;
  assign n446 = ( n365 & n443 ) | ( n365 & n445 ) | ( n443 & n445 ) ;
  assign n447 = ( n415 & ~n429 ) | ( n415 & n446 ) | ( ~n429 & n446 ) ;
  assign n448 = ~x0 & x9 ;
  assign n449 = n424 | n447 ;
  assign n450 = ~x5 & n449 ;
  assign n451 = n419 | n450 ;
  assign n452 = x8 & n448 ;
  assign n453 = n307 ^ x2 ^ 1'b0 ;
  assign n454 = ( n307 & n452 ) | ( n307 & n453 ) | ( n452 & n453 ) ;
  assign n455 = x4 & ~x7 ;
  assign n456 = x0 | n116 ;
  assign n457 = ( ~n22 & n455 ) | ( ~n22 & n456 ) | ( n455 & n456 ) ;
  assign n458 = ~n456 & n457 ;
  assign n459 = n359 & ~n458 ;
  assign n460 = ( ~x6 & n103 ) | ( ~x6 & n430 ) | ( n103 & n430 ) ;
  assign n461 = n430 & ~n460 ;
  assign n462 = ( ~x5 & x6 ) | ( ~x5 & n379 ) | ( x6 & n379 ) ;
  assign n463 = n448 & n462 ;
  assign n464 = ( n365 & n420 ) | ( n365 & n445 ) | ( n420 & n445 ) ;
  assign n465 = x3 & n451 ;
  assign n466 = n103 | n379 ;
  assign n467 = x9 ^ x0 ^ 1'b0 ;
  assign n468 = n86 & ~n467 ;
  assign n469 = ~n76 & n455 ;
  assign n470 = ( ~x8 & n463 ) | ( ~x8 & n468 ) | ( n463 & n468 ) ;
  assign n471 = x1 | n445 ;
  assign n472 = ( ~n274 & n445 ) | ( ~n274 & n471 ) | ( n445 & n471 ) ;
  assign n473 = ~x6 & n375 ;
  assign n474 = ( n375 & n470 ) | ( n375 & ~n473 ) | ( n470 & ~n473 ) ;
  assign n475 = n27 & n415 ;
  assign n476 = ( n431 & n466 ) | ( n431 & ~n469 ) | ( n466 & ~n469 ) ;
  assign n477 = x1 & ~n467 ;
  assign n478 = ( n464 & n471 ) | ( n464 & n472 ) | ( n471 & n472 ) ;
  assign n479 = n454 ^ x1 ^ 1'b0 ;
  assign n480 = ( n454 & n474 ) | ( n454 & n479 ) | ( n474 & n479 ) ;
  assign n481 = n431 & n476 ;
  assign n482 = n465 | n480 ;
  assign n483 = x5 | n211 ;
  assign n484 = ( x5 & ~n366 ) | ( x5 & n483 ) | ( ~n366 & n483 ) ;
  assign n485 = ~x7 & n435 ;
  assign n486 = ( x2 & x6 ) | ( x2 & n477 ) | ( x6 & n477 ) ;
  assign n487 = n397 & n444 ;
  assign n488 = x5 & n486 ;
  assign n489 = ( x6 & n484 ) | ( x6 & n488 ) | ( n484 & n488 ) ;
  assign n490 = x2 | n444 ;
  assign n491 = ( ~x8 & n95 ) | ( ~x8 & n490 ) | ( n95 & n490 ) ;
  assign n492 = x2 | n211 ;
  assign n493 = n303 & n490 ;
  assign n494 = ( x5 & n477 ) | ( x5 & n493 ) | ( n477 & n493 ) ;
  assign n495 = ( ~n28 & n493 ) | ( ~n28 & n494 ) | ( n493 & n494 ) ;
  assign n496 = n461 | n495 ;
  assign n497 = ( x1 & x7 ) | ( x1 & ~x9 ) | ( x7 & ~x9 ) ;
  assign n498 = ( x1 & n444 ) | ( x1 & ~n497 ) | ( n444 & ~n497 ) ;
  assign n499 = ~n497 & n498 ;
  assign n500 = x1 & ~n448 ;
  assign n501 = ( n22 & n492 ) | ( n22 & ~n500 ) | ( n492 & ~n500 ) ;
  assign n502 = n500 | n501 ;
  assign n503 = ( x2 & ~n499 ) | ( x2 & n502 ) | ( ~n499 & n502 ) ;
  assign n504 = x8 | n503 ;
  assign n505 = ( x8 & ~n485 ) | ( x8 & n504 ) | ( ~n485 & n504 ) ;
  assign n506 = ( ~x5 & x6 ) | ( ~x5 & n441 ) | ( x6 & n441 ) ;
  assign n507 = ~x1 & n177 ;
  assign n508 = x8 & ~n489 ;
  assign n509 = x0 | x1 ;
  assign n510 = ( ~x8 & n448 ) | ( ~x8 & n500 ) | ( n448 & n500 ) ;
  assign n511 = ~x5 & n510 ;
  assign n512 = ~x6 & n506 ;
  assign n513 = ( ~x5 & n487 ) | ( ~x5 & n511 ) | ( n487 & n511 ) ;
  assign n514 = x6 | n505 ;
  assign n515 = n152 & ~n509 ;
  assign n516 = n345 ^ x0 ^ 1'b0 ;
  assign n517 = ( x8 & ~n508 ) | ( x8 & n513 ) | ( ~n508 & n513 ) ;
  assign n518 = x2 & n177 ;
  assign n519 = ( ~n345 & n516 ) | ( ~n345 & n518 ) | ( n516 & n518 ) ;
  assign n520 = x8 | n117 ;
  assign n521 = x5 | n270 ;
  assign n522 = ( n270 & ~n520 ) | ( n270 & n521 ) | ( ~n520 & n521 ) ;
  assign n523 = ( x2 & n270 ) | ( x2 & n448 ) | ( n270 & n448 ) ;
  assign n524 = ( n521 & n522 ) | ( n521 & n523 ) | ( n522 & n523 ) ;
  assign n525 = ( x8 & n270 ) | ( x8 & n519 ) | ( n270 & n519 ) ;
  assign n526 = ~x5 & n420 ;
  assign n527 = n524 | n525 ;
  assign n528 = x7 & n527 ;
  assign n529 = ( n512 & n527 ) | ( n512 & ~n528 ) | ( n527 & ~n528 ) ;
  assign n530 = ( n497 & n507 ) | ( n497 & ~n526 ) | ( n507 & ~n526 ) ;
  assign n531 = x3 & n529 ;
  assign n532 = ~x7 & n482 ;
  assign n533 = ( n529 & ~n531 ) | ( n529 & n532 ) | ( ~n531 & n532 ) ;
  assign n534 = n475 | n491 ;
  assign n535 = n515 & n526 ;
  assign n536 = x4 | x6 ;
  assign n537 = x7 & ~n177 ;
  assign n538 = ( n507 & n530 ) | ( n507 & ~n537 ) | ( n530 & ~n537 ) ;
  assign n539 = x2 & n509 ;
  assign n540 = ( x8 & ~n475 ) | ( x8 & n539 ) | ( ~n475 & n539 ) ;
  assign n541 = ( n475 & n534 ) | ( n475 & ~n540 ) | ( n534 & ~n540 ) ;
  assign n542 = ~x7 & n541 ;
  assign n543 = ( n515 & n541 ) | ( n515 & ~n542 ) | ( n541 & ~n542 ) ;
  assign n544 = x7 & n410 ;
  assign n545 = ( ~n22 & n536 ) | ( ~n22 & n543 ) | ( n536 & n543 ) ;
  assign n546 = ( x0 & x2 ) | ( x0 & ~n538 ) | ( x2 & ~n538 ) ;
  assign n547 = ~n536 & n545 ;
  assign n548 = ( n410 & ~n544 ) | ( n410 & n547 ) | ( ~n544 & n547 ) ;
  assign n549 = ~x2 & n546 ;
  assign n550 = n535 | n549 ;
  assign n551 = ~x3 & n550 ;
  assign n552 = ( x6 & n514 ) | ( x6 & ~n551 ) | ( n514 & ~n551 ) ;
  assign n553 = x0 | n28 ;
  assign n554 = n520 | n553 ;
  assign n555 = x8 & n496 ;
  assign n556 = ( ~n305 & n554 ) | ( ~n305 & n555 ) | ( n554 & n555 ) ;
  assign n557 = n554 & ~n556 ;
  assign n558 = x3 & n557 ;
  assign n559 = n517 & n558 ;
  assign n560 = ( x7 & n557 ) | ( x7 & ~n559 ) | ( n557 & ~n559 ) ;
  assign n561 = ~n552 & n560 ;
  assign n562 = ~x7 & n368 ;
  assign n563 = ( x4 & n560 ) | ( x4 & ~n561 ) | ( n560 & ~n561 ) ;
  assign n564 = ~n562 & n563 ;
  assign n565 = ~x4 & n62 ;
  assign n566 = ( x2 & ~x5 ) | ( x2 & n195 ) | ( ~x5 & n195 ) ;
  assign n567 = x3 & ~x4 ;
  assign n568 = ~x1 & x4 ;
  assign n569 = ( x4 & ~n28 ) | ( x4 & n567 ) | ( ~n28 & n567 ) ;
  assign n570 = ( n567 & n568 ) | ( n567 & n569 ) | ( n568 & n569 ) ;
  assign n571 = ~n566 & n570 ;
  assign n572 = n565 | n571 ;
  assign n573 = ~x0 & n572 ;
  assign n574 = ~x4 & n413 ;
  assign n575 = n573 | n574 ;
  assign n576 = ( ~x4 & n28 ) | ( ~x4 & n478 ) | ( n28 & n478 ) ;
  assign n577 = ~n28 & n576 ;
  assign n578 = ( ~x5 & x6 ) | ( ~x5 & n577 ) | ( x6 & n577 ) ;
  assign n579 = ~x6 & n578 ;
  assign n580 = x7 & n575 ;
  assign n581 = ( n575 & n579 ) | ( n575 & ~n580 ) | ( n579 & ~n580 ) ;
  assign n582 = n310 & n569 ;
  assign n583 = x3 & ~n390 ;
  assign n584 = ( x2 & x4 ) | ( x2 & ~x6 ) | ( x4 & ~x6 ) ;
  assign n585 = x2 & ~n584 ;
  assign n586 = ( ~x4 & n583 ) | ( ~x4 & n585 ) | ( n583 & n585 ) ;
  assign n587 = n582 | n586 ;
  assign n588 = ~x1 & n587 ;
  assign n589 = ~x4 & n221 ;
  assign n590 = n588 | n589 ;
  assign n591 = ~x0 & n590 ;
  assign n592 = ~x4 & n237 ;
  assign n593 = n591 | n592 ;
  assign n594 = ~x7 & n593 ;
  assign n595 = ~x4 & n539 ;
  assign n596 = ( ~n456 & n567 ) | ( ~n456 & n569 ) | ( n567 & n569 ) ;
  assign n597 = n595 | n596 ;
  assign n598 = ~x7 & n303 ;
  assign n599 = n597 & n598 ;
  assign n600 = ~n553 & n568 ;
  assign n601 = ( ~x7 & n598 ) | ( ~x7 & n600 ) | ( n598 & n600 ) ;
  assign n602 = n597 ^ n595 ^ n567 ;
  assign n603 = n598 & n602 ;
  assign n604 = x4 & n533 ;
  assign n605 = ( n533 & n601 ) | ( n533 & ~n604 ) | ( n601 & ~n604 ) ;
  assign n606 = ( x2 & n567 ) | ( x2 & n600 ) | ( n567 & n600 ) ;
  assign n607 = ( n443 & n600 ) | ( n443 & n606 ) | ( n600 & n606 ) ;
  assign n608 = ( ~x7 & n600 ) | ( ~x7 & n607 ) | ( n600 & n607 ) ;
  assign n609 = ( ~x7 & n327 ) | ( ~x7 & n608 ) | ( n327 & n608 ) ;
  assign n610 = ~n327 & n609 ;
  assign y0 = ~n564 ;
  assign y1 = n548 ;
  assign y2 = n581 ;
  assign y3 = n594 ;
  assign y4 = n599 ;
  assign y5 = n603 ;
  assign y6 = ~n605 ;
  assign y7 = n481 ;
  assign y8 = n459 ;
  assign y9 = n342 ;
  assign y10 = n610 ;
endmodule
