module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 ;
  assign n129 = x105 | x106 ;
  assign n130 = x117 | x118 ;
  assign n131 = x119 | x120 ;
  assign n132 = n130 | n131 ;
  assign n133 = x113 | x114 ;
  assign n134 = n132 | n133 ;
  assign n135 = x107 | x108 ;
  assign n136 = x85 | x86 ;
  assign n137 = x87 | x88 ;
  assign n138 = x109 | x110 ;
  assign n139 = n136 | n137 ;
  assign n140 = x101 | x102 ;
  assign n141 = x93 | x94 ;
  assign n142 = x122 | x123 ;
  assign n143 = x95 | x96 ;
  assign n144 = x88 | x91 ;
  assign n145 = x115 | x116 ;
  assign n146 = x91 | x92 ;
  assign n147 = x126 | x127 ;
  assign n148 = x97 | x98 ;
  assign n149 = x99 | x100 ;
  assign n150 = x92 | x95 ;
  assign n151 = n129 | n135 ;
  assign n152 = x89 | x90 ;
  assign n153 = x125 | n147 ;
  assign n154 = x124 | n153 ;
  assign n155 = n142 | n154 ;
  assign n156 = x121 | n155 ;
  assign n157 = ( ~n134 & n145 ) | ( ~n134 & n156 ) | ( n145 & n156 ) ;
  assign n158 = n134 | n157 ;
  assign n159 = x111 | x112 ;
  assign n160 = n138 | n159 ;
  assign n161 = n151 | n160 ;
  assign n162 = n158 | n161 ;
  assign n163 = x120 | n156 ;
  assign n164 = x103 | x104 ;
  assign n165 = x84 | x87 ;
  assign n166 = n136 | n165 ;
  assign n167 = n140 | n164 ;
  assign n168 = n162 | n167 ;
  assign n169 = x35 & x64 ;
  assign n170 = x116 | x119 ;
  assign n171 = n132 | n156 ;
  assign n172 = x112 | x115 ;
  assign n173 = ( ~n130 & n163 ) | ( ~n130 & n170 ) | ( n163 & n170 ) ;
  assign n174 = n130 | n173 ;
  assign n175 = n141 | n143 ;
  assign n176 = n158 | n160 ;
  assign n177 = n135 | n176 ;
  assign n178 = n146 | n152 ;
  assign n179 = n175 | n178 ;
  assign n180 = ( ~x63 & x64 ) | ( ~x63 & x65 ) | ( x64 & x65 ) ;
  assign n181 = ( ~n133 & n172 ) | ( ~n133 & n174 ) | ( n172 & n174 ) ;
  assign n182 = n145 | n171 ;
  assign n183 = n133 | n181 ;
  assign n184 = n141 | n150 ;
  assign n185 = ( ~x65 & x66 ) | ( ~x65 & n180 ) | ( x66 & n180 ) ;
  assign n186 = ( ~x104 & x107 ) | ( ~x104 & n129 ) | ( x107 & n129 ) ;
  assign n187 = ( ~x100 & x103 ) | ( ~x100 & n140 ) | ( x103 & n140 ) ;
  assign n188 = x100 | n187 ;
  assign n189 = x104 | n186 ;
  assign n190 = x65 | n185 ;
  assign n191 = n149 | n167 ;
  assign n192 = ( ~x108 & x111 ) | ( ~x108 & n138 ) | ( x111 & n138 ) ;
  assign n193 = x108 | n192 ;
  assign n194 = n189 | n193 ;
  assign n195 = n139 | n179 ;
  assign n196 = ( ~x96 & x99 ) | ( ~x96 & n148 ) | ( x99 & n148 ) ;
  assign n197 = n148 | n149 ;
  assign n198 = n188 | n194 ;
  assign n199 = n183 | n198 ;
  assign n200 = ( ~n141 & n169 ) | ( ~n141 & n199 ) | ( n169 & n199 ) ;
  assign n201 = n144 | n152 ;
  assign n202 = n168 | n197 ;
  assign n203 = n179 | n202 ;
  assign n204 = n137 | n203 ;
  assign n205 = ~x62 & x64 ;
  assign n206 = x96 | n196 ;
  assign n207 = n198 | n206 ;
  assign n208 = ~n199 & n200 ;
  assign n209 = x76 | x77 ;
  assign n210 = x78 | x79 ;
  assign n211 = x74 | x75 ;
  assign n212 = x66 | x67 ;
  assign n213 = n209 | n210 ;
  assign n214 = x68 | x69 ;
  assign n215 = x70 | x71 ;
  assign n216 = x81 | x82 ;
  assign n217 = x72 | x73 ;
  assign n218 = n211 | n217 ;
  assign n219 = n213 | n218 ;
  assign n220 = n214 | n215 ;
  assign n221 = n212 | n220 ;
  assign n222 = x80 | x83 ;
  assign n223 = n216 | n222 ;
  assign n224 = n166 | n223 ;
  assign n225 = n184 | n201 ;
  assign n226 = n183 & ~n207 ;
  assign n227 = ( x64 & ~x65 ) | ( x64 & n207 ) | ( ~x65 & n207 ) ;
  assign n228 = n224 | n225 ;
  assign n229 = n219 | n228 ;
  assign n230 = ( ~n207 & n221 ) | ( ~n207 & n229 ) | ( n221 & n229 ) ;
  assign n231 = ( n207 & n227 ) | ( n207 & ~n230 ) | ( n227 & ~n230 ) ;
  assign n232 = ( n207 & ~n226 ) | ( n207 & n231 ) | ( ~n226 & n231 ) ;
  assign n233 = ( x65 & n205 ) | ( x65 & n225 ) | ( n205 & n225 ) ;
  assign n234 = ( x65 & n205 ) | ( x65 & ~n207 ) | ( n205 & ~n207 ) ;
  assign n235 = n219 | n224 ;
  assign n236 = ( ~n183 & n233 ) | ( ~n183 & n234 ) | ( n233 & n234 ) ;
  assign n237 = ~n233 & n236 ;
  assign n238 = ( ~n221 & n235 ) | ( ~n221 & n237 ) | ( n235 & n237 ) ;
  assign n239 = ( x63 & n207 ) | ( x63 & ~n232 ) | ( n207 & ~n232 ) ;
  assign n240 = n219 | n221 ;
  assign n241 = n235 & n239 ;
  assign n242 = ( x65 & n205 ) | ( x65 & ~n239 ) | ( n205 & ~n239 ) ;
  assign n243 = n183 | n207 ;
  assign n244 = n238 & ~n242 ;
  assign n245 = n229 | n243 ;
  assign n246 = ( n239 & n241 ) | ( n239 & ~n244 ) | ( n241 & ~n244 ) ;
  assign n247 = n206 | n225 ;
  assign n248 = n220 | n245 ;
  assign n249 = n166 | n247 ;
  assign n250 = n220 | n249 ;
  assign n251 = n219 | n223 ;
  assign n252 = ( n199 & ~n250 ) | ( n199 & n251 ) | ( ~n250 & n251 ) ;
  assign n253 = n250 | n252 ;
  assign n254 = n199 | n249 ;
  assign n255 = ( ~x69 & x72 ) | ( ~x69 & n215 ) | ( x72 & n215 ) ;
  assign n256 = x62 & ~x64 ;
  assign n257 = x69 | n255 ;
  assign n258 = x67 | x68 ;
  assign n259 = n257 | n258 ;
  assign n260 = ~x61 & x64 ;
  assign n261 = ( x62 & x66 ) | ( x62 & n202 ) | ( x66 & n202 ) ;
  assign n262 = x83 | x84 ;
  assign n263 = n216 | n262 ;
  assign n264 = n195 | n263 ;
  assign n265 = ( ~x77 & x80 ) | ( ~x77 & n210 ) | ( x80 & n210 ) ;
  assign n266 = x77 | n265 ;
  assign n267 = x73 | x76 ;
  assign n268 = ( ~n211 & n266 ) | ( ~n211 & n267 ) | ( n266 & n267 ) ;
  assign n269 = n211 | n268 ;
  assign n270 = n259 | n269 ;
  assign n271 = n264 | n270 ;
  assign n272 = ( x62 & n242 ) | ( x62 & n271 ) | ( n242 & n271 ) ;
  assign n273 = ( x62 & n261 ) | ( x62 & n272 ) | ( n261 & n272 ) ;
  assign n274 = ( x62 & n256 ) | ( x62 & n273 ) | ( n256 & n273 ) ;
  assign n275 = ( x65 & n260 ) | ( x65 & ~n274 ) | ( n260 & ~n274 ) ;
  assign n276 = ( x66 & ~n246 ) | ( x66 & n275 ) | ( ~n246 & n275 ) ;
  assign n277 = n228 | n243 ;
  assign n278 = ( n240 & ~n242 ) | ( n240 & n277 ) | ( ~n242 & n277 ) ;
  assign n279 = n242 | n278 ;
  assign n280 = n215 | n218 ;
  assign n281 = ( ~n202 & n271 ) | ( ~n202 & n276 ) | ( n271 & n276 ) ;
  assign n282 = n202 | n281 ;
  assign n283 = n246 & n282 ;
  assign n284 = ( ~x66 & n246 ) | ( ~x66 & n283 ) | ( n246 & n283 ) ;
  assign n285 = ( ~n275 & n283 ) | ( ~n275 & n284 ) | ( n283 & n284 ) ;
  assign n286 = n202 | n264 ;
  assign n287 = ( x65 & n260 ) | ( x65 & ~n286 ) | ( n260 & ~n286 ) ;
  assign n288 = ( x65 & n260 ) | ( x65 & n276 ) | ( n260 & n276 ) ;
  assign n289 = ( ~n270 & n287 ) | ( ~n270 & n288 ) | ( n287 & n288 ) ;
  assign n290 = ~n288 & n289 ;
  assign n291 = x61 & x64 ;
  assign n292 = n260 & ~n286 ;
  assign n293 = ( ~n270 & n276 ) | ( ~n270 & n292 ) | ( n276 & n292 ) ;
  assign n294 = n274 & ~n290 ;
  assign n295 = n290 ^ n274 ^ 1'b0 ;
  assign n296 = x67 | n276 ;
  assign n297 = ~n248 & n291 ;
  assign n298 = ~n296 & n297 ;
  assign n299 = ~n276 & n293 ;
  assign n300 = ( x61 & ~n298 ) | ( x61 & n299 ) | ( ~n298 & n299 ) ;
  assign n301 = n269 | n286 ;
  assign n302 = x66 & ~n294 ;
  assign n303 = n257 | n301 ;
  assign n304 = ( n190 & ~n258 ) | ( n190 & n303 ) | ( ~n258 & n303 ) ;
  assign n305 = n258 | n304 ;
  assign n306 = ~x60 & x64 ;
  assign n307 = ~x66 & n295 ;
  assign n308 = ( x65 & ~n300 ) | ( x65 & n306 ) | ( ~n300 & n306 ) ;
  assign n309 = ( n302 & ~n307 ) | ( n302 & n308 ) | ( ~n307 & n308 ) ;
  assign n310 = ( x67 & ~n285 ) | ( x67 & n309 ) | ( ~n285 & n309 ) ;
  assign n311 = n306 ^ x65 ^ 1'b0 ;
  assign n312 = ~n253 & n311 ;
  assign n313 = ( n248 & n306 ) | ( n248 & ~n310 ) | ( n306 & ~n310 ) ;
  assign n314 = n253 | n310 ;
  assign n315 = ~n248 & n313 ;
  assign n316 = n309 ^ n308 ^ n302 ;
  assign n317 = n285 & n314 ;
  assign n318 = n295 & n314 ;
  assign n319 = ( ~x66 & n295 ) | ( ~x66 & n318 ) | ( n295 & n318 ) ;
  assign n320 = ~x67 & n285 ;
  assign n321 = ( n253 & ~n309 ) | ( n253 & n320 ) | ( ~n309 & n320 ) ;
  assign n322 = ~n253 & n321 ;
  assign n323 = n310 & n312 ;
  assign n324 = ( ~n316 & n318 ) | ( ~n316 & n319 ) | ( n318 & n319 ) ;
  assign n325 = n323 ^ n312 ^ n300 ;
  assign n326 = ( n302 & n308 ) | ( n302 & ~n316 ) | ( n308 & ~n316 ) ;
  assign n327 = ( n310 & n316 ) | ( n310 & ~n324 ) | ( n316 & ~n324 ) ;
  assign n328 = x67 & ~n324 ;
  assign n329 = ~x59 & x64 ;
  assign n330 = ~x66 & n325 ;
  assign n331 = n330 ^ n325 ^ x66 ;
  assign n332 = ( x64 & x68 ) | ( x64 & ~n303 ) | ( x68 & ~n303 ) ;
  assign n333 = ~x68 & n332 ;
  assign n334 = ( x60 & n310 ) | ( x60 & ~n333 ) | ( n310 & ~n333 ) ;
  assign n335 = ~x60 & n334 ;
  assign n336 = ( n315 & n334 ) | ( n315 & ~n335 ) | ( n334 & ~n335 ) ;
  assign n337 = ( x65 & n329 ) | ( x65 & ~n336 ) | ( n329 & ~n336 ) ;
  assign n338 = n331 | n337 ;
  assign n339 = ( n324 & n326 ) | ( n324 & ~n327 ) | ( n326 & ~n327 ) ;
  assign n340 = ~n330 & n338 ;
  assign n341 = n253 & ~n324 ;
  assign n342 = ( n324 & n339 ) | ( n324 & ~n341 ) | ( n339 & ~n341 ) ;
  assign n343 = n328 | n340 ;
  assign n344 = ~x67 & n342 ;
  assign n345 = ( n328 & n340 ) | ( n328 & n344 ) | ( n340 & n344 ) ;
  assign n346 = n317 | n322 ;
  assign n347 = n343 & ~n344 ;
  assign n348 = ~n303 & n343 ;
  assign n349 = ( x68 & ~n317 ) | ( x68 & n347 ) | ( ~n317 & n347 ) ;
  assign n350 = ( x68 & ~n346 ) | ( x68 & n349 ) | ( ~n346 & n349 ) ;
  assign n351 = ~n345 & n348 ;
  assign n352 = ( n330 & n331 ) | ( n330 & n337 ) | ( n331 & n337 ) ;
  assign n353 = n303 | n350 ;
  assign n354 = n342 & n353 ;
  assign n355 = ( ~x67 & n342 ) | ( ~x67 & n354 ) | ( n342 & n354 ) ;
  assign n356 = ( ~n345 & n354 ) | ( ~n345 & n355 ) | ( n354 & n355 ) ;
  assign n357 = n350 & n351 ;
  assign n358 = n329 ^ x65 ^ 1'b0 ;
  assign n359 = ( n351 & n356 ) | ( n351 & ~n357 ) | ( n356 & ~n357 ) ;
  assign n360 = n353 & n358 ;
  assign n361 = n360 ^ n358 ^ n336 ;
  assign n362 = n325 & n353 ;
  assign n363 = ~n303 & n338 ;
  assign n364 = n213 | n223 ;
  assign n365 = ( ~x66 & n325 ) | ( ~x66 & n362 ) | ( n325 & n362 ) ;
  assign n366 = n254 | n364 ;
  assign n367 = n280 | n366 ;
  assign n368 = ~n352 & n363 ;
  assign n369 = ( ~n352 & n362 ) | ( ~n352 & n365 ) | ( n362 & n365 ) ;
  assign n370 = n346 & n353 ;
  assign n371 = n329 & ~n353 ;
  assign n372 = ( n303 & n346 ) | ( n303 & ~n347 ) | ( n346 & ~n347 ) ;
  assign n373 = x64 & ~x71 ;
  assign n374 = ( ~x68 & n346 ) | ( ~x68 & n370 ) | ( n346 & n370 ) ;
  assign n375 = ( ~n218 & n364 ) | ( ~n218 & n373 ) | ( n364 & n373 ) ;
  assign n376 = n350 & n368 ;
  assign n377 = ( n370 & n372 ) | ( n370 & n374 ) | ( n372 & n374 ) ;
  assign n378 = x69 | n350 ;
  assign n379 = ~n366 & n375 ;
  assign n380 = ~x58 & x64 ;
  assign n381 = x59 & x64 ;
  assign n382 = ~n367 & n381 ;
  assign n383 = ~n378 & n382 ;
  assign n384 = ( x59 & n371 ) | ( x59 & ~n383 ) | ( n371 & ~n383 ) ;
  assign n385 = n384 ^ n380 ^ x65 ;
  assign n386 = ( x65 & n380 ) | ( x65 & n385 ) | ( n380 & n385 ) ;
  assign n387 = n386 ^ n361 ^ x66 ;
  assign n388 = ( n368 & n369 ) | ( n368 & ~n376 ) | ( n369 & ~n376 ) ;
  assign n389 = ( x69 & n367 ) | ( x69 & ~n377 ) | ( n367 & ~n377 ) ;
  assign n390 = ( x66 & n386 ) | ( x66 & n387 ) | ( n386 & n387 ) ;
  assign n391 = n303 & n377 ;
  assign n392 = ( x67 & ~n388 ) | ( x67 & n390 ) | ( ~n388 & n390 ) ;
  assign n393 = ( x68 & ~n359 ) | ( x68 & n392 ) | ( ~n359 & n392 ) ;
  assign n394 = ( ~x69 & n377 ) | ( ~x69 & n393 ) | ( n377 & n393 ) ;
  assign n395 = n389 | n394 ;
  assign n396 = ( ~n377 & n391 ) | ( ~n377 & n395 ) | ( n391 & n395 ) ;
  assign n397 = n396 ^ n387 ^ 1'b0 ;
  assign n398 = ( n361 & n387 ) | ( n361 & n397 ) | ( n387 & n397 ) ;
  assign n399 = n396 ^ n385 ^ 1'b0 ;
  assign n400 = ( n384 & n385 ) | ( n384 & n399 ) | ( n385 & n399 ) ;
  assign n401 = n391 & ~n395 ;
  assign n402 = ( n322 & n391 ) | ( n322 & ~n401 ) | ( n391 & ~n401 ) ;
  assign n403 = n392 ^ n359 ^ x68 ;
  assign n404 = n390 ^ n388 ^ x67 ;
  assign n405 = n396 ^ n388 ^ 1'b0 ;
  assign n406 = ( n388 & n404 ) | ( n388 & ~n405 ) | ( n404 & ~n405 ) ;
  assign n407 = n396 ^ n359 ^ 1'b0 ;
  assign n408 = ( n359 & n403 ) | ( n359 & ~n407 ) | ( n403 & ~n407 ) ;
  assign n409 = ~x57 & x64 ;
  assign n410 = x71 | x72 ;
  assign n411 = x64 & n396 ;
  assign n412 = n411 ^ x64 ^ x58 ;
  assign n413 = n412 ^ n409 ^ x65 ;
  assign n414 = ( x65 & n409 ) | ( x65 & n413 ) | ( n409 & n413 ) ;
  assign n415 = n414 ^ n400 ^ x66 ;
  assign n416 = ( x66 & n414 ) | ( x66 & n415 ) | ( n414 & n415 ) ;
  assign n417 = ( x67 & ~n398 ) | ( x67 & n416 ) | ( ~n398 & n416 ) ;
  assign n418 = ( x68 & ~n406 ) | ( x68 & n417 ) | ( ~n406 & n417 ) ;
  assign n419 = ( x69 & ~n408 ) | ( x69 & n418 ) | ( ~n408 & n418 ) ;
  assign n420 = ( x70 & ~n402 ) | ( x70 & n419 ) | ( ~n402 & n419 ) ;
  assign n421 = ( ~n301 & n410 ) | ( ~n301 & n420 ) | ( n410 & n420 ) ;
  assign n422 = n301 | n421 ;
  assign n423 = ( n322 & n402 ) | ( n322 & n422 ) | ( n402 & n422 ) ;
  assign n424 = ~x56 & x64 ;
  assign n425 = n422 ^ n415 ^ 1'b0 ;
  assign n426 = ( n400 & n415 ) | ( n400 & n425 ) | ( n415 & n425 ) ;
  assign n427 = n418 ^ n408 ^ x69 ;
  assign n428 = n422 ^ n406 ^ 1'b0 ;
  assign n429 = ~n218 & n424 ;
  assign n430 = ( x57 & ~n379 ) | ( x57 & n420 ) | ( ~n379 & n420 ) ;
  assign n431 = n427 ^ n422 ^ 1'b0 ;
  assign n432 = ( n408 & n427 ) | ( n408 & n431 ) | ( n427 & n431 ) ;
  assign n433 = n409 & ~n422 ;
  assign n434 = x57 & ~n430 ;
  assign n435 = ( x57 & n433 ) | ( x57 & ~n434 ) | ( n433 & ~n434 ) ;
  assign n436 = n422 ^ n413 ^ 1'b0 ;
  assign n437 = n435 ^ n424 ^ x65 ;
  assign n438 = n422 ^ n398 ^ 1'b0 ;
  assign n439 = n416 ^ n398 ^ x67 ;
  assign n440 = ( x65 & n424 ) | ( x65 & n437 ) | ( n424 & n437 ) ;
  assign n441 = ( n412 & n413 ) | ( n412 & n436 ) | ( n413 & n436 ) ;
  assign n442 = n441 ^ n440 ^ x66 ;
  assign n443 = ( n398 & ~n438 ) | ( n398 & n439 ) | ( ~n438 & n439 ) ;
  assign n444 = n417 ^ n406 ^ x68 ;
  assign n445 = ( n406 & ~n428 ) | ( n406 & n444 ) | ( ~n428 & n444 ) ;
  assign n446 = ( x66 & n440 ) | ( x66 & n442 ) | ( n440 & n442 ) ;
  assign n447 = ( x67 & ~n426 ) | ( x67 & n446 ) | ( ~n426 & n446 ) ;
  assign n448 = ( x68 & ~n443 ) | ( x68 & n447 ) | ( ~n443 & n447 ) ;
  assign n449 = ( x69 & ~n445 ) | ( x69 & n448 ) | ( ~n445 & n448 ) ;
  assign n450 = ( x70 & ~n432 ) | ( x70 & n449 ) | ( ~n432 & n449 ) ;
  assign n451 = ( x71 & ~n423 ) | ( x71 & n450 ) | ( ~n423 & n450 ) ;
  assign n452 = n245 | n451 ;
  assign n453 = n448 ^ n445 ^ x69 ;
  assign n454 = n446 ^ n426 ^ x67 ;
  assign n455 = n452 ^ n437 ^ 1'b0 ;
  assign n456 = ( n435 & n437 ) | ( n435 & n455 ) | ( n437 & n455 ) ;
  assign n457 = n449 ^ n432 ^ x70 ;
  assign n458 = n452 ^ n442 ^ 1'b0 ;
  assign n459 = n457 ^ n452 ^ 1'b0 ;
  assign n460 = ( n441 & n442 ) | ( n441 & n458 ) | ( n442 & n458 ) ;
  assign n461 = n452 ^ n426 ^ 1'b0 ;
  assign n462 = n452 ^ n443 ^ 1'b0 ;
  assign n463 = ( n426 & n454 ) | ( n426 & ~n461 ) | ( n454 & ~n461 ) ;
  assign n464 = n447 ^ n443 ^ x68 ;
  assign n465 = ( n443 & ~n462 ) | ( n443 & n464 ) | ( ~n462 & n464 ) ;
  assign n466 = ( n432 & n457 ) | ( n432 & n459 ) | ( n457 & n459 ) ;
  assign n467 = n452 ^ n445 ^ 1'b0 ;
  assign n468 = ( n445 & n453 ) | ( n445 & ~n467 ) | ( n453 & ~n467 ) ;
  assign n469 = ~x55 & x64 ;
  assign n470 = n195 | n202 ;
  assign n471 = n263 | n470 ;
  assign n472 = x56 & x64 ;
  assign n473 = ( ~x72 & n451 ) | ( ~x72 & n472 ) | ( n451 & n472 ) ;
  assign n474 = ( ~n366 & n429 ) | ( ~n366 & n451 ) | ( n429 & n451 ) ;
  assign n475 = ~n451 & n474 ;
  assign n476 = n423 & n452 ;
  assign n477 = n322 | n476 ;
  assign n478 = ~n451 & n473 ;
  assign n479 = ( ~n269 & n471 ) | ( ~n269 & n478 ) | ( n471 & n478 ) ;
  assign n480 = ~n471 & n479 ;
  assign n481 = ( x56 & n475 ) | ( x56 & ~n480 ) | ( n475 & ~n480 ) ;
  assign n482 = n481 ^ n469 ^ x65 ;
  assign n483 = ( x65 & n469 ) | ( x65 & n482 ) | ( n469 & n482 ) ;
  assign n484 = n483 ^ n456 ^ x66 ;
  assign n485 = ( x66 & n483 ) | ( x66 & n484 ) | ( n483 & n484 ) ;
  assign n486 = ( x67 & ~n460 ) | ( x67 & n485 ) | ( ~n460 & n485 ) ;
  assign n487 = ( x68 & ~n463 ) | ( x68 & n486 ) | ( ~n463 & n486 ) ;
  assign n488 = ( x69 & ~n465 ) | ( x69 & n487 ) | ( ~n465 & n487 ) ;
  assign n489 = ( x70 & ~n468 ) | ( x70 & n488 ) | ( ~n468 & n488 ) ;
  assign n490 = n489 ^ n466 ^ x71 ;
  assign n491 = ( x71 & ~n466 ) | ( x71 & n489 ) | ( ~n466 & n489 ) ;
  assign n492 = ( x72 & n301 ) | ( x72 & ~n476 ) | ( n301 & ~n476 ) ;
  assign n493 = ( ~x72 & n301 ) | ( ~x72 & n477 ) | ( n301 & n477 ) ;
  assign n494 = ( ~n491 & n492 ) | ( ~n491 & n493 ) | ( n492 & n493 ) ;
  assign n495 = n491 | n494 ;
  assign n496 = n245 & n477 ;
  assign n497 = ( ~n477 & n495 ) | ( ~n477 & n496 ) | ( n495 & n496 ) ;
  assign n498 = n497 ^ n466 ^ 1'b0 ;
  assign n499 = ( n466 & n490 ) | ( n466 & ~n498 ) | ( n490 & ~n498 ) ;
  assign n500 = n488 ^ n468 ^ x70 ;
  assign n501 = n497 ^ n468 ^ 1'b0 ;
  assign n502 = ( n468 & n500 ) | ( n468 & ~n501 ) | ( n500 & ~n501 ) ;
  assign n503 = n487 ^ n465 ^ x69 ;
  assign n504 = n497 ^ n465 ^ 1'b0 ;
  assign n505 = ( n465 & n503 ) | ( n465 & ~n504 ) | ( n503 & ~n504 ) ;
  assign n506 = n486 ^ n463 ^ x68 ;
  assign n507 = n497 ^ n463 ^ 1'b0 ;
  assign n508 = ( n463 & n506 ) | ( n463 & ~n507 ) | ( n506 & ~n507 ) ;
  assign n509 = n485 ^ n460 ^ x67 ;
  assign n510 = n497 ^ n460 ^ 1'b0 ;
  assign n511 = ( n460 & n509 ) | ( n460 & ~n510 ) | ( n509 & ~n510 ) ;
  assign n512 = n497 ^ n484 ^ 1'b0 ;
  assign n513 = ( n456 & n484 ) | ( n456 & n512 ) | ( n484 & n512 ) ;
  assign n514 = n497 ^ n482 ^ 1'b0 ;
  assign n515 = ( n481 & n482 ) | ( n481 & n514 ) | ( n482 & n514 ) ;
  assign n516 = ( n245 & n322 ) | ( n245 & n423 ) | ( n322 & n423 ) ;
  assign n517 = n322 | n495 ;
  assign n518 = ( n322 & n516 ) | ( n322 & n517 ) | ( n516 & n517 ) ;
  assign n519 = x64 & n497 ;
  assign n520 = n519 ^ x64 ^ x55 ;
  assign n521 = ~x54 & x64 ;
  assign n522 = n521 ^ n520 ^ x65 ;
  assign n523 = ( x65 & n521 ) | ( x65 & n522 ) | ( n521 & n522 ) ;
  assign n524 = n523 ^ n515 ^ x66 ;
  assign n525 = ( x66 & n523 ) | ( x66 & n524 ) | ( n523 & n524 ) ;
  assign n526 = ( x67 & ~n513 ) | ( x67 & n525 ) | ( ~n513 & n525 ) ;
  assign n527 = ( x68 & ~n511 ) | ( x68 & n526 ) | ( ~n511 & n526 ) ;
  assign n528 = ( x69 & ~n508 ) | ( x69 & n527 ) | ( ~n508 & n527 ) ;
  assign n529 = ( x70 & ~n505 ) | ( x70 & n528 ) | ( ~n505 & n528 ) ;
  assign n530 = ( x71 & ~n502 ) | ( x71 & n529 ) | ( ~n502 & n529 ) ;
  assign n531 = ( x72 & ~n499 ) | ( x72 & n530 ) | ( ~n499 & n530 ) ;
  assign n532 = ( x73 & ~n518 ) | ( x73 & n531 ) | ( ~n518 & n531 ) ;
  assign n533 = x74 | n532 ;
  assign n534 = n526 ^ n511 ^ x68 ;
  assign n535 = n525 ^ n513 ^ x67 ;
  assign n536 = n211 | n213 ;
  assign n537 = n527 ^ n508 ^ x69 ;
  assign n538 = ( n277 & n532 ) | ( n277 & ~n536 ) | ( n532 & ~n536 ) ;
  assign n539 = n536 | n538 ;
  assign n540 = x75 | x76 ;
  assign n541 = ( ~n266 & n286 ) | ( ~n266 & n540 ) | ( n286 & n540 ) ;
  assign n542 = n530 ^ n499 ^ x72 ;
  assign n543 = n266 | n541 ;
  assign n544 = n542 ^ n539 ^ 1'b0 ;
  assign n545 = ( n499 & n542 ) | ( n499 & n544 ) | ( n542 & n544 ) ;
  assign n546 = n528 ^ n505 ^ x70 ;
  assign n547 = n539 ^ n511 ^ 1'b0 ;
  assign n548 = ( n511 & n534 ) | ( n511 & ~n547 ) | ( n534 & ~n547 ) ;
  assign n549 = x54 & x64 ;
  assign n550 = ~n543 & n549 ;
  assign n551 = ~n533 & n550 ;
  assign n552 = ~x53 & x64 ;
  assign n553 = n529 ^ n502 ^ x71 ;
  assign n554 = n539 ^ n513 ^ 1'b0 ;
  assign n555 = n539 ^ n505 ^ 1'b0 ;
  assign n556 = ( n513 & n535 ) | ( n513 & ~n554 ) | ( n535 & ~n554 ) ;
  assign n557 = ( n505 & n546 ) | ( n505 & ~n555 ) | ( n546 & ~n555 ) ;
  assign n558 = n521 & ~n539 ;
  assign n559 = ( x54 & ~n551 ) | ( x54 & n558 ) | ( ~n551 & n558 ) ;
  assign n560 = n559 ^ n552 ^ x65 ;
  assign n561 = n539 ^ n522 ^ 1'b0 ;
  assign n562 = ( n520 & n522 ) | ( n520 & n561 ) | ( n522 & n561 ) ;
  assign n563 = ( n322 & n518 ) | ( n322 & n539 ) | ( n518 & n539 ) ;
  assign n564 = n539 ^ n524 ^ 1'b0 ;
  assign n565 = ( x65 & n552 ) | ( x65 & n560 ) | ( n552 & n560 ) ;
  assign n566 = n565 ^ n562 ^ x66 ;
  assign n567 = ( x66 & n565 ) | ( x66 & n566 ) | ( n565 & n566 ) ;
  assign n568 = n539 ^ n508 ^ 1'b0 ;
  assign n569 = ( n515 & n524 ) | ( n515 & n564 ) | ( n524 & n564 ) ;
  assign n570 = ( x67 & n567 ) | ( x67 & ~n569 ) | ( n567 & ~n569 ) ;
  assign n571 = ( n508 & n537 ) | ( n508 & ~n568 ) | ( n537 & ~n568 ) ;
  assign n572 = ( x68 & ~n556 ) | ( x68 & n570 ) | ( ~n556 & n570 ) ;
  assign n573 = ( x69 & ~n548 ) | ( x69 & n572 ) | ( ~n548 & n572 ) ;
  assign n574 = ( x70 & ~n571 ) | ( x70 & n573 ) | ( ~n571 & n573 ) ;
  assign n575 = ( x71 & ~n557 ) | ( x71 & n574 ) | ( ~n557 & n574 ) ;
  assign n576 = n539 ^ n502 ^ 1'b0 ;
  assign n577 = ( n502 & n553 ) | ( n502 & ~n576 ) | ( n553 & ~n576 ) ;
  assign n578 = ( x72 & n575 ) | ( x72 & ~n577 ) | ( n575 & ~n577 ) ;
  assign n579 = ( x73 & ~n545 ) | ( x73 & n578 ) | ( ~n545 & n578 ) ;
  assign n580 = ( x74 & ~n563 ) | ( x74 & n579 ) | ( ~n563 & n579 ) ;
  assign n581 = ( x64 & ~x75 ) | ( x64 & n580 ) | ( ~x75 & n580 ) ;
  assign n582 = ( ~n213 & n228 ) | ( ~n213 & n581 ) | ( n228 & n581 ) ;
  assign n583 = n572 ^ n548 ^ x69 ;
  assign n584 = n277 & ~n580 ;
  assign n585 = n543 | n580 ;
  assign n586 = n552 | n585 ;
  assign n587 = ( n580 & n582 ) | ( n580 & ~n584 ) | ( n582 & ~n584 ) ;
  assign n588 = n585 ^ n548 ^ 1'b0 ;
  assign n589 = n577 ^ n575 ^ x72 ;
  assign n590 = ( n548 & n583 ) | ( n548 & ~n588 ) | ( n583 & ~n588 ) ;
  assign n591 = n585 ^ n566 ^ 1'b0 ;
  assign n592 = ( n562 & n566 ) | ( n562 & n591 ) | ( n566 & n591 ) ;
  assign n593 = n585 ^ n560 ^ 1'b0 ;
  assign n594 = n585 ^ n577 ^ 1'b0 ;
  assign n595 = ( x53 & n580 ) | ( x53 & ~n587 ) | ( n580 & ~n587 ) ;
  assign n596 = ( ~n585 & n586 ) | ( ~n585 & n595 ) | ( n586 & n595 ) ;
  assign n597 = ( n577 & n589 ) | ( n577 & ~n594 ) | ( n589 & ~n594 ) ;
  assign n598 = ( n559 & n560 ) | ( n559 & n593 ) | ( n560 & n593 ) ;
  assign n599 = n578 ^ n545 ^ x73 ;
  assign n600 = n599 ^ n585 ^ 1'b0 ;
  assign n601 = ( n545 & n599 ) | ( n545 & n600 ) | ( n599 & n600 ) ;
  assign n602 = n574 ^ n557 ^ x71 ;
  assign n603 = n573 ^ n571 ^ x70 ;
  assign n604 = n585 ^ n571 ^ 1'b0 ;
  assign n605 = ( n571 & n603 ) | ( n571 & ~n604 ) | ( n603 & ~n604 ) ;
  assign n606 = n570 ^ n556 ^ x68 ;
  assign n607 = n585 ^ n556 ^ 1'b0 ;
  assign n608 = ( n556 & n606 ) | ( n556 & ~n607 ) | ( n606 & ~n607 ) ;
  assign n609 = n569 ^ n567 ^ x67 ;
  assign n610 = n585 ^ n557 ^ 1'b0 ;
  assign n611 = ( n557 & n602 ) | ( n557 & ~n610 ) | ( n602 & ~n610 ) ;
  assign n612 = n585 ^ n569 ^ 1'b0 ;
  assign n613 = ( n569 & n609 ) | ( n569 & ~n612 ) | ( n609 & ~n612 ) ;
  assign n614 = ~x52 & x64 ;
  assign n615 = n614 ^ n596 ^ x65 ;
  assign n616 = ( x65 & n614 ) | ( x65 & n615 ) | ( n614 & n615 ) ;
  assign n617 = n616 ^ n598 ^ x66 ;
  assign n618 = ( x66 & n616 ) | ( x66 & n617 ) | ( n616 & n617 ) ;
  assign n619 = ( x67 & ~n592 ) | ( x67 & n618 ) | ( ~n592 & n618 ) ;
  assign n620 = ( x68 & ~n613 ) | ( x68 & n619 ) | ( ~n613 & n619 ) ;
  assign n621 = ( x69 & ~n608 ) | ( x69 & n620 ) | ( ~n608 & n620 ) ;
  assign n622 = ( x70 & ~n590 ) | ( x70 & n621 ) | ( ~n590 & n621 ) ;
  assign n623 = ( x71 & ~n605 ) | ( x71 & n622 ) | ( ~n605 & n622 ) ;
  assign n624 = ( x72 & ~n611 ) | ( x72 & n623 ) | ( ~n611 & n623 ) ;
  assign n625 = ( x73 & ~n597 ) | ( x73 & n624 ) | ( ~n597 & n624 ) ;
  assign n626 = n625 ^ n601 ^ x74 ;
  assign n627 = n563 & n585 ;
  assign n628 = n322 | n627 ;
  assign n629 = ( x74 & ~n601 ) | ( x74 & n625 ) | ( ~n601 & n625 ) ;
  assign n630 = ( x75 & n366 ) | ( x75 & ~n627 ) | ( n366 & ~n627 ) ;
  assign n631 = ( ~x75 & n366 ) | ( ~x75 & n628 ) | ( n366 & n628 ) ;
  assign n632 = ( ~n629 & n630 ) | ( ~n629 & n631 ) | ( n630 & n631 ) ;
  assign n633 = n629 | n632 ;
  assign n634 = n543 & n628 ;
  assign n635 = ( ~n628 & n633 ) | ( ~n628 & n634 ) | ( n633 & n634 ) ;
  assign n636 = n635 ^ n601 ^ 1'b0 ;
  assign n637 = ( n601 & n626 ) | ( n601 & ~n636 ) | ( n626 & ~n636 ) ;
  assign n638 = n624 ^ n597 ^ x73 ;
  assign n639 = n635 ^ n597 ^ 1'b0 ;
  assign n640 = ( n597 & n638 ) | ( n597 & ~n639 ) | ( n638 & ~n639 ) ;
  assign n641 = n623 ^ n611 ^ x72 ;
  assign n642 = n635 ^ n611 ^ 1'b0 ;
  assign n643 = ( n611 & n641 ) | ( n611 & ~n642 ) | ( n641 & ~n642 ) ;
  assign n644 = n622 ^ n605 ^ x71 ;
  assign n645 = n635 ^ n605 ^ 1'b0 ;
  assign n646 = ( n605 & n644 ) | ( n605 & ~n645 ) | ( n644 & ~n645 ) ;
  assign n647 = n621 ^ n590 ^ x70 ;
  assign n648 = n635 ^ n590 ^ 1'b0 ;
  assign n649 = ( n590 & n647 ) | ( n590 & ~n648 ) | ( n647 & ~n648 ) ;
  assign n650 = n620 ^ n608 ^ x69 ;
  assign n651 = n635 ^ n608 ^ 1'b0 ;
  assign n652 = ( n608 & n650 ) | ( n608 & ~n651 ) | ( n650 & ~n651 ) ;
  assign n653 = n619 ^ n613 ^ x68 ;
  assign n654 = n635 ^ n613 ^ 1'b0 ;
  assign n655 = ( n613 & n653 ) | ( n613 & ~n654 ) | ( n653 & ~n654 ) ;
  assign n656 = n618 ^ n592 ^ x67 ;
  assign n657 = n635 ^ n592 ^ 1'b0 ;
  assign n658 = ( n592 & n656 ) | ( n592 & ~n657 ) | ( n656 & ~n657 ) ;
  assign n659 = n635 ^ n617 ^ 1'b0 ;
  assign n660 = ( n598 & n617 ) | ( n598 & n659 ) | ( n617 & n659 ) ;
  assign n661 = n635 ^ n615 ^ 1'b0 ;
  assign n662 = ( n596 & n615 ) | ( n596 & n661 ) | ( n615 & n661 ) ;
  assign n663 = ( n322 & n563 ) | ( n322 & n633 ) | ( n563 & n633 ) ;
  assign n664 = n322 | n543 ;
  assign n665 = ( n322 & n663 ) | ( n322 & n664 ) | ( n663 & n664 ) ;
  assign n666 = ( ~n210 & n223 ) | ( ~n210 & n254 ) | ( n223 & n254 ) ;
  assign n667 = n210 | n666 ;
  assign n668 = ~x51 & x64 ;
  assign n669 = x64 & n635 ;
  assign n670 = n669 ^ x64 ^ x52 ;
  assign n671 = n670 ^ n668 ^ x65 ;
  assign n672 = ( x65 & n668 ) | ( x65 & n671 ) | ( n668 & n671 ) ;
  assign n673 = n672 ^ n662 ^ x66 ;
  assign n674 = ( x66 & n672 ) | ( x66 & n673 ) | ( n672 & n673 ) ;
  assign n675 = ( x67 & ~n660 ) | ( x67 & n674 ) | ( ~n660 & n674 ) ;
  assign n676 = ( x68 & ~n658 ) | ( x68 & n675 ) | ( ~n658 & n675 ) ;
  assign n677 = ( x69 & ~n655 ) | ( x69 & n676 ) | ( ~n655 & n676 ) ;
  assign n678 = ( x70 & ~n652 ) | ( x70 & n677 ) | ( ~n652 & n677 ) ;
  assign n679 = ( x71 & ~n649 ) | ( x71 & n678 ) | ( ~n649 & n678 ) ;
  assign n680 = ( x72 & ~n646 ) | ( x72 & n679 ) | ( ~n646 & n679 ) ;
  assign n681 = ( x73 & ~n643 ) | ( x73 & n680 ) | ( ~n643 & n680 ) ;
  assign n682 = ( x74 & ~n640 ) | ( x74 & n681 ) | ( ~n640 & n681 ) ;
  assign n683 = ( x75 & ~n637 ) | ( x75 & n682 ) | ( ~n637 & n682 ) ;
  assign n684 = ( x76 & ~n665 ) | ( x76 & n683 ) | ( ~n665 & n683 ) ;
  assign n685 = ( ~n266 & n471 ) | ( ~n266 & n684 ) | ( n471 & n684 ) ;
  assign n686 = n266 | n685 ;
  assign n687 = n674 ^ n660 ^ x67 ;
  assign n688 = ~n286 & n668 ;
  assign n689 = n679 ^ n646 ^ x72 ;
  assign n690 = n677 ^ n652 ^ x70 ;
  assign n691 = ( ~n266 & n684 ) | ( ~n266 & n688 ) | ( n684 & n688 ) ;
  assign n692 = n686 ^ n646 ^ 1'b0 ;
  assign n693 = ( n646 & n689 ) | ( n646 & ~n692 ) | ( n689 & ~n692 ) ;
  assign n694 = n676 ^ n655 ^ x69 ;
  assign n695 = n686 ^ n671 ^ 1'b0 ;
  assign n696 = ( n670 & n671 ) | ( n670 & n695 ) | ( n671 & n695 ) ;
  assign n697 = ~n684 & n691 ;
  assign n698 = n686 ^ n660 ^ 1'b0 ;
  assign n699 = n680 ^ n643 ^ x73 ;
  assign n700 = n678 ^ n649 ^ x71 ;
  assign n701 = n675 ^ n658 ^ x68 ;
  assign n702 = n682 ^ n637 ^ x75 ;
  assign n703 = n686 ^ n643 ^ 1'b0 ;
  assign n704 = ( n322 & n665 ) | ( n322 & n686 ) | ( n665 & n686 ) ;
  assign n705 = n686 ^ n649 ^ 1'b0 ;
  assign n706 = ( n649 & n700 ) | ( n649 & ~n705 ) | ( n700 & ~n705 ) ;
  assign n707 = n681 ^ n640 ^ x74 ;
  assign n708 = ( n660 & n687 ) | ( n660 & ~n698 ) | ( n687 & ~n698 ) ;
  assign n709 = n686 ^ n640 ^ 1'b0 ;
  assign n710 = n702 ^ n686 ^ 1'b0 ;
  assign n711 = n686 ^ n673 ^ 1'b0 ;
  assign n712 = n686 ^ n658 ^ 1'b0 ;
  assign n713 = ( n662 & n673 ) | ( n662 & n711 ) | ( n673 & n711 ) ;
  assign n714 = n686 ^ n652 ^ 1'b0 ;
  assign n715 = ( n643 & n699 ) | ( n643 & ~n703 ) | ( n699 & ~n703 ) ;
  assign n716 = n686 ^ n655 ^ 1'b0 ;
  assign n717 = ( n637 & n702 ) | ( n637 & n710 ) | ( n702 & n710 ) ;
  assign n718 = ( n655 & n694 ) | ( n655 & ~n716 ) | ( n694 & ~n716 ) ;
  assign n719 = ( n640 & n707 ) | ( n640 & ~n709 ) | ( n707 & ~n709 ) ;
  assign n720 = ( n652 & n690 ) | ( n652 & ~n714 ) | ( n690 & ~n714 ) ;
  assign n721 = ( n658 & n701 ) | ( n658 & ~n712 ) | ( n701 & ~n712 ) ;
  assign n722 = x77 | n684 ;
  assign n723 = ~x50 & x64 ;
  assign n724 = x51 & x64 ;
  assign n725 = ~n667 & n724 ;
  assign n726 = ~n722 & n725 ;
  assign n727 = ( x51 & n697 ) | ( x51 & ~n726 ) | ( n697 & ~n726 ) ;
  assign n728 = n727 ^ n723 ^ x65 ;
  assign n729 = ( x65 & n723 ) | ( x65 & n728 ) | ( n723 & n728 ) ;
  assign n730 = n729 ^ n696 ^ x66 ;
  assign n731 = ( x66 & n729 ) | ( x66 & n730 ) | ( n729 & n730 ) ;
  assign n732 = ( x67 & ~n713 ) | ( x67 & n731 ) | ( ~n713 & n731 ) ;
  assign n733 = ( x68 & ~n708 ) | ( x68 & n732 ) | ( ~n708 & n732 ) ;
  assign n734 = ( x69 & ~n721 ) | ( x69 & n733 ) | ( ~n721 & n733 ) ;
  assign n735 = ( x70 & ~n718 ) | ( x70 & n734 ) | ( ~n718 & n734 ) ;
  assign n736 = ( x71 & ~n720 ) | ( x71 & n735 ) | ( ~n720 & n735 ) ;
  assign n737 = ( x72 & ~n706 ) | ( x72 & n736 ) | ( ~n706 & n736 ) ;
  assign n738 = ( x73 & ~n693 ) | ( x73 & n737 ) | ( ~n693 & n737 ) ;
  assign n739 = ( x74 & ~n715 ) | ( x74 & n738 ) | ( ~n715 & n738 ) ;
  assign n740 = ( x75 & ~n719 ) | ( x75 & n739 ) | ( ~n719 & n739 ) ;
  assign n741 = n740 ^ n717 ^ x76 ;
  assign n742 = ( x76 & ~n717 ) | ( x76 & n740 ) | ( ~n717 & n740 ) ;
  assign n743 = ( x77 & ~n704 ) | ( x77 & n742 ) | ( ~n704 & n742 ) ;
  assign n744 = n667 | n743 ;
  assign n745 = n744 ^ n741 ^ 1'b0 ;
  assign n746 = ( n717 & n741 ) | ( n717 & n745 ) | ( n741 & n745 ) ;
  assign n747 = n739 ^ n719 ^ x75 ;
  assign n748 = n744 ^ n719 ^ 1'b0 ;
  assign n749 = ( n719 & n747 ) | ( n719 & ~n748 ) | ( n747 & ~n748 ) ;
  assign n750 = n738 ^ n715 ^ x74 ;
  assign n751 = n744 ^ n715 ^ 1'b0 ;
  assign n752 = ( n715 & n750 ) | ( n715 & ~n751 ) | ( n750 & ~n751 ) ;
  assign n753 = n737 ^ n693 ^ x73 ;
  assign n754 = n744 ^ n693 ^ 1'b0 ;
  assign n755 = ( n693 & n753 ) | ( n693 & ~n754 ) | ( n753 & ~n754 ) ;
  assign n756 = n736 ^ n706 ^ x72 ;
  assign n757 = n744 ^ n706 ^ 1'b0 ;
  assign n758 = ( n706 & n756 ) | ( n706 & ~n757 ) | ( n756 & ~n757 ) ;
  assign n759 = n735 ^ n720 ^ x71 ;
  assign n760 = n744 ^ n720 ^ 1'b0 ;
  assign n761 = ( n720 & n759 ) | ( n720 & ~n760 ) | ( n759 & ~n760 ) ;
  assign n762 = n734 ^ n718 ^ x70 ;
  assign n763 = n744 ^ n718 ^ 1'b0 ;
  assign n764 = ( n718 & n762 ) | ( n718 & ~n763 ) | ( n762 & ~n763 ) ;
  assign n765 = n733 ^ n721 ^ x69 ;
  assign n766 = n744 ^ n728 ^ 1'b0 ;
  assign n767 = ( n727 & n728 ) | ( n727 & n766 ) | ( n728 & n766 ) ;
  assign n768 = ( ~x79 & x80 ) | ( ~x79 & n471 ) | ( x80 & n471 ) ;
  assign n769 = x78 | n743 ;
  assign n770 = n744 ^ n730 ^ 1'b0 ;
  assign n771 = n731 ^ n713 ^ x67 ;
  assign n772 = x50 & x64 ;
  assign n773 = x79 | n768 ;
  assign n774 = n772 & ~n773 ;
  assign n775 = ~x49 & x64 ;
  assign n776 = n744 ^ n713 ^ 1'b0 ;
  assign n777 = ( n696 & n730 ) | ( n696 & n770 ) | ( n730 & n770 ) ;
  assign n778 = ~n769 & n774 ;
  assign n779 = n723 & ~n744 ;
  assign n780 = ( x50 & ~n778 ) | ( x50 & n779 ) | ( ~n778 & n779 ) ;
  assign n781 = n780 ^ n775 ^ x65 ;
  assign n782 = ( x65 & n775 ) | ( x65 & n781 ) | ( n775 & n781 ) ;
  assign n783 = n782 ^ n767 ^ x66 ;
  assign n784 = ( x66 & n782 ) | ( x66 & n783 ) | ( n782 & n783 ) ;
  assign n785 = ( x67 & ~n777 ) | ( x67 & n784 ) | ( ~n777 & n784 ) ;
  assign n786 = n744 ^ n708 ^ 1'b0 ;
  assign n787 = ( n713 & n771 ) | ( n713 & ~n776 ) | ( n771 & ~n776 ) ;
  assign n788 = ( x68 & n785 ) | ( x68 & ~n787 ) | ( n785 & ~n787 ) ;
  assign n789 = n784 ^ n777 ^ x67 ;
  assign n790 = n732 ^ n708 ^ x68 ;
  assign n791 = ( n708 & ~n786 ) | ( n708 & n790 ) | ( ~n786 & n790 ) ;
  assign n792 = ( x69 & n788 ) | ( x69 & ~n791 ) | ( n788 & ~n791 ) ;
  assign n793 = n791 ^ n788 ^ x69 ;
  assign n794 = n744 ^ n721 ^ 1'b0 ;
  assign n795 = ( n721 & n765 ) | ( n721 & ~n794 ) | ( n765 & ~n794 ) ;
  assign n796 = ( x70 & n792 ) | ( x70 & ~n795 ) | ( n792 & ~n795 ) ;
  assign n797 = ( x71 & ~n764 ) | ( x71 & n796 ) | ( ~n764 & n796 ) ;
  assign n798 = ( x72 & ~n761 ) | ( x72 & n797 ) | ( ~n761 & n797 ) ;
  assign n799 = ( x73 & ~n758 ) | ( x73 & n798 ) | ( ~n758 & n798 ) ;
  assign n800 = n787 ^ n785 ^ x68 ;
  assign n801 = n797 ^ n761 ^ x72 ;
  assign n802 = n796 ^ n764 ^ x71 ;
  assign n803 = n798 ^ n758 ^ x73 ;
  assign n804 = n795 ^ n792 ^ x70 ;
  assign n805 = ( x74 & ~n755 ) | ( x74 & n799 ) | ( ~n755 & n799 ) ;
  assign n806 = ( x75 & ~n752 ) | ( x75 & n805 ) | ( ~n752 & n805 ) ;
  assign n807 = ( x76 & ~n749 ) | ( x76 & n806 ) | ( ~n749 & n806 ) ;
  assign n808 = n807 ^ n746 ^ x77 ;
  assign n809 = n704 & n744 ;
  assign n810 = n322 | n809 ;
  assign n811 = ( x77 & ~n746 ) | ( x77 & n807 ) | ( ~n746 & n807 ) ;
  assign n812 = ( x78 & n810 ) | ( x78 & ~n811 ) | ( n810 & ~n811 ) ;
  assign n813 = ( x78 & n809 ) | ( x78 & n811 ) | ( n809 & n811 ) ;
  assign n814 = ( n773 & n812 ) | ( n773 & ~n813 ) | ( n812 & ~n813 ) ;
  assign n815 = n811 | n814 ;
  assign n816 = n667 & n810 ;
  assign n817 = ( ~n810 & n815 ) | ( ~n810 & n816 ) | ( n815 & n816 ) ;
  assign n818 = n817 ^ n746 ^ 1'b0 ;
  assign n819 = ( n746 & n808 ) | ( n746 & ~n818 ) | ( n808 & ~n818 ) ;
  assign n820 = n806 ^ n749 ^ x76 ;
  assign n821 = n817 ^ n749 ^ 1'b0 ;
  assign n822 = ( n749 & n820 ) | ( n749 & ~n821 ) | ( n820 & ~n821 ) ;
  assign n823 = n805 ^ n752 ^ x75 ;
  assign n824 = n817 ^ n752 ^ 1'b0 ;
  assign n825 = ( n752 & n823 ) | ( n752 & ~n824 ) | ( n823 & ~n824 ) ;
  assign n826 = n799 ^ n755 ^ x74 ;
  assign n827 = n817 ^ n755 ^ 1'b0 ;
  assign n828 = ( n755 & n826 ) | ( n755 & ~n827 ) | ( n826 & ~n827 ) ;
  assign n829 = n817 ^ n758 ^ 1'b0 ;
  assign n830 = ( n758 & n803 ) | ( n758 & ~n829 ) | ( n803 & ~n829 ) ;
  assign n831 = n817 ^ n761 ^ 1'b0 ;
  assign n832 = ( n761 & n801 ) | ( n761 & ~n831 ) | ( n801 & ~n831 ) ;
  assign n833 = n817 ^ n764 ^ 1'b0 ;
  assign n834 = ( n764 & n802 ) | ( n764 & ~n833 ) | ( n802 & ~n833 ) ;
  assign n835 = n817 ^ n795 ^ 1'b0 ;
  assign n836 = ( n795 & n804 ) | ( n795 & ~n835 ) | ( n804 & ~n835 ) ;
  assign n837 = n817 ^ n791 ^ 1'b0 ;
  assign n838 = ( n791 & n793 ) | ( n791 & ~n837 ) | ( n793 & ~n837 ) ;
  assign n839 = n817 ^ n787 ^ 1'b0 ;
  assign n840 = ( n787 & n800 ) | ( n787 & ~n839 ) | ( n800 & ~n839 ) ;
  assign n841 = n817 ^ n777 ^ 1'b0 ;
  assign n842 = ( n777 & n789 ) | ( n777 & ~n841 ) | ( n789 & ~n841 ) ;
  assign n843 = n817 ^ n783 ^ 1'b0 ;
  assign n844 = ( n767 & n783 ) | ( n767 & n843 ) | ( n783 & n843 ) ;
  assign n845 = n817 ^ n781 ^ 1'b0 ;
  assign n846 = ( n780 & n781 ) | ( n780 & n845 ) | ( n781 & n845 ) ;
  assign n847 = ( n322 & n704 ) | ( n322 & n815 ) | ( n704 & n815 ) ;
  assign n848 = n322 | n667 ;
  assign n849 = ( n322 & n847 ) | ( n322 & n848 ) | ( n847 & n848 ) ;
  assign n850 = x64 & n817 ;
  assign n851 = ~x48 & x64 ;
  assign n852 = n850 ^ x64 ^ x49 ;
  assign n853 = n852 ^ n851 ^ x65 ;
  assign n854 = ( x65 & n851 ) | ( x65 & n853 ) | ( n851 & n853 ) ;
  assign n855 = n854 ^ n846 ^ x66 ;
  assign n856 = ( x66 & n854 ) | ( x66 & n855 ) | ( n854 & n855 ) ;
  assign n857 = ( x67 & ~n844 ) | ( x67 & n856 ) | ( ~n844 & n856 ) ;
  assign n858 = ( x68 & ~n842 ) | ( x68 & n857 ) | ( ~n842 & n857 ) ;
  assign n859 = ( x69 & ~n840 ) | ( x69 & n858 ) | ( ~n840 & n858 ) ;
  assign n860 = ( x70 & ~n838 ) | ( x70 & n859 ) | ( ~n838 & n859 ) ;
  assign n861 = ( x71 & ~n836 ) | ( x71 & n860 ) | ( ~n836 & n860 ) ;
  assign n862 = ( x72 & ~n834 ) | ( x72 & n861 ) | ( ~n834 & n861 ) ;
  assign n863 = n860 ^ n836 ^ x71 ;
  assign n864 = ~n223 & n851 ;
  assign n865 = ( x73 & ~n832 ) | ( x73 & n862 ) | ( ~n832 & n862 ) ;
  assign n866 = ( x74 & ~n830 ) | ( x74 & n865 ) | ( ~n830 & n865 ) ;
  assign n867 = ( x75 & ~n828 ) | ( x75 & n866 ) | ( ~n828 & n866 ) ;
  assign n868 = ( x76 & ~n825 ) | ( x76 & n867 ) | ( ~n825 & n867 ) ;
  assign n869 = ( x77 & ~n822 ) | ( x77 & n868 ) | ( ~n822 & n868 ) ;
  assign n870 = ( x78 & ~n819 ) | ( x78 & n869 ) | ( ~n819 & n869 ) ;
  assign n871 = ( x79 & ~n849 ) | ( x79 & n870 ) | ( ~n849 & n870 ) ;
  assign n872 = n277 | n871 ;
  assign n873 = n859 ^ n838 ^ x70 ;
  assign n874 = n856 ^ n844 ^ x67 ;
  assign n875 = n872 ^ n838 ^ 1'b0 ;
  assign n876 = ( n838 & n873 ) | ( n838 & ~n875 ) | ( n873 & ~n875 ) ;
  assign n877 = n872 ^ n834 ^ 1'b0 ;
  assign n878 = n858 ^ n840 ^ x69 ;
  assign n879 = n872 ^ n822 ^ 1'b0 ;
  assign n880 = n861 ^ n834 ^ x72 ;
  assign n881 = ( n834 & ~n877 ) | ( n834 & n880 ) | ( ~n877 & n880 ) ;
  assign n882 = n872 ^ n853 ^ 1'b0 ;
  assign n883 = n869 ^ n819 ^ x78 ;
  assign n884 = n872 ^ n840 ^ 1'b0 ;
  assign n885 = ( n840 & n878 ) | ( n840 & ~n884 ) | ( n878 & ~n884 ) ;
  assign n886 = n857 ^ n842 ^ x68 ;
  assign n887 = n872 ^ n828 ^ 1'b0 ;
  assign n888 = n872 ^ n830 ^ 1'b0 ;
  assign n889 = ( n852 & n853 ) | ( n852 & n882 ) | ( n853 & n882 ) ;
  assign n890 = n872 ^ n832 ^ 1'b0 ;
  assign n891 = n872 ^ n842 ^ 1'b0 ;
  assign n892 = ( n842 & n886 ) | ( n842 & ~n891 ) | ( n886 & ~n891 ) ;
  assign n893 = n867 ^ n825 ^ x76 ;
  assign n894 = n883 ^ n872 ^ 1'b0 ;
  assign n895 = n866 ^ n828 ^ x75 ;
  assign n896 = n862 ^ n832 ^ x73 ;
  assign n897 = ( n832 & ~n890 ) | ( n832 & n896 ) | ( ~n890 & n896 ) ;
  assign n898 = n872 ^ n855 ^ 1'b0 ;
  assign n899 = n865 ^ n830 ^ x74 ;
  assign n900 = n872 ^ n836 ^ 1'b0 ;
  assign n901 = n872 ^ n844 ^ 1'b0 ;
  assign n902 = ( n844 & n874 ) | ( n844 & ~n901 ) | ( n874 & ~n901 ) ;
  assign n903 = ( n828 & ~n887 ) | ( n828 & n895 ) | ( ~n887 & n895 ) ;
  assign n904 = n868 ^ n822 ^ x77 ;
  assign n905 = ( n822 & ~n879 ) | ( n822 & n904 ) | ( ~n879 & n904 ) ;
  assign n906 = ( n846 & n855 ) | ( n846 & n898 ) | ( n855 & n898 ) ;
  assign n907 = ( n830 & ~n888 ) | ( n830 & n899 ) | ( ~n888 & n899 ) ;
  assign n908 = ( n836 & n863 ) | ( n836 & ~n900 ) | ( n863 & ~n900 ) ;
  assign n909 = ( n819 & n883 ) | ( n819 & n894 ) | ( n883 & n894 ) ;
  assign n910 = n872 ^ n825 ^ 1'b0 ;
  assign n911 = ( n825 & n893 ) | ( n825 & ~n910 ) | ( n893 & ~n910 ) ;
  assign n912 = ( ~n254 & n864 ) | ( ~n254 & n871 ) | ( n864 & n871 ) ;
  assign n913 = ~n871 & n912 ;
  assign n914 = ( ~x48 & x64 ) | ( ~x48 & n871 ) | ( x64 & n871 ) ;
  assign n915 = x64 & ~n914 ;
  assign n916 = ( ~x80 & n471 ) | ( ~x80 & n915 ) | ( n471 & n915 ) ;
  assign n917 = ~x47 & x64 ;
  assign n918 = ( n322 & n849 ) | ( n322 & n872 ) | ( n849 & n872 ) ;
  assign n919 = ~n471 & n916 ;
  assign n920 = ( x48 & n913 ) | ( x48 & ~n919 ) | ( n913 & ~n919 ) ;
  assign n921 = n920 ^ n917 ^ x65 ;
  assign n922 = ( x65 & n917 ) | ( x65 & n921 ) | ( n917 & n921 ) ;
  assign n923 = n922 ^ n889 ^ x66 ;
  assign n924 = ( x66 & n922 ) | ( x66 & n923 ) | ( n922 & n923 ) ;
  assign n925 = ( x67 & ~n906 ) | ( x67 & n924 ) | ( ~n906 & n924 ) ;
  assign n926 = ( x68 & ~n902 ) | ( x68 & n925 ) | ( ~n902 & n925 ) ;
  assign n927 = ( x69 & ~n892 ) | ( x69 & n926 ) | ( ~n892 & n926 ) ;
  assign n928 = ( x70 & ~n885 ) | ( x70 & n927 ) | ( ~n885 & n927 ) ;
  assign n929 = ( x71 & ~n876 ) | ( x71 & n928 ) | ( ~n876 & n928 ) ;
  assign n930 = ( x72 & ~n908 ) | ( x72 & n929 ) | ( ~n908 & n929 ) ;
  assign n931 = ( x73 & ~n881 ) | ( x73 & n930 ) | ( ~n881 & n930 ) ;
  assign n932 = ( x74 & ~n897 ) | ( x74 & n931 ) | ( ~n897 & n931 ) ;
  assign n933 = ( x75 & ~n907 ) | ( x75 & n932 ) | ( ~n907 & n932 ) ;
  assign n934 = ( x76 & ~n903 ) | ( x76 & n933 ) | ( ~n903 & n933 ) ;
  assign n935 = ( x77 & ~n911 ) | ( x77 & n934 ) | ( ~n911 & n934 ) ;
  assign n936 = ( x78 & ~n905 ) | ( x78 & n935 ) | ( ~n905 & n935 ) ;
  assign n937 = ( x79 & ~n909 ) | ( x79 & n936 ) | ( ~n909 & n936 ) ;
  assign n938 = n933 ^ n903 ^ x76 ;
  assign n939 = n932 ^ n907 ^ x75 ;
  assign n940 = n934 ^ n911 ^ x77 ;
  assign n941 = ( x80 & ~n918 ) | ( x80 & n937 ) | ( ~n918 & n937 ) ;
  assign n942 = n286 | n941 ;
  assign n943 = n917 & ~n941 ;
  assign n944 = ~n471 & n943 ;
  assign n945 = n942 ^ n923 ^ 1'b0 ;
  assign n946 = n931 ^ n897 ^ x74 ;
  assign n947 = ( n889 & n923 ) | ( n889 & n945 ) | ( n923 & n945 ) ;
  assign n948 = n942 ^ n911 ^ 1'b0 ;
  assign n949 = n942 ^ n921 ^ 1'b0 ;
  assign n950 = n935 ^ n905 ^ x78 ;
  assign n951 = ( n920 & n921 ) | ( n920 & n949 ) | ( n921 & n949 ) ;
  assign n952 = n942 ^ n909 ^ 1'b0 ;
  assign n953 = n936 ^ n909 ^ x79 ;
  assign n954 = n942 ^ n897 ^ 1'b0 ;
  assign n955 = ( n909 & ~n952 ) | ( n909 & n953 ) | ( ~n952 & n953 ) ;
  assign n956 = n942 ^ n903 ^ 1'b0 ;
  assign n957 = n942 ^ n907 ^ 1'b0 ;
  assign n958 = ( n903 & n938 ) | ( n903 & ~n956 ) | ( n938 & ~n956 ) ;
  assign n959 = n942 ^ n905 ^ 1'b0 ;
  assign n960 = ( n897 & n946 ) | ( n897 & ~n954 ) | ( n946 & ~n954 ) ;
  assign n961 = ( n911 & n940 ) | ( n911 & ~n948 ) | ( n940 & ~n948 ) ;
  assign n962 = ( n907 & n939 ) | ( n907 & ~n957 ) | ( n939 & ~n957 ) ;
  assign n963 = ( n905 & n950 ) | ( n905 & ~n959 ) | ( n950 & ~n959 ) ;
  assign n964 = n928 ^ n876 ^ x71 ;
  assign n965 = n924 ^ n906 ^ x67 ;
  assign n966 = n930 ^ n881 ^ x73 ;
  assign n967 = n927 ^ n885 ^ x70 ;
  assign n968 = n926 ^ n892 ^ x69 ;
  assign n969 = n929 ^ n908 ^ x72 ;
  assign n970 = x81 | n941 ;
  assign n971 = n942 ^ n885 ^ 1'b0 ;
  assign n972 = ( n885 & n967 ) | ( n885 & ~n971 ) | ( n967 & ~n971 ) ;
  assign n973 = ( n286 & n322 ) | ( n286 & n918 ) | ( n322 & n918 ) ;
  assign n974 = n942 ^ n908 ^ 1'b0 ;
  assign n975 = n918 & n942 ;
  assign n976 = ( n908 & n969 ) | ( n908 & ~n974 ) | ( n969 & ~n974 ) ;
  assign n977 = ~x46 & x64 ;
  assign n978 = n942 ^ n876 ^ 1'b0 ;
  assign n979 = ( n876 & n964 ) | ( n876 & ~n978 ) | ( n964 & ~n978 ) ;
  assign n980 = n942 ^ n881 ^ 1'b0 ;
  assign n981 = x81 & n975 ;
  assign n982 = ( n881 & n966 ) | ( n881 & ~n980 ) | ( n966 & ~n980 ) ;
  assign n983 = n942 ^ n892 ^ 1'b0 ;
  assign n984 = n225 | n243 ;
  assign n985 = ( n892 & n968 ) | ( n892 & ~n983 ) | ( n968 & ~n983 ) ;
  assign n986 = x82 | x83 ;
  assign n987 = ( ~n166 & n984 ) | ( ~n166 & n986 ) | ( n984 & n986 ) ;
  assign n988 = n322 | n975 ;
  assign n989 = n942 ^ n906 ^ 1'b0 ;
  assign n990 = ( n906 & n965 ) | ( n906 & ~n989 ) | ( n965 & ~n989 ) ;
  assign n991 = n942 ^ n902 ^ 1'b0 ;
  assign n992 = n925 ^ n902 ^ x68 ;
  assign n993 = ( n902 & ~n991 ) | ( n902 & n992 ) | ( ~n991 & n992 ) ;
  assign n994 = n166 | n987 ;
  assign n995 = x47 & x64 ;
  assign n996 = n286 & n988 ;
  assign n997 = ~n994 & n995 ;
  assign n998 = ~n970 & n997 ;
  assign n999 = ( x47 & n944 ) | ( x47 & ~n998 ) | ( n944 & ~n998 ) ;
  assign n1000 = x81 | n988 ;
  assign n1001 = n999 ^ n977 ^ x65 ;
  assign n1002 = ( x65 & n977 ) | ( x65 & n1001 ) | ( n977 & n1001 ) ;
  assign n1003 = n1002 ^ n951 ^ x66 ;
  assign n1004 = ( ~n981 & n994 ) | ( ~n981 & n1000 ) | ( n994 & n1000 ) ;
  assign n1005 = ( x66 & n1002 ) | ( x66 & n1003 ) | ( n1002 & n1003 ) ;
  assign n1006 = ( x67 & ~n947 ) | ( x67 & n1005 ) | ( ~n947 & n1005 ) ;
  assign n1007 = ( x68 & ~n990 ) | ( x68 & n1006 ) | ( ~n990 & n1006 ) ;
  assign n1008 = ( x69 & ~n993 ) | ( x69 & n1007 ) | ( ~n993 & n1007 ) ;
  assign n1009 = ( x70 & ~n985 ) | ( x70 & n1008 ) | ( ~n985 & n1008 ) ;
  assign n1010 = ( x71 & ~n972 ) | ( x71 & n1009 ) | ( ~n972 & n1009 ) ;
  assign n1011 = ( x72 & ~n979 ) | ( x72 & n1010 ) | ( ~n979 & n1010 ) ;
  assign n1012 = ( x73 & ~n976 ) | ( x73 & n1011 ) | ( ~n976 & n1011 ) ;
  assign n1013 = ( x74 & ~n982 ) | ( x74 & n1012 ) | ( ~n982 & n1012 ) ;
  assign n1014 = ( x75 & ~n960 ) | ( x75 & n1013 ) | ( ~n960 & n1013 ) ;
  assign n1015 = ( x76 & ~n962 ) | ( x76 & n1014 ) | ( ~n962 & n1014 ) ;
  assign n1016 = ( x77 & ~n958 ) | ( x77 & n1015 ) | ( ~n958 & n1015 ) ;
  assign n1017 = ( x78 & ~n961 ) | ( x78 & n1016 ) | ( ~n961 & n1016 ) ;
  assign n1018 = ( x79 & ~n963 ) | ( x79 & n1017 ) | ( ~n963 & n1017 ) ;
  assign n1019 = ( x80 & ~n955 ) | ( x80 & n1018 ) | ( ~n955 & n1018 ) ;
  assign n1020 = n1004 | n1019 ;
  assign n1021 = ( ~n988 & n996 ) | ( ~n988 & n1020 ) | ( n996 & n1020 ) ;
  assign n1022 = n1017 ^ n963 ^ x79 ;
  assign n1023 = n1021 ^ n963 ^ 1'b0 ;
  assign n1024 = ( n963 & n1022 ) | ( n963 & ~n1023 ) | ( n1022 & ~n1023 ) ;
  assign n1025 = n1016 ^ n961 ^ x78 ;
  assign n1026 = n1021 ^ n961 ^ 1'b0 ;
  assign n1027 = ( n961 & n1025 ) | ( n961 & ~n1026 ) | ( n1025 & ~n1026 ) ;
  assign n1028 = n1015 ^ n958 ^ x77 ;
  assign n1029 = n1021 ^ n958 ^ 1'b0 ;
  assign n1030 = ( n958 & n1028 ) | ( n958 & ~n1029 ) | ( n1028 & ~n1029 ) ;
  assign n1031 = n1014 ^ n962 ^ x76 ;
  assign n1032 = n1021 ^ n962 ^ 1'b0 ;
  assign n1033 = ( n962 & n1031 ) | ( n962 & ~n1032 ) | ( n1031 & ~n1032 ) ;
  assign n1034 = n1013 ^ n960 ^ x75 ;
  assign n1035 = n1021 ^ n960 ^ 1'b0 ;
  assign n1036 = ( n960 & n1034 ) | ( n960 & ~n1035 ) | ( n1034 & ~n1035 ) ;
  assign n1037 = n1012 ^ n982 ^ x74 ;
  assign n1038 = n1021 ^ n982 ^ 1'b0 ;
  assign n1039 = ( n982 & n1037 ) | ( n982 & ~n1038 ) | ( n1037 & ~n1038 ) ;
  assign n1040 = n1011 ^ n976 ^ x73 ;
  assign n1041 = n1021 ^ n976 ^ 1'b0 ;
  assign n1042 = ( n976 & n1040 ) | ( n976 & ~n1041 ) | ( n1040 & ~n1041 ) ;
  assign n1043 = n1010 ^ n979 ^ x72 ;
  assign n1044 = n1021 ^ n979 ^ 1'b0 ;
  assign n1045 = ( n979 & n1043 ) | ( n979 & ~n1044 ) | ( n1043 & ~n1044 ) ;
  assign n1046 = n1009 ^ n972 ^ x71 ;
  assign n1047 = n1021 ^ n972 ^ 1'b0 ;
  assign n1048 = ( n972 & n1046 ) | ( n972 & ~n1047 ) | ( n1046 & ~n1047 ) ;
  assign n1049 = n1008 ^ n985 ^ x70 ;
  assign n1050 = n1021 ^ n985 ^ 1'b0 ;
  assign n1051 = ( n985 & n1049 ) | ( n985 & ~n1050 ) | ( n1049 & ~n1050 ) ;
  assign n1052 = n1021 ^ n1003 ^ 1'b0 ;
  assign n1053 = ( n951 & n1003 ) | ( n951 & n1052 ) | ( n1003 & n1052 ) ;
  assign n1054 = n1021 ^ n1001 ^ 1'b0 ;
  assign n1055 = ( n999 & n1001 ) | ( n999 & n1054 ) | ( n1001 & n1054 ) ;
  assign n1056 = n322 | n1020 ;
  assign n1057 = ( n322 & n973 ) | ( n322 & n1056 ) | ( n973 & n1056 ) ;
  assign n1058 = n1018 ^ n955 ^ x80 ;
  assign n1059 = n1021 ^ n955 ^ 1'b0 ;
  assign n1060 = ( n955 & n1058 ) | ( n955 & ~n1059 ) | ( n1058 & ~n1059 ) ;
  assign n1061 = n1007 ^ n993 ^ x69 ;
  assign n1062 = n1021 ^ n993 ^ 1'b0 ;
  assign n1063 = ( n993 & n1061 ) | ( n993 & ~n1062 ) | ( n1061 & ~n1062 ) ;
  assign n1064 = n1006 ^ n990 ^ x68 ;
  assign n1065 = n1021 ^ n990 ^ 1'b0 ;
  assign n1066 = ( n990 & n1064 ) | ( n990 & ~n1065 ) | ( n1064 & ~n1065 ) ;
  assign n1067 = n1005 ^ n947 ^ x67 ;
  assign n1068 = n1021 ^ n947 ^ 1'b0 ;
  assign n1069 = ( n947 & n1067 ) | ( n947 & ~n1068 ) | ( n1067 & ~n1068 ) ;
  assign n1070 = ~x45 & x64 ;
  assign n1071 = x64 & n1021 ;
  assign n1072 = n1071 ^ x64 ^ x46 ;
  assign n1073 = n1072 ^ n1070 ^ x65 ;
  assign n1074 = ( x65 & n1070 ) | ( x65 & n1073 ) | ( n1070 & n1073 ) ;
  assign n1075 = n1074 ^ n1055 ^ x66 ;
  assign n1076 = ( x66 & n1074 ) | ( x66 & n1075 ) | ( n1074 & n1075 ) ;
  assign n1077 = ( x67 & ~n1053 ) | ( x67 & n1076 ) | ( ~n1053 & n1076 ) ;
  assign n1078 = ( x68 & ~n1069 ) | ( x68 & n1077 ) | ( ~n1069 & n1077 ) ;
  assign n1079 = ( x69 & ~n1066 ) | ( x69 & n1078 ) | ( ~n1066 & n1078 ) ;
  assign n1080 = ( x70 & ~n1063 ) | ( x70 & n1079 ) | ( ~n1063 & n1079 ) ;
  assign n1081 = ( x71 & ~n1051 ) | ( x71 & n1080 ) | ( ~n1051 & n1080 ) ;
  assign n1082 = ( x72 & ~n1048 ) | ( x72 & n1081 ) | ( ~n1048 & n1081 ) ;
  assign n1083 = ( x73 & ~n1045 ) | ( x73 & n1082 ) | ( ~n1045 & n1082 ) ;
  assign n1084 = ( x74 & ~n1042 ) | ( x74 & n1083 ) | ( ~n1042 & n1083 ) ;
  assign n1085 = ( x75 & ~n1039 ) | ( x75 & n1084 ) | ( ~n1039 & n1084 ) ;
  assign n1086 = ( x76 & ~n1036 ) | ( x76 & n1085 ) | ( ~n1036 & n1085 ) ;
  assign n1087 = ( x77 & ~n1033 ) | ( x77 & n1086 ) | ( ~n1033 & n1086 ) ;
  assign n1088 = ( x78 & ~n1030 ) | ( x78 & n1087 ) | ( ~n1030 & n1087 ) ;
  assign n1089 = ( x79 & ~n1027 ) | ( x79 & n1088 ) | ( ~n1027 & n1088 ) ;
  assign n1090 = ( x80 & ~n1024 ) | ( x80 & n1089 ) | ( ~n1024 & n1089 ) ;
  assign n1091 = n202 | n262 ;
  assign n1092 = ( x81 & ~n1060 ) | ( x81 & n1090 ) | ( ~n1060 & n1090 ) ;
  assign n1093 = ( x82 & ~n1057 ) | ( x82 & n1092 ) | ( ~n1057 & n1092 ) ;
  assign n1094 = ( ~n195 & n1091 ) | ( ~n195 & n1093 ) | ( n1091 & n1093 ) ;
  assign n1095 = n195 | n1094 ;
  assign n1096 = n1086 ^ n1033 ^ x77 ;
  assign n1097 = n1095 ^ n1033 ^ 1'b0 ;
  assign n1098 = ( n1033 & n1096 ) | ( n1033 & ~n1097 ) | ( n1096 & ~n1097 ) ;
  assign n1099 = n1084 ^ n1039 ^ x75 ;
  assign n1100 = n1095 ^ n1039 ^ 1'b0 ;
  assign n1101 = ( n1039 & n1099 ) | ( n1039 & ~n1100 ) | ( n1099 & ~n1100 ) ;
  assign n1102 = n1080 ^ n1051 ^ x71 ;
  assign n1103 = n1095 ^ n1051 ^ 1'b0 ;
  assign n1104 = ( n1051 & n1102 ) | ( n1051 & ~n1103 ) | ( n1102 & ~n1103 ) ;
  assign n1105 = n1076 ^ n1053 ^ x67 ;
  assign n1106 = n1095 ^ n1053 ^ 1'b0 ;
  assign n1107 = ( n1053 & n1105 ) | ( n1053 & ~n1106 ) | ( n1105 & ~n1106 ) ;
  assign n1108 = n1095 ^ n1073 ^ 1'b0 ;
  assign n1109 = ( n1072 & n1073 ) | ( n1072 & n1108 ) | ( n1073 & n1108 ) ;
  assign n1110 = n1090 ^ n1060 ^ x81 ;
  assign n1111 = n1110 ^ n1095 ^ 1'b0 ;
  assign n1112 = ( n1060 & n1110 ) | ( n1060 & n1111 ) | ( n1110 & n1111 ) ;
  assign n1113 = n1089 ^ n1024 ^ x80 ;
  assign n1114 = n1095 ^ n1024 ^ 1'b0 ;
  assign n1115 = ( n1024 & n1113 ) | ( n1024 & ~n1114 ) | ( n1113 & ~n1114 ) ;
  assign n1116 = n1088 ^ n1027 ^ x79 ;
  assign n1117 = n1095 ^ n1027 ^ 1'b0 ;
  assign n1118 = ( n1027 & n1116 ) | ( n1027 & ~n1117 ) | ( n1116 & ~n1117 ) ;
  assign n1119 = n1087 ^ n1030 ^ x78 ;
  assign n1120 = n1095 ^ n1030 ^ 1'b0 ;
  assign n1121 = ( n1030 & n1119 ) | ( n1030 & ~n1120 ) | ( n1119 & ~n1120 ) ;
  assign n1122 = n1085 ^ n1036 ^ x76 ;
  assign n1123 = n1095 ^ n1036 ^ 1'b0 ;
  assign n1124 = ( n1036 & n1122 ) | ( n1036 & ~n1123 ) | ( n1122 & ~n1123 ) ;
  assign n1125 = n1083 ^ n1042 ^ x74 ;
  assign n1126 = n1095 ^ n1042 ^ 1'b0 ;
  assign n1127 = ( n1042 & n1125 ) | ( n1042 & ~n1126 ) | ( n1125 & ~n1126 ) ;
  assign n1128 = n1082 ^ n1045 ^ x73 ;
  assign n1129 = n1095 ^ n1045 ^ 1'b0 ;
  assign n1130 = ( n1045 & n1128 ) | ( n1045 & ~n1129 ) | ( n1128 & ~n1129 ) ;
  assign n1131 = n1081 ^ n1048 ^ x72 ;
  assign n1132 = n1095 ^ n1048 ^ 1'b0 ;
  assign n1133 = ( n1048 & n1131 ) | ( n1048 & ~n1132 ) | ( n1131 & ~n1132 ) ;
  assign n1134 = n1079 ^ n1063 ^ x70 ;
  assign n1135 = n1095 ^ n1063 ^ 1'b0 ;
  assign n1136 = ( n1063 & n1134 ) | ( n1063 & ~n1135 ) | ( n1134 & ~n1135 ) ;
  assign n1137 = n1078 ^ n1066 ^ x69 ;
  assign n1138 = n1095 ^ n1066 ^ 1'b0 ;
  assign n1139 = ( n1066 & n1137 ) | ( n1066 & ~n1138 ) | ( n1137 & ~n1138 ) ;
  assign n1140 = n1077 ^ n1069 ^ x68 ;
  assign n1141 = n1095 ^ n1069 ^ 1'b0 ;
  assign n1142 = ( n1069 & n1140 ) | ( n1069 & ~n1141 ) | ( n1140 & ~n1141 ) ;
  assign n1143 = n1095 ^ n1075 ^ 1'b0 ;
  assign n1144 = ( n1055 & n1075 ) | ( n1055 & n1143 ) | ( n1075 & n1143 ) ;
  assign n1145 = n1070 & ~n1095 ;
  assign n1146 = x64 & ~x83 ;
  assign n1147 = ( ~n166 & n225 ) | ( ~n166 & n1146 ) | ( n225 & n1146 ) ;
  assign n1148 = ~n984 & n1147 ;
  assign n1149 = ( x45 & n1093 ) | ( x45 & ~n1148 ) | ( n1093 & ~n1148 ) ;
  assign n1150 = x45 & ~n1149 ;
  assign n1151 = ( x45 & n1145 ) | ( x45 & ~n1150 ) | ( n1145 & ~n1150 ) ;
  assign n1152 = ( n322 & n1057 ) | ( n322 & n1095 ) | ( n1057 & n1095 ) ;
  assign n1153 = ~x44 & x64 ;
  assign n1154 = n1153 ^ n1151 ^ x65 ;
  assign n1155 = ( x65 & n1153 ) | ( x65 & n1154 ) | ( n1153 & n1154 ) ;
  assign n1156 = n1155 ^ n1109 ^ x66 ;
  assign n1157 = ( x66 & n1155 ) | ( x66 & n1156 ) | ( n1155 & n1156 ) ;
  assign n1158 = ( x67 & ~n1144 ) | ( x67 & n1157 ) | ( ~n1144 & n1157 ) ;
  assign n1159 = ( x68 & ~n1107 ) | ( x68 & n1158 ) | ( ~n1107 & n1158 ) ;
  assign n1160 = ( x69 & ~n1142 ) | ( x69 & n1159 ) | ( ~n1142 & n1159 ) ;
  assign n1161 = ( x70 & ~n1139 ) | ( x70 & n1160 ) | ( ~n1139 & n1160 ) ;
  assign n1162 = ( x71 & ~n1136 ) | ( x71 & n1161 ) | ( ~n1136 & n1161 ) ;
  assign n1163 = ( x72 & ~n1104 ) | ( x72 & n1162 ) | ( ~n1104 & n1162 ) ;
  assign n1164 = ( x73 & ~n1133 ) | ( x73 & n1163 ) | ( ~n1133 & n1163 ) ;
  assign n1165 = ( x74 & ~n1130 ) | ( x74 & n1164 ) | ( ~n1130 & n1164 ) ;
  assign n1166 = ( x75 & ~n1127 ) | ( x75 & n1165 ) | ( ~n1127 & n1165 ) ;
  assign n1167 = ( x76 & ~n1101 ) | ( x76 & n1166 ) | ( ~n1101 & n1166 ) ;
  assign n1168 = ( x77 & ~n1124 ) | ( x77 & n1167 ) | ( ~n1124 & n1167 ) ;
  assign n1169 = ( x78 & ~n1098 ) | ( x78 & n1168 ) | ( ~n1098 & n1168 ) ;
  assign n1170 = ( x79 & ~n1121 ) | ( x79 & n1169 ) | ( ~n1121 & n1169 ) ;
  assign n1171 = ( x80 & ~n1118 ) | ( x80 & n1170 ) | ( ~n1118 & n1170 ) ;
  assign n1172 = ( x81 & ~n1115 ) | ( x81 & n1171 ) | ( ~n1115 & n1171 ) ;
  assign n1173 = ( x82 & ~n1112 ) | ( x82 & n1172 ) | ( ~n1112 & n1172 ) ;
  assign n1174 = ( x83 & ~n1152 ) | ( x83 & n1173 ) | ( ~n1152 & n1173 ) ;
  assign n1175 = n254 | n1174 ;
  assign n1176 = ~n166 & n1153 ;
  assign n1177 = n1175 ^ n1118 ^ 1'b0 ;
  assign n1178 = n1171 ^ n1115 ^ x81 ;
  assign n1179 = n1169 ^ n1121 ^ x79 ;
  assign n1180 = n1170 ^ n1118 ^ x80 ;
  assign n1181 = ( n1118 & ~n1177 ) | ( n1118 & n1180 ) | ( ~n1177 & n1180 ) ;
  assign n1182 = n1175 ^ n1156 ^ 1'b0 ;
  assign n1183 = n1175 ^ n1124 ^ 1'b0 ;
  assign n1184 = ( n1109 & n1156 ) | ( n1109 & n1182 ) | ( n1156 & n1182 ) ;
  assign n1185 = n1175 ^ n1154 ^ 1'b0 ;
  assign n1186 = n1175 ^ n1144 ^ 1'b0 ;
  assign n1187 = n1157 ^ n1144 ^ x67 ;
  assign n1188 = n1167 ^ n1124 ^ x77 ;
  assign n1189 = n1165 ^ n1127 ^ x75 ;
  assign n1190 = ( n1124 & ~n1183 ) | ( n1124 & n1188 ) | ( ~n1183 & n1188 ) ;
  assign n1191 = n1175 ^ n1127 ^ 1'b0 ;
  assign n1192 = n1175 ^ n1121 ^ 1'b0 ;
  assign n1193 = ( n1151 & n1154 ) | ( n1151 & n1185 ) | ( n1154 & n1185 ) ;
  assign n1194 = ( n1121 & n1179 ) | ( n1121 & ~n1192 ) | ( n1179 & ~n1192 ) ;
  assign n1195 = ( n1144 & ~n1186 ) | ( n1144 & n1187 ) | ( ~n1186 & n1187 ) ;
  assign n1196 = n1175 ^ n1115 ^ 1'b0 ;
  assign n1197 = ( n1127 & n1189 ) | ( n1127 & ~n1191 ) | ( n1189 & ~n1191 ) ;
  assign n1198 = ( n1115 & n1178 ) | ( n1115 & ~n1196 ) | ( n1178 & ~n1196 ) ;
  assign n1199 = n1172 ^ n1112 ^ x82 ;
  assign n1200 = n1175 ^ n1112 ^ 1'b0 ;
  assign n1201 = ( n1112 & n1199 ) | ( n1112 & ~n1200 ) | ( n1199 & ~n1200 ) ;
  assign n1202 = n1168 ^ n1098 ^ x78 ;
  assign n1203 = n1175 ^ n1098 ^ 1'b0 ;
  assign n1204 = ( n1098 & n1202 ) | ( n1098 & ~n1203 ) | ( n1202 & ~n1203 ) ;
  assign n1205 = n1175 ^ n1101 ^ 1'b0 ;
  assign n1206 = n1164 ^ n1130 ^ x74 ;
  assign n1207 = n1175 ^ n1130 ^ 1'b0 ;
  assign n1208 = ( n1130 & n1206 ) | ( n1130 & ~n1207 ) | ( n1206 & ~n1207 ) ;
  assign n1209 = n1163 ^ n1133 ^ x73 ;
  assign n1210 = n1175 ^ n1133 ^ 1'b0 ;
  assign n1211 = n1166 ^ n1101 ^ x76 ;
  assign n1212 = ( n1101 & ~n1205 ) | ( n1101 & n1211 ) | ( ~n1205 & n1211 ) ;
  assign n1213 = ( n1133 & n1209 ) | ( n1133 & ~n1210 ) | ( n1209 & ~n1210 ) ;
  assign n1214 = n1162 ^ n1104 ^ x72 ;
  assign n1215 = n1175 ^ n1104 ^ 1'b0 ;
  assign n1216 = ( n1104 & n1214 ) | ( n1104 & ~n1215 ) | ( n1214 & ~n1215 ) ;
  assign n1217 = n1161 ^ n1136 ^ x71 ;
  assign n1218 = n1175 ^ n1136 ^ 1'b0 ;
  assign n1219 = ( n1136 & n1217 ) | ( n1136 & ~n1218 ) | ( n1217 & ~n1218 ) ;
  assign n1220 = n1160 ^ n1139 ^ x70 ;
  assign n1221 = n1175 ^ n1139 ^ 1'b0 ;
  assign n1222 = ( n1139 & n1220 ) | ( n1139 & ~n1221 ) | ( n1220 & ~n1221 ) ;
  assign n1223 = n1159 ^ n1142 ^ x69 ;
  assign n1224 = n1175 ^ n1142 ^ 1'b0 ;
  assign n1225 = ( n1142 & n1223 ) | ( n1142 & ~n1224 ) | ( n1223 & ~n1224 ) ;
  assign n1226 = n1158 ^ n1107 ^ x68 ;
  assign n1227 = n1175 ^ n1107 ^ 1'b0 ;
  assign n1228 = ( n1107 & n1226 ) | ( n1107 & ~n1227 ) | ( n1226 & ~n1227 ) ;
  assign n1229 = ( ~n984 & n1174 ) | ( ~n984 & n1176 ) | ( n1174 & n1176 ) ;
  assign n1230 = ~n1174 & n1229 ;
  assign n1231 = x44 & x64 ;
  assign n1232 = ( ~x84 & n202 ) | ( ~x84 & n1231 ) | ( n202 & n1231 ) ;
  assign n1233 = ~n202 & n1232 ;
  assign n1234 = ( ~n195 & n1174 ) | ( ~n195 & n1233 ) | ( n1174 & n1233 ) ;
  assign n1235 = ~n1174 & n1234 ;
  assign n1236 = ( x44 & n1230 ) | ( x44 & ~n1235 ) | ( n1230 & ~n1235 ) ;
  assign n1237 = ~x43 & x64 ;
  assign n1238 = n1237 ^ n1236 ^ x65 ;
  assign n1239 = ( x65 & n1237 ) | ( x65 & n1238 ) | ( n1237 & n1238 ) ;
  assign n1240 = n1239 ^ n1193 ^ x66 ;
  assign n1241 = ( x66 & n1239 ) | ( x66 & n1240 ) | ( n1239 & n1240 ) ;
  assign n1242 = ( x67 & ~n1184 ) | ( x67 & n1241 ) | ( ~n1184 & n1241 ) ;
  assign n1243 = ( x68 & ~n1195 ) | ( x68 & n1242 ) | ( ~n1195 & n1242 ) ;
  assign n1244 = ( x69 & ~n1228 ) | ( x69 & n1243 ) | ( ~n1228 & n1243 ) ;
  assign n1245 = ( x70 & ~n1225 ) | ( x70 & n1244 ) | ( ~n1225 & n1244 ) ;
  assign n1246 = ( x71 & ~n1222 ) | ( x71 & n1245 ) | ( ~n1222 & n1245 ) ;
  assign n1247 = ( x72 & ~n1219 ) | ( x72 & n1246 ) | ( ~n1219 & n1246 ) ;
  assign n1248 = ( x73 & ~n1216 ) | ( x73 & n1247 ) | ( ~n1216 & n1247 ) ;
  assign n1249 = ( x74 & ~n1213 ) | ( x74 & n1248 ) | ( ~n1213 & n1248 ) ;
  assign n1250 = ( x75 & ~n1208 ) | ( x75 & n1249 ) | ( ~n1208 & n1249 ) ;
  assign n1251 = ( x76 & ~n1197 ) | ( x76 & n1250 ) | ( ~n1197 & n1250 ) ;
  assign n1252 = ( x77 & ~n1212 ) | ( x77 & n1251 ) | ( ~n1212 & n1251 ) ;
  assign n1253 = ( x78 & ~n1190 ) | ( x78 & n1252 ) | ( ~n1190 & n1252 ) ;
  assign n1254 = ( x79 & ~n1204 ) | ( x79 & n1253 ) | ( ~n1204 & n1253 ) ;
  assign n1255 = ( x80 & ~n1194 ) | ( x80 & n1254 ) | ( ~n1194 & n1254 ) ;
  assign n1256 = ( x81 & ~n1181 ) | ( x81 & n1255 ) | ( ~n1181 & n1255 ) ;
  assign n1257 = ( x82 & ~n1198 ) | ( x82 & n1256 ) | ( ~n1198 & n1256 ) ;
  assign n1258 = n1152 & n1175 ;
  assign n1259 = n322 | n1258 ;
  assign n1260 = ( x83 & ~n1201 ) | ( x83 & n1257 ) | ( ~n1201 & n1257 ) ;
  assign n1261 = ( x84 & n470 ) | ( x84 & ~n1258 ) | ( n470 & ~n1258 ) ;
  assign n1262 = ( ~x84 & n470 ) | ( ~x84 & n1259 ) | ( n470 & n1259 ) ;
  assign n1263 = ( ~n1260 & n1261 ) | ( ~n1260 & n1262 ) | ( n1261 & n1262 ) ;
  assign n1264 = n1260 | n1263 ;
  assign n1265 = n254 & n1259 ;
  assign n1266 = ( ~n1259 & n1264 ) | ( ~n1259 & n1265 ) | ( n1264 & n1265 ) ;
  assign n1267 = n1247 ^ n1216 ^ x73 ;
  assign n1268 = n1266 ^ n1216 ^ 1'b0 ;
  assign n1269 = ( n1216 & n1267 ) | ( n1216 & ~n1268 ) | ( n1267 & ~n1268 ) ;
  assign n1270 = n1244 ^ n1225 ^ x70 ;
  assign n1271 = n1266 ^ n1225 ^ 1'b0 ;
  assign n1272 = ( n1225 & n1270 ) | ( n1225 & ~n1271 ) | ( n1270 & ~n1271 ) ;
  assign n1273 = n1243 ^ n1228 ^ x69 ;
  assign n1274 = n1266 ^ n1228 ^ 1'b0 ;
  assign n1275 = ( n1228 & n1273 ) | ( n1228 & ~n1274 ) | ( n1273 & ~n1274 ) ;
  assign n1276 = n1241 ^ n1184 ^ x67 ;
  assign n1277 = n1266 ^ n1184 ^ 1'b0 ;
  assign n1278 = ( n1184 & n1276 ) | ( n1184 & ~n1277 ) | ( n1276 & ~n1277 ) ;
  assign n1279 = n1266 ^ n1240 ^ 1'b0 ;
  assign n1280 = ( n1193 & n1240 ) | ( n1193 & n1279 ) | ( n1240 & n1279 ) ;
  assign n1281 = n1266 ^ n1238 ^ 1'b0 ;
  assign n1282 = ( n1236 & n1238 ) | ( n1236 & n1281 ) | ( n1238 & n1281 ) ;
  assign n1283 = ( n254 & n322 ) | ( n254 & n1152 ) | ( n322 & n1152 ) ;
  assign n1284 = n322 | n1264 ;
  assign n1285 = ( n322 & n1283 ) | ( n322 & n1284 ) | ( n1283 & n1284 ) ;
  assign n1286 = n1253 ^ n1204 ^ x79 ;
  assign n1287 = n1248 ^ n1213 ^ x74 ;
  assign n1288 = n1256 ^ n1198 ^ x82 ;
  assign n1289 = n1246 ^ n1219 ^ x72 ;
  assign n1290 = n1266 ^ n1204 ^ 1'b0 ;
  assign n1291 = ( n1204 & n1286 ) | ( n1204 & ~n1290 ) | ( n1286 & ~n1290 ) ;
  assign n1292 = n1266 ^ n1197 ^ 1'b0 ;
  assign n1293 = n1266 ^ n1181 ^ 1'b0 ;
  assign n1294 = n1254 ^ n1194 ^ x80 ;
  assign n1295 = n1250 ^ n1197 ^ x76 ;
  assign n1296 = n131 | n156 ;
  assign n1297 = n151 | n164 ;
  assign n1298 = n158 | n159 ;
  assign n1299 = n1252 ^ n1190 ^ x78 ;
  assign n1300 = n1249 ^ n1208 ^ x75 ;
  assign n1301 = n1255 ^ n1181 ^ x81 ;
  assign n1302 = n199 | n247 ;
  assign n1303 = n1245 ^ n1222 ^ x71 ;
  assign n1304 = ( n1181 & ~n1293 ) | ( n1181 & n1301 ) | ( ~n1293 & n1301 ) ;
  assign n1305 = n1266 ^ n1212 ^ 1'b0 ;
  assign n1306 = n1251 ^ n1212 ^ x77 ;
  assign n1307 = n1266 ^ n1194 ^ 1'b0 ;
  assign n1308 = ( n1194 & n1294 ) | ( n1194 & ~n1307 ) | ( n1294 & ~n1307 ) ;
  assign n1309 = n1266 ^ n1198 ^ 1'b0 ;
  assign n1310 = n143 | n202 ;
  assign n1311 = n1266 ^ n1190 ^ 1'b0 ;
  assign n1312 = ( n1190 & n1299 ) | ( n1190 & ~n1311 ) | ( n1299 & ~n1311 ) ;
  assign n1313 = n1266 ^ n1195 ^ 1'b0 ;
  assign n1314 = n1266 ^ n1219 ^ 1'b0 ;
  assign n1315 = ( n1198 & n1288 ) | ( n1198 & ~n1309 ) | ( n1288 & ~n1309 ) ;
  assign n1316 = n1257 ^ n1201 ^ x83 ;
  assign n1317 = n1266 ^ n1213 ^ 1'b0 ;
  assign n1318 = n1266 ^ n1208 ^ 1'b0 ;
  assign n1319 = n1242 ^ n1195 ^ x68 ;
  assign n1320 = ( n1213 & n1287 ) | ( n1213 & ~n1317 ) | ( n1287 & ~n1317 ) ;
  assign n1321 = n1266 ^ n1222 ^ 1'b0 ;
  assign n1322 = n1266 ^ n1201 ^ 1'b0 ;
  assign n1323 = ( n1219 & n1289 ) | ( n1219 & ~n1314 ) | ( n1289 & ~n1314 ) ;
  assign n1324 = ( n1201 & n1316 ) | ( n1201 & ~n1322 ) | ( n1316 & ~n1322 ) ;
  assign n1325 = ( n1212 & ~n1305 ) | ( n1212 & n1306 ) | ( ~n1305 & n1306 ) ;
  assign n1326 = ( n1197 & ~n1292 ) | ( n1197 & n1295 ) | ( ~n1292 & n1295 ) ;
  assign n1327 = ( n1208 & n1300 ) | ( n1208 & ~n1318 ) | ( n1300 & ~n1318 ) ;
  assign n1328 = ( n1195 & ~n1313 ) | ( n1195 & n1319 ) | ( ~n1313 & n1319 ) ;
  assign n1329 = ( n1222 & n1303 ) | ( n1222 & ~n1321 ) | ( n1303 & ~n1321 ) ;
  assign n1330 = ~x42 & x64 ;
  assign n1331 = x64 & n1266 ;
  assign n1332 = n1331 ^ x64 ^ x43 ;
  assign n1333 = n1332 ^ n1330 ^ x65 ;
  assign n1334 = ( x65 & n1330 ) | ( x65 & n1333 ) | ( n1330 & n1333 ) ;
  assign n1335 = n1334 ^ n1282 ^ x66 ;
  assign n1336 = ( x66 & n1334 ) | ( x66 & n1335 ) | ( n1334 & n1335 ) ;
  assign n1337 = ( x67 & ~n1280 ) | ( x67 & n1336 ) | ( ~n1280 & n1336 ) ;
  assign n1338 = ( x68 & ~n1278 ) | ( x68 & n1337 ) | ( ~n1278 & n1337 ) ;
  assign n1339 = ( x69 & ~n1328 ) | ( x69 & n1338 ) | ( ~n1328 & n1338 ) ;
  assign n1340 = ( x70 & ~n1275 ) | ( x70 & n1339 ) | ( ~n1275 & n1339 ) ;
  assign n1341 = ( x71 & ~n1272 ) | ( x71 & n1340 ) | ( ~n1272 & n1340 ) ;
  assign n1342 = ( x72 & ~n1329 ) | ( x72 & n1341 ) | ( ~n1329 & n1341 ) ;
  assign n1343 = ( x73 & ~n1323 ) | ( x73 & n1342 ) | ( ~n1323 & n1342 ) ;
  assign n1344 = ( x74 & ~n1269 ) | ( x74 & n1343 ) | ( ~n1269 & n1343 ) ;
  assign n1345 = ( x75 & ~n1320 ) | ( x75 & n1344 ) | ( ~n1320 & n1344 ) ;
  assign n1346 = x86 | x87 ;
  assign n1347 = n1343 ^ n1269 ^ x74 ;
  assign n1348 = ( x76 & ~n1327 ) | ( x76 & n1345 ) | ( ~n1327 & n1345 ) ;
  assign n1349 = ( x77 & ~n1326 ) | ( x77 & n1348 ) | ( ~n1326 & n1348 ) ;
  assign n1350 = ( x78 & ~n1325 ) | ( x78 & n1349 ) | ( ~n1325 & n1349 ) ;
  assign n1351 = ( x79 & ~n1312 ) | ( x79 & n1350 ) | ( ~n1312 & n1350 ) ;
  assign n1352 = ( x80 & ~n1291 ) | ( x80 & n1351 ) | ( ~n1291 & n1351 ) ;
  assign n1353 = ( x81 & ~n1308 ) | ( x81 & n1352 ) | ( ~n1308 & n1352 ) ;
  assign n1354 = ( x82 & ~n1304 ) | ( x82 & n1353 ) | ( ~n1304 & n1353 ) ;
  assign n1355 = ( x83 & ~n1315 ) | ( x83 & n1354 ) | ( ~n1315 & n1354 ) ;
  assign n1356 = ( x84 & ~n1324 ) | ( x84 & n1355 ) | ( ~n1324 & n1355 ) ;
  assign n1357 = ( x85 & ~n1285 ) | ( x85 & n1356 ) | ( ~n1285 & n1356 ) ;
  assign n1358 = ( ~n1302 & n1346 ) | ( ~n1302 & n1357 ) | ( n1346 & n1357 ) ;
  assign n1359 = n1302 | n1358 ;
  assign n1360 = n1359 ^ n1269 ^ 1'b0 ;
  assign n1361 = ( n1269 & n1347 ) | ( n1269 & ~n1360 ) | ( n1347 & ~n1360 ) ;
  assign n1362 = n1341 ^ n1329 ^ x72 ;
  assign n1363 = n1359 ^ n1329 ^ 1'b0 ;
  assign n1364 = ( n1329 & n1362 ) | ( n1329 & ~n1363 ) | ( n1362 & ~n1363 ) ;
  assign n1365 = n1340 ^ n1272 ^ x71 ;
  assign n1366 = n1359 ^ n1272 ^ 1'b0 ;
  assign n1367 = ( n1272 & n1365 ) | ( n1272 & ~n1366 ) | ( n1365 & ~n1366 ) ;
  assign n1368 = n1339 ^ n1275 ^ x70 ;
  assign n1369 = n1359 ^ n1275 ^ 1'b0 ;
  assign n1370 = ( n1275 & n1368 ) | ( n1275 & ~n1369 ) | ( n1368 & ~n1369 ) ;
  assign n1371 = n1337 ^ n1278 ^ x68 ;
  assign n1372 = n1359 ^ n1278 ^ 1'b0 ;
  assign n1373 = ( n1278 & n1371 ) | ( n1278 & ~n1372 ) | ( n1371 & ~n1372 ) ;
  assign n1374 = n1336 ^ n1280 ^ x67 ;
  assign n1375 = n1359 ^ n1280 ^ 1'b0 ;
  assign n1376 = ( n1280 & n1374 ) | ( n1280 & ~n1375 ) | ( n1374 & ~n1375 ) ;
  assign n1377 = n1359 ^ n1335 ^ 1'b0 ;
  assign n1378 = ( n1282 & n1335 ) | ( n1282 & n1377 ) | ( n1335 & n1377 ) ;
  assign n1379 = n1359 ^ n1333 ^ 1'b0 ;
  assign n1380 = ( n1332 & n1333 ) | ( n1332 & n1379 ) | ( n1333 & n1379 ) ;
  assign n1381 = n1355 ^ n1324 ^ x84 ;
  assign n1382 = n1381 ^ n1359 ^ 1'b0 ;
  assign n1383 = ( n1324 & n1381 ) | ( n1324 & n1382 ) | ( n1381 & n1382 ) ;
  assign n1384 = n1359 ^ n1315 ^ 1'b0 ;
  assign n1385 = n1353 ^ n1304 ^ x82 ;
  assign n1386 = n1359 ^ n1304 ^ 1'b0 ;
  assign n1387 = ( n1304 & n1385 ) | ( n1304 & ~n1386 ) | ( n1385 & ~n1386 ) ;
  assign n1388 = n1352 ^ n1308 ^ x81 ;
  assign n1389 = n1359 ^ n1308 ^ 1'b0 ;
  assign n1390 = ( n1308 & n1388 ) | ( n1308 & ~n1389 ) | ( n1388 & ~n1389 ) ;
  assign n1391 = n1351 ^ n1291 ^ x80 ;
  assign n1392 = n1359 ^ n1291 ^ 1'b0 ;
  assign n1393 = ( n1291 & n1391 ) | ( n1291 & ~n1392 ) | ( n1391 & ~n1392 ) ;
  assign n1394 = n1350 ^ n1312 ^ x79 ;
  assign n1395 = n1359 ^ n1312 ^ 1'b0 ;
  assign n1396 = ( n1312 & n1394 ) | ( n1312 & ~n1395 ) | ( n1394 & ~n1395 ) ;
  assign n1397 = n1349 ^ n1325 ^ x78 ;
  assign n1398 = n1359 ^ n1325 ^ 1'b0 ;
  assign n1399 = ( n1325 & n1397 ) | ( n1325 & ~n1398 ) | ( n1397 & ~n1398 ) ;
  assign n1400 = n1348 ^ n1326 ^ x77 ;
  assign n1401 = n1359 ^ n1326 ^ 1'b0 ;
  assign n1402 = ( n1326 & n1400 ) | ( n1326 & ~n1401 ) | ( n1400 & ~n1401 ) ;
  assign n1403 = n1345 ^ n1327 ^ x76 ;
  assign n1404 = n1359 ^ n1327 ^ 1'b0 ;
  assign n1405 = ( n1327 & n1403 ) | ( n1327 & ~n1404 ) | ( n1403 & ~n1404 ) ;
  assign n1406 = n1344 ^ n1320 ^ x75 ;
  assign n1407 = n1359 ^ n1320 ^ 1'b0 ;
  assign n1408 = ( n1320 & n1406 ) | ( n1320 & ~n1407 ) | ( n1406 & ~n1407 ) ;
  assign n1409 = n1342 ^ n1323 ^ x73 ;
  assign n1410 = n1359 ^ n1323 ^ 1'b0 ;
  assign n1411 = ( n1323 & n1409 ) | ( n1323 & ~n1410 ) | ( n1409 & ~n1410 ) ;
  assign n1412 = n1338 ^ n1328 ^ x69 ;
  assign n1413 = n1359 ^ n1328 ^ 1'b0 ;
  assign n1414 = n1354 ^ n1315 ^ x83 ;
  assign n1415 = ( n1315 & ~n1384 ) | ( n1315 & n1414 ) | ( ~n1384 & n1414 ) ;
  assign n1416 = ( n1328 & n1412 ) | ( n1328 & ~n1413 ) | ( n1412 & ~n1413 ) ;
  assign n1417 = n1330 & ~n1359 ;
  assign n1418 = x86 | n1357 ;
  assign n1419 = x42 & x64 ;
  assign n1420 = ~n204 & n1419 ;
  assign n1421 = ~n1418 & n1420 ;
  assign n1422 = ( x42 & n1417 ) | ( x42 & ~n1421 ) | ( n1417 & ~n1421 ) ;
  assign n1423 = ( n322 & n1285 ) | ( n322 & n1359 ) | ( n1285 & n1359 ) ;
  assign n1424 = ~x41 & x64 ;
  assign n1425 = n1424 ^ n1422 ^ x65 ;
  assign n1426 = ( x65 & n1424 ) | ( x65 & n1425 ) | ( n1424 & n1425 ) ;
  assign n1427 = n1426 ^ n1380 ^ x66 ;
  assign n1428 = ( x66 & n1426 ) | ( x66 & n1427 ) | ( n1426 & n1427 ) ;
  assign n1429 = ( x67 & ~n1378 ) | ( x67 & n1428 ) | ( ~n1378 & n1428 ) ;
  assign n1430 = ( x68 & ~n1376 ) | ( x68 & n1429 ) | ( ~n1376 & n1429 ) ;
  assign n1431 = ( x69 & ~n1373 ) | ( x69 & n1430 ) | ( ~n1373 & n1430 ) ;
  assign n1432 = ( x70 & ~n1416 ) | ( x70 & n1431 ) | ( ~n1416 & n1431 ) ;
  assign n1433 = ( x71 & ~n1370 ) | ( x71 & n1432 ) | ( ~n1370 & n1432 ) ;
  assign n1434 = ( x72 & ~n1367 ) | ( x72 & n1433 ) | ( ~n1367 & n1433 ) ;
  assign n1435 = ( x73 & ~n1364 ) | ( x73 & n1434 ) | ( ~n1364 & n1434 ) ;
  assign n1436 = ( x74 & ~n1411 ) | ( x74 & n1435 ) | ( ~n1411 & n1435 ) ;
  assign n1437 = ( x75 & ~n1361 ) | ( x75 & n1436 ) | ( ~n1361 & n1436 ) ;
  assign n1438 = ( x76 & ~n1408 ) | ( x76 & n1437 ) | ( ~n1408 & n1437 ) ;
  assign n1439 = ( x77 & ~n1405 ) | ( x77 & n1438 ) | ( ~n1405 & n1438 ) ;
  assign n1440 = ( x78 & ~n1402 ) | ( x78 & n1439 ) | ( ~n1402 & n1439 ) ;
  assign n1441 = ( x79 & ~n1399 ) | ( x79 & n1440 ) | ( ~n1399 & n1440 ) ;
  assign n1442 = ( x80 & ~n1396 ) | ( x80 & n1441 ) | ( ~n1396 & n1441 ) ;
  assign n1443 = ( x81 & ~n1393 ) | ( x81 & n1442 ) | ( ~n1393 & n1442 ) ;
  assign n1444 = ( x82 & ~n1390 ) | ( x82 & n1443 ) | ( ~n1390 & n1443 ) ;
  assign n1445 = ( x83 & ~n1387 ) | ( x83 & n1444 ) | ( ~n1387 & n1444 ) ;
  assign n1446 = ( x84 & ~n1415 ) | ( x84 & n1445 ) | ( ~n1415 & n1445 ) ;
  assign n1447 = ( x85 & ~n1383 ) | ( x85 & n1446 ) | ( ~n1383 & n1446 ) ;
  assign n1448 = ( x86 & ~n1423 ) | ( x86 & n1447 ) | ( ~n1423 & n1447 ) ;
  assign n1449 = n204 | n1448 ;
  assign n1450 = n1438 ^ n1405 ^ x77 ;
  assign n1451 = n1449 ^ n1405 ^ 1'b0 ;
  assign n1452 = ( n1405 & n1450 ) | ( n1405 & ~n1451 ) | ( n1450 & ~n1451 ) ;
  assign n1453 = n1437 ^ n1408 ^ x76 ;
  assign n1454 = n1449 ^ n1408 ^ 1'b0 ;
  assign n1455 = n1434 ^ n1364 ^ x73 ;
  assign n1456 = n1449 ^ n1364 ^ 1'b0 ;
  assign n1457 = ( n1364 & n1455 ) | ( n1364 & ~n1456 ) | ( n1455 & ~n1456 ) ;
  assign n1458 = n1433 ^ n1367 ^ x72 ;
  assign n1459 = ( n1408 & n1453 ) | ( n1408 & ~n1454 ) | ( n1453 & ~n1454 ) ;
  assign n1460 = n1449 ^ n1367 ^ 1'b0 ;
  assign n1461 = ( n1367 & n1458 ) | ( n1367 & ~n1460 ) | ( n1458 & ~n1460 ) ;
  assign n1462 = n1432 ^ n1370 ^ x71 ;
  assign n1463 = n1449 ^ n1370 ^ 1'b0 ;
  assign n1464 = ( n1370 & n1462 ) | ( n1370 & ~n1463 ) | ( n1462 & ~n1463 ) ;
  assign n1465 = n1431 ^ n1416 ^ x70 ;
  assign n1466 = n1449 ^ n1416 ^ 1'b0 ;
  assign n1467 = ( n1416 & n1465 ) | ( n1416 & ~n1466 ) | ( n1465 & ~n1466 ) ;
  assign n1468 = n1430 ^ n1373 ^ x69 ;
  assign n1469 = n1449 ^ n1373 ^ 1'b0 ;
  assign n1470 = ( n1373 & n1468 ) | ( n1373 & ~n1469 ) | ( n1468 & ~n1469 ) ;
  assign n1471 = n1428 ^ n1378 ^ x67 ;
  assign n1472 = n1449 ^ n1378 ^ 1'b0 ;
  assign n1473 = ( n1378 & n1471 ) | ( n1378 & ~n1472 ) | ( n1471 & ~n1472 ) ;
  assign n1474 = n1449 ^ n1425 ^ 1'b0 ;
  assign n1475 = ( n1422 & n1425 ) | ( n1422 & n1474 ) | ( n1425 & n1474 ) ;
  assign n1476 = n1446 ^ n1383 ^ x85 ;
  assign n1477 = n1476 ^ n1449 ^ 1'b0 ;
  assign n1478 = ( n1383 & n1476 ) | ( n1383 & n1477 ) | ( n1476 & n1477 ) ;
  assign n1479 = n1449 ^ n1415 ^ 1'b0 ;
  assign n1480 = n1445 ^ n1415 ^ x84 ;
  assign n1481 = ( n1415 & ~n1479 ) | ( n1415 & n1480 ) | ( ~n1479 & n1480 ) ;
  assign n1482 = n1444 ^ n1387 ^ x83 ;
  assign n1483 = n1449 ^ n1387 ^ 1'b0 ;
  assign n1484 = ( n1387 & n1482 ) | ( n1387 & ~n1483 ) | ( n1482 & ~n1483 ) ;
  assign n1485 = n1443 ^ n1390 ^ x82 ;
  assign n1486 = n1449 ^ n1390 ^ 1'b0 ;
  assign n1487 = ( n1390 & n1485 ) | ( n1390 & ~n1486 ) | ( n1485 & ~n1486 ) ;
  assign n1488 = n1442 ^ n1393 ^ x81 ;
  assign n1489 = n1449 ^ n1393 ^ 1'b0 ;
  assign n1490 = ( n1393 & n1488 ) | ( n1393 & ~n1489 ) | ( n1488 & ~n1489 ) ;
  assign n1491 = n1441 ^ n1396 ^ x80 ;
  assign n1492 = n1449 ^ n1396 ^ 1'b0 ;
  assign n1493 = ( n1396 & n1491 ) | ( n1396 & ~n1492 ) | ( n1491 & ~n1492 ) ;
  assign n1494 = n1440 ^ n1399 ^ x79 ;
  assign n1495 = n1449 ^ n1399 ^ 1'b0 ;
  assign n1496 = ( n1399 & n1494 ) | ( n1399 & ~n1495 ) | ( n1494 & ~n1495 ) ;
  assign n1497 = n1439 ^ n1402 ^ x78 ;
  assign n1498 = n1449 ^ n1402 ^ 1'b0 ;
  assign n1499 = ( n1402 & n1497 ) | ( n1402 & ~n1498 ) | ( n1497 & ~n1498 ) ;
  assign n1500 = n1436 ^ n1361 ^ x75 ;
  assign n1501 = n1449 ^ n1361 ^ 1'b0 ;
  assign n1502 = ( n1361 & n1500 ) | ( n1361 & ~n1501 ) | ( n1500 & ~n1501 ) ;
  assign n1503 = n1435 ^ n1411 ^ x74 ;
  assign n1504 = n1449 ^ n1411 ^ 1'b0 ;
  assign n1505 = ( n1411 & n1503 ) | ( n1411 & ~n1504 ) | ( n1503 & ~n1504 ) ;
  assign n1506 = n1429 ^ n1376 ^ x68 ;
  assign n1507 = n1449 ^ n1376 ^ 1'b0 ;
  assign n1508 = ( n1376 & n1506 ) | ( n1376 & ~n1507 ) | ( n1506 & ~n1507 ) ;
  assign n1509 = n1449 ^ n1427 ^ 1'b0 ;
  assign n1510 = ( n1380 & n1427 ) | ( n1380 & n1509 ) | ( n1427 & n1509 ) ;
  assign n1511 = n184 | n206 ;
  assign n1512 = n199 | n201 ;
  assign n1513 = x64 & ~x87 ;
  assign n1514 = ( n1511 & ~n1512 ) | ( n1511 & n1513 ) | ( ~n1512 & n1513 ) ;
  assign n1515 = ~n1511 & n1514 ;
  assign n1516 = ( x41 & n1448 ) | ( x41 & ~n1515 ) | ( n1448 & ~n1515 ) ;
  assign n1517 = x41 & ~n1516 ;
  assign n1518 = n1424 & ~n1449 ;
  assign n1519 = ( x41 & ~n1517 ) | ( x41 & n1518 ) | ( ~n1517 & n1518 ) ;
  assign n1520 = n199 | n1511 ;
  assign n1521 = ~x40 & x64 ;
  assign n1522 = n1521 ^ n1519 ^ x65 ;
  assign n1523 = ( x65 & n1521 ) | ( x65 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1524 = n1523 ^ n1475 ^ x66 ;
  assign n1525 = ( x66 & n1523 ) | ( x66 & n1524 ) | ( n1523 & n1524 ) ;
  assign n1526 = ( x67 & ~n1510 ) | ( x67 & n1525 ) | ( ~n1510 & n1525 ) ;
  assign n1527 = ( x68 & ~n1473 ) | ( x68 & n1526 ) | ( ~n1473 & n1526 ) ;
  assign n1528 = ( x69 & ~n1508 ) | ( x69 & n1527 ) | ( ~n1508 & n1527 ) ;
  assign n1529 = ( x70 & ~n1470 ) | ( x70 & n1528 ) | ( ~n1470 & n1528 ) ;
  assign n1530 = ( x71 & ~n1467 ) | ( x71 & n1529 ) | ( ~n1467 & n1529 ) ;
  assign n1531 = ( x72 & ~n1464 ) | ( x72 & n1530 ) | ( ~n1464 & n1530 ) ;
  assign n1532 = ( x73 & ~n1461 ) | ( x73 & n1531 ) | ( ~n1461 & n1531 ) ;
  assign n1533 = ( x74 & ~n1457 ) | ( x74 & n1532 ) | ( ~n1457 & n1532 ) ;
  assign n1534 = ( x75 & ~n1505 ) | ( x75 & n1533 ) | ( ~n1505 & n1533 ) ;
  assign n1535 = ( x76 & ~n1502 ) | ( x76 & n1534 ) | ( ~n1502 & n1534 ) ;
  assign n1536 = ( x77 & ~n1459 ) | ( x77 & n1535 ) | ( ~n1459 & n1535 ) ;
  assign n1537 = ( x78 & ~n1452 ) | ( x78 & n1536 ) | ( ~n1452 & n1536 ) ;
  assign n1538 = ( x79 & ~n1499 ) | ( x79 & n1537 ) | ( ~n1499 & n1537 ) ;
  assign n1539 = ( x80 & ~n1496 ) | ( x80 & n1538 ) | ( ~n1496 & n1538 ) ;
  assign n1540 = ( x81 & ~n1493 ) | ( x81 & n1539 ) | ( ~n1493 & n1539 ) ;
  assign n1541 = ( x82 & ~n1490 ) | ( x82 & n1540 ) | ( ~n1490 & n1540 ) ;
  assign n1542 = ( x83 & ~n1487 ) | ( x83 & n1541 ) | ( ~n1487 & n1541 ) ;
  assign n1543 = ( x84 & ~n1484 ) | ( x84 & n1542 ) | ( ~n1484 & n1542 ) ;
  assign n1544 = ( x85 & ~n1481 ) | ( x85 & n1543 ) | ( ~n1481 & n1543 ) ;
  assign n1545 = n1544 ^ n1478 ^ x86 ;
  assign n1546 = n1423 & n1449 ;
  assign n1547 = n322 | n1546 ;
  assign n1548 = ( x86 & ~n1478 ) | ( x86 & n1544 ) | ( ~n1478 & n1544 ) ;
  assign n1549 = ( x87 & n984 ) | ( x87 & ~n1546 ) | ( n984 & ~n1546 ) ;
  assign n1550 = ( ~x87 & n984 ) | ( ~x87 & n1547 ) | ( n984 & n1547 ) ;
  assign n1551 = ( ~n1548 & n1549 ) | ( ~n1548 & n1550 ) | ( n1549 & n1550 ) ;
  assign n1552 = n1548 | n1551 ;
  assign n1553 = n204 & n1547 ;
  assign n1554 = ( ~n1547 & n1552 ) | ( ~n1547 & n1553 ) | ( n1552 & n1553 ) ;
  assign n1555 = n1554 ^ n1478 ^ 1'b0 ;
  assign n1556 = ( n1478 & n1545 ) | ( n1478 & ~n1555 ) | ( n1545 & ~n1555 ) ;
  assign n1557 = n1543 ^ n1481 ^ x85 ;
  assign n1558 = n1554 ^ n1481 ^ 1'b0 ;
  assign n1559 = ( n1481 & n1557 ) | ( n1481 & ~n1558 ) | ( n1557 & ~n1558 ) ;
  assign n1560 = n1542 ^ n1484 ^ x84 ;
  assign n1561 = n1554 ^ n1484 ^ 1'b0 ;
  assign n1562 = ( n1484 & n1560 ) | ( n1484 & ~n1561 ) | ( n1560 & ~n1561 ) ;
  assign n1563 = n1531 ^ n1461 ^ x73 ;
  assign n1564 = n1554 ^ n1461 ^ 1'b0 ;
  assign n1565 = ( n1461 & n1563 ) | ( n1461 & ~n1564 ) | ( n1563 & ~n1564 ) ;
  assign n1566 = n1525 ^ n1510 ^ x67 ;
  assign n1567 = n1554 ^ n1510 ^ 1'b0 ;
  assign n1568 = ( n1510 & n1566 ) | ( n1510 & ~n1567 ) | ( n1566 & ~n1567 ) ;
  assign n1569 = n1554 ^ n1524 ^ 1'b0 ;
  assign n1570 = ( n1475 & n1524 ) | ( n1475 & n1569 ) | ( n1524 & n1569 ) ;
  assign n1571 = n1554 ^ n1522 ^ 1'b0 ;
  assign n1572 = ( n1519 & n1522 ) | ( n1519 & n1571 ) | ( n1522 & n1571 ) ;
  assign n1573 = ( n204 & n322 ) | ( n204 & n1423 ) | ( n322 & n1423 ) ;
  assign n1574 = n322 | n1552 ;
  assign n1575 = ( n322 & n1573 ) | ( n322 & n1574 ) | ( n1573 & n1574 ) ;
  assign n1576 = n1541 ^ n1487 ^ x83 ;
  assign n1577 = n1554 ^ n1487 ^ 1'b0 ;
  assign n1578 = ( n1487 & n1576 ) | ( n1487 & ~n1577 ) | ( n1576 & ~n1577 ) ;
  assign n1579 = n1540 ^ n1490 ^ x82 ;
  assign n1580 = n1554 ^ n1490 ^ 1'b0 ;
  assign n1581 = ( n1490 & n1579 ) | ( n1490 & ~n1580 ) | ( n1579 & ~n1580 ) ;
  assign n1582 = n1539 ^ n1493 ^ x81 ;
  assign n1583 = n1554 ^ n1493 ^ 1'b0 ;
  assign n1584 = ( n1493 & n1582 ) | ( n1493 & ~n1583 ) | ( n1582 & ~n1583 ) ;
  assign n1585 = n1538 ^ n1496 ^ x80 ;
  assign n1586 = n1554 ^ n1496 ^ 1'b0 ;
  assign n1587 = ( n1496 & n1585 ) | ( n1496 & ~n1586 ) | ( n1585 & ~n1586 ) ;
  assign n1588 = n1537 ^ n1499 ^ x79 ;
  assign n1589 = n1554 ^ n1499 ^ 1'b0 ;
  assign n1590 = ( n1499 & n1588 ) | ( n1499 & ~n1589 ) | ( n1588 & ~n1589 ) ;
  assign n1591 = n1536 ^ n1452 ^ x78 ;
  assign n1592 = n1554 ^ n1452 ^ 1'b0 ;
  assign n1593 = ( n1452 & n1591 ) | ( n1452 & ~n1592 ) | ( n1591 & ~n1592 ) ;
  assign n1594 = n1535 ^ n1459 ^ x77 ;
  assign n1595 = n1554 ^ n1459 ^ 1'b0 ;
  assign n1596 = ( n1459 & n1594 ) | ( n1459 & ~n1595 ) | ( n1594 & ~n1595 ) ;
  assign n1597 = n1534 ^ n1502 ^ x76 ;
  assign n1598 = n1554 ^ n1502 ^ 1'b0 ;
  assign n1599 = ( n1502 & n1597 ) | ( n1502 & ~n1598 ) | ( n1597 & ~n1598 ) ;
  assign n1600 = n1533 ^ n1505 ^ x75 ;
  assign n1601 = n1554 ^ n1505 ^ 1'b0 ;
  assign n1602 = ( n1505 & n1600 ) | ( n1505 & ~n1601 ) | ( n1600 & ~n1601 ) ;
  assign n1603 = n1532 ^ n1457 ^ x74 ;
  assign n1604 = n1554 ^ n1457 ^ 1'b0 ;
  assign n1605 = ( n1457 & n1603 ) | ( n1457 & ~n1604 ) | ( n1603 & ~n1604 ) ;
  assign n1606 = n1530 ^ n1464 ^ x72 ;
  assign n1607 = n1554 ^ n1464 ^ 1'b0 ;
  assign n1608 = ( n1464 & n1606 ) | ( n1464 & ~n1607 ) | ( n1606 & ~n1607 ) ;
  assign n1609 = n1529 ^ n1467 ^ x71 ;
  assign n1610 = n1554 ^ n1467 ^ 1'b0 ;
  assign n1611 = ( n1467 & n1609 ) | ( n1467 & ~n1610 ) | ( n1609 & ~n1610 ) ;
  assign n1612 = n1528 ^ n1470 ^ x70 ;
  assign n1613 = n1554 ^ n1470 ^ 1'b0 ;
  assign n1614 = ( n1470 & n1612 ) | ( n1470 & ~n1613 ) | ( n1612 & ~n1613 ) ;
  assign n1615 = n1527 ^ n1508 ^ x69 ;
  assign n1616 = n1554 ^ n1508 ^ 1'b0 ;
  assign n1617 = ( n1508 & n1615 ) | ( n1508 & ~n1616 ) | ( n1615 & ~n1616 ) ;
  assign n1618 = n1526 ^ n1473 ^ x68 ;
  assign n1619 = n1554 ^ n1473 ^ 1'b0 ;
  assign n1620 = ( n1473 & n1618 ) | ( n1473 & ~n1619 ) | ( n1618 & ~n1619 ) ;
  assign n1621 = x64 & n1554 ;
  assign n1622 = ~x39 & x64 ;
  assign n1623 = n1621 ^ x64 ^ x40 ;
  assign n1624 = n1623 ^ n1622 ^ x65 ;
  assign n1625 = ( x65 & n1622 ) | ( x65 & n1624 ) | ( n1622 & n1624 ) ;
  assign n1626 = n1625 ^ n1572 ^ x66 ;
  assign n1627 = ( x66 & n1625 ) | ( x66 & n1626 ) | ( n1625 & n1626 ) ;
  assign n1628 = ( x67 & ~n1570 ) | ( x67 & n1627 ) | ( ~n1570 & n1627 ) ;
  assign n1629 = ( x68 & ~n1568 ) | ( x68 & n1628 ) | ( ~n1568 & n1628 ) ;
  assign n1630 = ( x69 & ~n1620 ) | ( x69 & n1629 ) | ( ~n1620 & n1629 ) ;
  assign n1631 = ( x70 & ~n1617 ) | ( x70 & n1630 ) | ( ~n1617 & n1630 ) ;
  assign n1632 = ( x71 & ~n1614 ) | ( x71 & n1631 ) | ( ~n1614 & n1631 ) ;
  assign n1633 = ( x72 & ~n1611 ) | ( x72 & n1632 ) | ( ~n1611 & n1632 ) ;
  assign n1634 = ( x73 & ~n1608 ) | ( x73 & n1633 ) | ( ~n1608 & n1633 ) ;
  assign n1635 = ( x74 & ~n1565 ) | ( x74 & n1634 ) | ( ~n1565 & n1634 ) ;
  assign n1636 = ( x75 & ~n1605 ) | ( x75 & n1635 ) | ( ~n1605 & n1635 ) ;
  assign n1637 = ( x76 & ~n1602 ) | ( x76 & n1636 ) | ( ~n1602 & n1636 ) ;
  assign n1638 = ( x77 & ~n1599 ) | ( x77 & n1637 ) | ( ~n1599 & n1637 ) ;
  assign n1639 = ( x78 & ~n1596 ) | ( x78 & n1638 ) | ( ~n1596 & n1638 ) ;
  assign n1640 = ( x79 & ~n1593 ) | ( x79 & n1639 ) | ( ~n1593 & n1639 ) ;
  assign n1641 = n1630 ^ n1617 ^ x70 ;
  assign n1642 = ( x80 & ~n1590 ) | ( x80 & n1640 ) | ( ~n1590 & n1640 ) ;
  assign n1643 = ( x81 & ~n1587 ) | ( x81 & n1642 ) | ( ~n1587 & n1642 ) ;
  assign n1644 = n1638 ^ n1596 ^ x78 ;
  assign n1645 = ( x82 & ~n1584 ) | ( x82 & n1643 ) | ( ~n1584 & n1643 ) ;
  assign n1646 = ( x83 & ~n1581 ) | ( x83 & n1645 ) | ( ~n1581 & n1645 ) ;
  assign n1647 = ( x84 & ~n1578 ) | ( x84 & n1646 ) | ( ~n1578 & n1646 ) ;
  assign n1648 = ( x85 & ~n1562 ) | ( x85 & n1647 ) | ( ~n1562 & n1647 ) ;
  assign n1649 = ( x86 & ~n1559 ) | ( x86 & n1648 ) | ( ~n1559 & n1648 ) ;
  assign n1650 = ( x87 & ~n1556 ) | ( x87 & n1649 ) | ( ~n1556 & n1649 ) ;
  assign n1651 = ~n178 & n1622 ;
  assign n1652 = ( x88 & ~n1575 ) | ( x88 & n1650 ) | ( ~n1575 & n1650 ) ;
  assign n1653 = n203 | n1652 ;
  assign n1654 = n1653 ^ n1617 ^ 1'b0 ;
  assign n1655 = ( n1617 & n1641 ) | ( n1617 & ~n1654 ) | ( n1641 & ~n1654 ) ;
  assign n1656 = n1637 ^ n1599 ^ x77 ;
  assign n1657 = n1653 ^ n1624 ^ 1'b0 ;
  assign n1658 = n1653 ^ n1596 ^ 1'b0 ;
  assign n1659 = ( n1596 & n1644 ) | ( n1596 & ~n1658 ) | ( n1644 & ~n1658 ) ;
  assign n1660 = n1653 ^ n1599 ^ 1'b0 ;
  assign n1661 = ( n1599 & n1656 ) | ( n1599 & ~n1660 ) | ( n1656 & ~n1660 ) ;
  assign n1662 = n1653 ^ n1626 ^ 1'b0 ;
  assign n1663 = n1653 ^ n1614 ^ 1'b0 ;
  assign n1664 = ( n1572 & n1626 ) | ( n1572 & n1662 ) | ( n1626 & n1662 ) ;
  assign n1665 = n1631 ^ n1614 ^ x71 ;
  assign n1666 = ( n1614 & ~n1663 ) | ( n1614 & n1665 ) | ( ~n1663 & n1665 ) ;
  assign n1667 = n1628 ^ n1568 ^ x68 ;
  assign n1668 = n1653 ^ n1568 ^ 1'b0 ;
  assign n1669 = ( n1568 & n1667 ) | ( n1568 & ~n1668 ) | ( n1667 & ~n1668 ) ;
  assign n1670 = n1627 ^ n1570 ^ x67 ;
  assign n1671 = n1653 ^ n1570 ^ 1'b0 ;
  assign n1672 = ( n1570 & n1670 ) | ( n1570 & ~n1671 ) | ( n1670 & ~n1671 ) ;
  assign n1673 = ( n1623 & n1624 ) | ( n1623 & n1657 ) | ( n1624 & n1657 ) ;
  assign n1674 = n1649 ^ n1556 ^ x87 ;
  assign n1675 = n1674 ^ n1653 ^ 1'b0 ;
  assign n1676 = ( n1556 & n1674 ) | ( n1556 & n1675 ) | ( n1674 & n1675 ) ;
  assign n1677 = n1648 ^ n1559 ^ x86 ;
  assign n1678 = n1653 ^ n1559 ^ 1'b0 ;
  assign n1679 = ( n1559 & n1677 ) | ( n1559 & ~n1678 ) | ( n1677 & ~n1678 ) ;
  assign n1680 = n1647 ^ n1562 ^ x85 ;
  assign n1681 = n1653 ^ n1562 ^ 1'b0 ;
  assign n1682 = ( n1562 & n1680 ) | ( n1562 & ~n1681 ) | ( n1680 & ~n1681 ) ;
  assign n1683 = n1646 ^ n1578 ^ x84 ;
  assign n1684 = n1653 ^ n1578 ^ 1'b0 ;
  assign n1685 = ( n1578 & n1683 ) | ( n1578 & ~n1684 ) | ( n1683 & ~n1684 ) ;
  assign n1686 = n1645 ^ n1581 ^ x83 ;
  assign n1687 = n1653 ^ n1581 ^ 1'b0 ;
  assign n1688 = ( n1581 & n1686 ) | ( n1581 & ~n1687 ) | ( n1686 & ~n1687 ) ;
  assign n1689 = n1643 ^ n1584 ^ x82 ;
  assign n1690 = n1653 ^ n1584 ^ 1'b0 ;
  assign n1691 = ( n1584 & n1689 ) | ( n1584 & ~n1690 ) | ( n1689 & ~n1690 ) ;
  assign n1692 = n1642 ^ n1587 ^ x81 ;
  assign n1693 = n1653 ^ n1587 ^ 1'b0 ;
  assign n1694 = ( n1587 & n1692 ) | ( n1587 & ~n1693 ) | ( n1692 & ~n1693 ) ;
  assign n1695 = n1640 ^ n1590 ^ x80 ;
  assign n1696 = n1653 ^ n1590 ^ 1'b0 ;
  assign n1697 = ( n1590 & n1695 ) | ( n1590 & ~n1696 ) | ( n1695 & ~n1696 ) ;
  assign n1698 = n1639 ^ n1593 ^ x79 ;
  assign n1699 = n1653 ^ n1593 ^ 1'b0 ;
  assign n1700 = ( n1593 & n1698 ) | ( n1593 & ~n1699 ) | ( n1698 & ~n1699 ) ;
  assign n1701 = n1636 ^ n1602 ^ x76 ;
  assign n1702 = n1653 ^ n1602 ^ 1'b0 ;
  assign n1703 = ( n1602 & n1701 ) | ( n1602 & ~n1702 ) | ( n1701 & ~n1702 ) ;
  assign n1704 = n1635 ^ n1605 ^ x75 ;
  assign n1705 = n1653 ^ n1605 ^ 1'b0 ;
  assign n1706 = ( n1605 & n1704 ) | ( n1605 & ~n1705 ) | ( n1704 & ~n1705 ) ;
  assign n1707 = n1634 ^ n1565 ^ x74 ;
  assign n1708 = n1653 ^ n1565 ^ 1'b0 ;
  assign n1709 = ( n1565 & n1707 ) | ( n1565 & ~n1708 ) | ( n1707 & ~n1708 ) ;
  assign n1710 = n1633 ^ n1608 ^ x73 ;
  assign n1711 = n1653 ^ n1608 ^ 1'b0 ;
  assign n1712 = ( n1608 & n1710 ) | ( n1608 & ~n1711 ) | ( n1710 & ~n1711 ) ;
  assign n1713 = n1632 ^ n1611 ^ x72 ;
  assign n1714 = n1653 ^ n1611 ^ 1'b0 ;
  assign n1715 = ( n1611 & n1713 ) | ( n1611 & ~n1714 ) | ( n1713 & ~n1714 ) ;
  assign n1716 = n1629 ^ n1620 ^ x69 ;
  assign n1717 = n1653 ^ n1620 ^ 1'b0 ;
  assign n1718 = ( n1620 & n1716 ) | ( n1620 & ~n1717 ) | ( n1716 & ~n1717 ) ;
  assign n1719 = x39 & x64 ;
  assign n1720 = ~x38 & x64 ;
  assign n1721 = x90 | x91 ;
  assign n1722 = x89 | n1652 ;
  assign n1723 = ( ~n184 & n243 ) | ( ~n184 & n1721 ) | ( n243 & n1721 ) ;
  assign n1724 = n184 | n1723 ;
  assign n1725 = n1719 & ~n1724 ;
  assign n1726 = ~n1722 & n1725 ;
  assign n1727 = n175 | n202 ;
  assign n1728 = n1651 & ~n1727 ;
  assign n1729 = ~n1652 & n1728 ;
  assign n1730 = ( x39 & ~n1726 ) | ( x39 & n1729 ) | ( ~n1726 & n1729 ) ;
  assign n1731 = n1730 ^ n1720 ^ x65 ;
  assign n1732 = ( x65 & n1720 ) | ( x65 & n1731 ) | ( n1720 & n1731 ) ;
  assign n1733 = n1732 ^ n1673 ^ x66 ;
  assign n1734 = ( x66 & n1732 ) | ( x66 & n1733 ) | ( n1732 & n1733 ) ;
  assign n1735 = ( x67 & ~n1664 ) | ( x67 & n1734 ) | ( ~n1664 & n1734 ) ;
  assign n1736 = n1735 ^ n1672 ^ x68 ;
  assign n1737 = ( n322 & n1575 ) | ( n322 & n1653 ) | ( n1575 & n1653 ) ;
  assign n1738 = n1734 ^ n1664 ^ x67 ;
  assign n1739 = ( x68 & ~n1672 ) | ( x68 & n1735 ) | ( ~n1672 & n1735 ) ;
  assign n1740 = ( x69 & ~n1669 ) | ( x69 & n1739 ) | ( ~n1669 & n1739 ) ;
  assign n1741 = ( x70 & ~n1718 ) | ( x70 & n1740 ) | ( ~n1718 & n1740 ) ;
  assign n1742 = ( x71 & ~n1655 ) | ( x71 & n1741 ) | ( ~n1655 & n1741 ) ;
  assign n1743 = ( x72 & ~n1666 ) | ( x72 & n1742 ) | ( ~n1666 & n1742 ) ;
  assign n1744 = n1739 ^ n1669 ^ x69 ;
  assign n1745 = ( x73 & ~n1715 ) | ( x73 & n1743 ) | ( ~n1715 & n1743 ) ;
  assign n1746 = ( x74 & ~n1712 ) | ( x74 & n1745 ) | ( ~n1712 & n1745 ) ;
  assign n1747 = ( x75 & ~n1709 ) | ( x75 & n1746 ) | ( ~n1709 & n1746 ) ;
  assign n1748 = ( x76 & ~n1706 ) | ( x76 & n1747 ) | ( ~n1706 & n1747 ) ;
  assign n1749 = ( x77 & ~n1703 ) | ( x77 & n1748 ) | ( ~n1703 & n1748 ) ;
  assign n1750 = ( x78 & ~n1661 ) | ( x78 & n1749 ) | ( ~n1661 & n1749 ) ;
  assign n1751 = ( x79 & ~n1659 ) | ( x79 & n1750 ) | ( ~n1659 & n1750 ) ;
  assign n1752 = n1751 ^ n1700 ^ x80 ;
  assign n1753 = ( x80 & ~n1700 ) | ( x80 & n1751 ) | ( ~n1700 & n1751 ) ;
  assign n1754 = n1753 ^ n1697 ^ x81 ;
  assign n1755 = ( x81 & ~n1697 ) | ( x81 & n1753 ) | ( ~n1697 & n1753 ) ;
  assign n1756 = ( x82 & ~n1694 ) | ( x82 & n1755 ) | ( ~n1694 & n1755 ) ;
  assign n1757 = ( x83 & ~n1691 ) | ( x83 & n1756 ) | ( ~n1691 & n1756 ) ;
  assign n1758 = ( x84 & ~n1688 ) | ( x84 & n1757 ) | ( ~n1688 & n1757 ) ;
  assign n1759 = ( x85 & ~n1685 ) | ( x85 & n1758 ) | ( ~n1685 & n1758 ) ;
  assign n1760 = ( x86 & ~n1682 ) | ( x86 & n1759 ) | ( ~n1682 & n1759 ) ;
  assign n1761 = ( x87 & ~n1679 ) | ( x87 & n1760 ) | ( ~n1679 & n1760 ) ;
  assign n1762 = n1761 ^ n1676 ^ x88 ;
  assign n1763 = ( x88 & ~n1676 ) | ( x88 & n1761 ) | ( ~n1676 & n1761 ) ;
  assign n1764 = ( x89 & ~n1737 ) | ( x89 & n1763 ) | ( ~n1737 & n1763 ) ;
  assign n1765 = n1724 | n1764 ;
  assign n1766 = n1765 ^ n1762 ^ 1'b0 ;
  assign n1767 = ( n1676 & n1762 ) | ( n1676 & n1766 ) | ( n1762 & n1766 ) ;
  assign n1768 = n1760 ^ n1679 ^ x87 ;
  assign n1769 = n1765 ^ n1679 ^ 1'b0 ;
  assign n1770 = ( n1679 & n1768 ) | ( n1679 & ~n1769 ) | ( n1768 & ~n1769 ) ;
  assign n1771 = n1765 ^ n1682 ^ 1'b0 ;
  assign n1772 = n1758 ^ n1685 ^ x85 ;
  assign n1773 = n1765 ^ n1685 ^ 1'b0 ;
  assign n1774 = ( n1685 & n1772 ) | ( n1685 & ~n1773 ) | ( n1772 & ~n1773 ) ;
  assign n1775 = n1757 ^ n1688 ^ x84 ;
  assign n1776 = n1765 ^ n1688 ^ 1'b0 ;
  assign n1777 = ( n1688 & n1775 ) | ( n1688 & ~n1776 ) | ( n1775 & ~n1776 ) ;
  assign n1778 = n1756 ^ n1691 ^ x83 ;
  assign n1779 = n1765 ^ n1691 ^ 1'b0 ;
  assign n1780 = ( n1691 & n1778 ) | ( n1691 & ~n1779 ) | ( n1778 & ~n1779 ) ;
  assign n1781 = n1755 ^ n1694 ^ x82 ;
  assign n1782 = n1765 ^ n1694 ^ 1'b0 ;
  assign n1783 = ( n1694 & n1781 ) | ( n1694 & ~n1782 ) | ( n1781 & ~n1782 ) ;
  assign n1784 = n1765 ^ n1697 ^ 1'b0 ;
  assign n1785 = ( n1697 & n1754 ) | ( n1697 & ~n1784 ) | ( n1754 & ~n1784 ) ;
  assign n1786 = n1765 ^ n1700 ^ 1'b0 ;
  assign n1787 = ( n1700 & n1752 ) | ( n1700 & ~n1786 ) | ( n1752 & ~n1786 ) ;
  assign n1788 = n1765 ^ n1669 ^ 1'b0 ;
  assign n1789 = ( n1669 & n1744 ) | ( n1669 & ~n1788 ) | ( n1744 & ~n1788 ) ;
  assign n1790 = n1765 ^ n1672 ^ 1'b0 ;
  assign n1791 = n1759 ^ n1682 ^ x86 ;
  assign n1792 = ( n1682 & ~n1771 ) | ( n1682 & n1791 ) | ( ~n1771 & n1791 ) ;
  assign n1793 = ( n1672 & n1736 ) | ( n1672 & ~n1790 ) | ( n1736 & ~n1790 ) ;
  assign n1794 = n1765 ^ n1664 ^ 1'b0 ;
  assign n1795 = ( n1664 & n1738 ) | ( n1664 & ~n1794 ) | ( n1738 & ~n1794 ) ;
  assign n1796 = n1765 ^ n1733 ^ 1'b0 ;
  assign n1797 = ( n1673 & n1733 ) | ( n1673 & n1796 ) | ( n1733 & n1796 ) ;
  assign n1798 = n1765 ^ n1731 ^ 1'b0 ;
  assign n1799 = ( n1730 & n1731 ) | ( n1730 & n1798 ) | ( n1731 & n1798 ) ;
  assign n1800 = n1741 ^ n1655 ^ x71 ;
  assign n1801 = n1765 ^ n1661 ^ 1'b0 ;
  assign n1802 = n1765 ^ n1659 ^ 1'b0 ;
  assign n1803 = n1765 ^ n1706 ^ 1'b0 ;
  assign n1804 = n1765 ^ n1712 ^ 1'b0 ;
  assign n1805 = n1746 ^ n1709 ^ x75 ;
  assign n1806 = n1765 ^ n1709 ^ 1'b0 ;
  assign n1807 = n1749 ^ n1661 ^ x78 ;
  assign n1808 = n1750 ^ n1659 ^ x79 ;
  assign n1809 = n1720 & ~n1765 ;
  assign n1810 = ( n1659 & ~n1802 ) | ( n1659 & n1808 ) | ( ~n1802 & n1808 ) ;
  assign n1811 = n1765 ^ n1655 ^ 1'b0 ;
  assign n1812 = ( n1655 & n1800 ) | ( n1655 & ~n1811 ) | ( n1800 & ~n1811 ) ;
  assign n1813 = n1743 ^ n1715 ^ x73 ;
  assign n1814 = x90 | n1764 ;
  assign n1815 = n1742 ^ n1666 ^ x72 ;
  assign n1816 = n1765 ^ n1666 ^ 1'b0 ;
  assign n1817 = ( n1666 & n1815 ) | ( n1666 & ~n1816 ) | ( n1815 & ~n1816 ) ;
  assign n1818 = n1765 ^ n1715 ^ 1'b0 ;
  assign n1819 = ( n1715 & n1813 ) | ( n1715 & ~n1818 ) | ( n1813 & ~n1818 ) ;
  assign n1820 = ~x37 & x64 ;
  assign n1821 = x38 & x64 ;
  assign n1822 = n146 | n1727 ;
  assign n1823 = n1821 & ~n1822 ;
  assign n1824 = ~n1814 & n1823 ;
  assign n1825 = ( x38 & n1809 ) | ( x38 & ~n1824 ) | ( n1809 & ~n1824 ) ;
  assign n1826 = n1825 ^ n1820 ^ x65 ;
  assign n1827 = ( x65 & n1820 ) | ( x65 & n1826 ) | ( n1820 & n1826 ) ;
  assign n1828 = n1827 ^ n1799 ^ x66 ;
  assign n1829 = ( x66 & n1827 ) | ( x66 & n1828 ) | ( n1827 & n1828 ) ;
  assign n1830 = ( x67 & ~n1797 ) | ( x67 & n1829 ) | ( ~n1797 & n1829 ) ;
  assign n1831 = ( x68 & ~n1795 ) | ( x68 & n1830 ) | ( ~n1795 & n1830 ) ;
  assign n1832 = ( n1709 & n1805 ) | ( n1709 & ~n1806 ) | ( n1805 & ~n1806 ) ;
  assign n1833 = ( x69 & ~n1793 ) | ( x69 & n1831 ) | ( ~n1793 & n1831 ) ;
  assign n1834 = ( x70 & ~n1789 ) | ( x70 & n1833 ) | ( ~n1789 & n1833 ) ;
  assign n1835 = n1765 ^ n1718 ^ 1'b0 ;
  assign n1836 = n1740 ^ n1718 ^ x70 ;
  assign n1837 = ( n1718 & ~n1835 ) | ( n1718 & n1836 ) | ( ~n1835 & n1836 ) ;
  assign n1838 = ( x71 & n1834 ) | ( x71 & ~n1837 ) | ( n1834 & ~n1837 ) ;
  assign n1839 = ( x72 & ~n1812 ) | ( x72 & n1838 ) | ( ~n1812 & n1838 ) ;
  assign n1840 = n1745 ^ n1712 ^ x74 ;
  assign n1841 = ( n1712 & ~n1804 ) | ( n1712 & n1840 ) | ( ~n1804 & n1840 ) ;
  assign n1842 = ( n1661 & ~n1801 ) | ( n1661 & n1807 ) | ( ~n1801 & n1807 ) ;
  assign n1843 = n1747 ^ n1706 ^ x76 ;
  assign n1844 = ( n1706 & ~n1803 ) | ( n1706 & n1843 ) | ( ~n1803 & n1843 ) ;
  assign n1845 = n1765 ^ n1703 ^ 1'b0 ;
  assign n1846 = n1748 ^ n1703 ^ x77 ;
  assign n1847 = ( n1703 & ~n1845 ) | ( n1703 & n1846 ) | ( ~n1845 & n1846 ) ;
  assign n1848 = ( x73 & ~n1817 ) | ( x73 & n1839 ) | ( ~n1817 & n1839 ) ;
  assign n1849 = ( x74 & ~n1819 ) | ( x74 & n1848 ) | ( ~n1819 & n1848 ) ;
  assign n1850 = ( x75 & ~n1841 ) | ( x75 & n1849 ) | ( ~n1841 & n1849 ) ;
  assign n1851 = ( x76 & ~n1832 ) | ( x76 & n1850 ) | ( ~n1832 & n1850 ) ;
  assign n1852 = ( x77 & ~n1844 ) | ( x77 & n1851 ) | ( ~n1844 & n1851 ) ;
  assign n1853 = ( x78 & ~n1847 ) | ( x78 & n1852 ) | ( ~n1847 & n1852 ) ;
  assign n1854 = n1829 ^ n1797 ^ x67 ;
  assign n1855 = n1830 ^ n1795 ^ x68 ;
  assign n1856 = n1831 ^ n1793 ^ x69 ;
  assign n1857 = ( x79 & ~n1842 ) | ( x79 & n1853 ) | ( ~n1842 & n1853 ) ;
  assign n1858 = n1837 ^ n1834 ^ x71 ;
  assign n1859 = n1838 ^ n1812 ^ x72 ;
  assign n1860 = n1839 ^ n1817 ^ x73 ;
  assign n1861 = n1848 ^ n1819 ^ x74 ;
  assign n1862 = n1833 ^ n1789 ^ x70 ;
  assign n1863 = n1850 ^ n1832 ^ x76 ;
  assign n1864 = n1851 ^ n1844 ^ x77 ;
  assign n1865 = n1852 ^ n1847 ^ x78 ;
  assign n1866 = n1853 ^ n1842 ^ x79 ;
  assign n1867 = n1849 ^ n1841 ^ x75 ;
  assign n1868 = ( x80 & ~n1810 ) | ( x80 & n1857 ) | ( ~n1810 & n1857 ) ;
  assign n1869 = ( x81 & ~n1787 ) | ( x81 & n1868 ) | ( ~n1787 & n1868 ) ;
  assign n1870 = ( x82 & ~n1785 ) | ( x82 & n1869 ) | ( ~n1785 & n1869 ) ;
  assign n1871 = ( x83 & ~n1783 ) | ( x83 & n1870 ) | ( ~n1783 & n1870 ) ;
  assign n1872 = ( x84 & ~n1780 ) | ( x84 & n1871 ) | ( ~n1780 & n1871 ) ;
  assign n1873 = ( x85 & ~n1777 ) | ( x85 & n1872 ) | ( ~n1777 & n1872 ) ;
  assign n1874 = ( x86 & ~n1774 ) | ( x86 & n1873 ) | ( ~n1774 & n1873 ) ;
  assign n1875 = ( x87 & ~n1792 ) | ( x87 & n1874 ) | ( ~n1792 & n1874 ) ;
  assign n1876 = ( x88 & ~n1770 ) | ( x88 & n1875 ) | ( ~n1770 & n1875 ) ;
  assign n1877 = n1737 & n1765 ;
  assign n1878 = n322 | n1877 ;
  assign n1879 = ( x89 & ~n1767 ) | ( x89 & n1876 ) | ( ~n1767 & n1876 ) ;
  assign n1880 = ( x90 & n1822 ) | ( x90 & ~n1877 ) | ( n1822 & ~n1877 ) ;
  assign n1881 = ( ~x90 & n1822 ) | ( ~x90 & n1878 ) | ( n1822 & n1878 ) ;
  assign n1882 = ( ~n1879 & n1880 ) | ( ~n1879 & n1881 ) | ( n1880 & n1881 ) ;
  assign n1883 = n1879 | n1882 ;
  assign n1884 = n1724 & n1878 ;
  assign n1885 = ( ~n1878 & n1883 ) | ( ~n1878 & n1884 ) | ( n1883 & n1884 ) ;
  assign n1886 = n1885 ^ n1842 ^ 1'b0 ;
  assign n1887 = ( n1842 & n1866 ) | ( n1842 & ~n1886 ) | ( n1866 & ~n1886 ) ;
  assign n1888 = n1885 ^ n1847 ^ 1'b0 ;
  assign n1889 = ( n1847 & n1865 ) | ( n1847 & ~n1888 ) | ( n1865 & ~n1888 ) ;
  assign n1890 = n1885 ^ n1844 ^ 1'b0 ;
  assign n1891 = ( n1844 & n1864 ) | ( n1844 & ~n1890 ) | ( n1864 & ~n1890 ) ;
  assign n1892 = n1885 ^ n1832 ^ 1'b0 ;
  assign n1893 = ( n1832 & n1863 ) | ( n1832 & ~n1892 ) | ( n1863 & ~n1892 ) ;
  assign n1894 = n1885 ^ n1841 ^ 1'b0 ;
  assign n1895 = ( n1841 & n1867 ) | ( n1841 & ~n1894 ) | ( n1867 & ~n1894 ) ;
  assign n1896 = n1885 ^ n1819 ^ 1'b0 ;
  assign n1897 = ( n1819 & n1861 ) | ( n1819 & ~n1896 ) | ( n1861 & ~n1896 ) ;
  assign n1898 = n1885 ^ n1789 ^ 1'b0 ;
  assign n1899 = ( n1789 & n1862 ) | ( n1789 & ~n1898 ) | ( n1862 & ~n1898 ) ;
  assign n1900 = n1885 ^ n1793 ^ 1'b0 ;
  assign n1901 = ( n1793 & n1856 ) | ( n1793 & ~n1900 ) | ( n1856 & ~n1900 ) ;
  assign n1902 = n1885 ^ n1795 ^ 1'b0 ;
  assign n1903 = ( n1795 & n1855 ) | ( n1795 & ~n1902 ) | ( n1855 & ~n1902 ) ;
  assign n1904 = n1885 ^ n1797 ^ 1'b0 ;
  assign n1905 = ( n1797 & n1854 ) | ( n1797 & ~n1904 ) | ( n1854 & ~n1904 ) ;
  assign n1906 = n1885 ^ n1828 ^ 1'b0 ;
  assign n1907 = ( n1799 & n1828 ) | ( n1799 & n1906 ) | ( n1828 & n1906 ) ;
  assign n1908 = n1885 ^ n1826 ^ 1'b0 ;
  assign n1909 = ( n1825 & n1826 ) | ( n1825 & n1908 ) | ( n1826 & n1908 ) ;
  assign n1910 = ( n322 & n1737 ) | ( n322 & n1883 ) | ( n1737 & n1883 ) ;
  assign n1911 = n1875 ^ n1770 ^ x88 ;
  assign n1912 = n1870 ^ n1783 ^ x83 ;
  assign n1913 = n1873 ^ n1774 ^ x86 ;
  assign n1914 = n322 | n1724 ;
  assign n1915 = ( n322 & n1910 ) | ( n322 & n1914 ) | ( n1910 & n1914 ) ;
  assign n1916 = n1874 ^ n1792 ^ x87 ;
  assign n1917 = n1885 ^ n1837 ^ 1'b0 ;
  assign n1918 = ( n1837 & n1858 ) | ( n1837 & ~n1917 ) | ( n1858 & ~n1917 ) ;
  assign n1919 = n1868 ^ n1787 ^ x81 ;
  assign n1920 = n1885 ^ n1792 ^ 1'b0 ;
  assign n1921 = n1871 ^ n1780 ^ x84 ;
  assign n1922 = n1869 ^ n1785 ^ x82 ;
  assign n1923 = n1872 ^ n1777 ^ x85 ;
  assign n1924 = n1885 ^ n1810 ^ 1'b0 ;
  assign n1925 = ( n1792 & n1916 ) | ( n1792 & ~n1920 ) | ( n1916 & ~n1920 ) ;
  assign n1926 = n1885 ^ n1787 ^ 1'b0 ;
  assign n1927 = n1885 ^ n1780 ^ 1'b0 ;
  assign n1928 = ( n1780 & n1921 ) | ( n1780 & ~n1927 ) | ( n1921 & ~n1927 ) ;
  assign n1929 = n1885 ^ n1770 ^ 1'b0 ;
  assign n1930 = n1885 ^ n1812 ^ 1'b0 ;
  assign n1931 = ( n1812 & n1859 ) | ( n1812 & ~n1930 ) | ( n1859 & ~n1930 ) ;
  assign n1932 = n1885 ^ n1817 ^ 1'b0 ;
  assign n1933 = n1885 ^ n1774 ^ 1'b0 ;
  assign n1934 = ( n1770 & n1911 ) | ( n1770 & ~n1929 ) | ( n1911 & ~n1929 ) ;
  assign n1935 = n1885 ^ n1777 ^ 1'b0 ;
  assign n1936 = n1885 ^ n1783 ^ 1'b0 ;
  assign n1937 = n1857 ^ n1810 ^ x80 ;
  assign n1938 = n1876 ^ n1767 ^ x89 ;
  assign n1939 = ( n1810 & ~n1924 ) | ( n1810 & n1937 ) | ( ~n1924 & n1937 ) ;
  assign n1940 = n1885 ^ n1767 ^ 1'b0 ;
  assign n1941 = ( n1767 & n1938 ) | ( n1767 & ~n1940 ) | ( n1938 & ~n1940 ) ;
  assign n1942 = ( n1787 & n1919 ) | ( n1787 & ~n1926 ) | ( n1919 & ~n1926 ) ;
  assign n1943 = n1885 ^ n1785 ^ 1'b0 ;
  assign n1944 = ( n1785 & n1922 ) | ( n1785 & ~n1943 ) | ( n1922 & ~n1943 ) ;
  assign n1945 = ( n1774 & n1913 ) | ( n1774 & ~n1933 ) | ( n1913 & ~n1933 ) ;
  assign n1946 = ( n1777 & n1923 ) | ( n1777 & ~n1935 ) | ( n1923 & ~n1935 ) ;
  assign n1947 = ( n1817 & n1860 ) | ( n1817 & ~n1932 ) | ( n1860 & ~n1932 ) ;
  assign n1948 = ( n1783 & n1912 ) | ( n1783 & ~n1936 ) | ( n1912 & ~n1936 ) ;
  assign n1949 = x64 & n1885 ;
  assign n1950 = ~x36 & x64 ;
  assign n1951 = n1949 ^ x64 ^ x37 ;
  assign n1952 = n1951 ^ n1950 ^ x65 ;
  assign n1953 = ( x65 & n1950 ) | ( x65 & n1952 ) | ( n1950 & n1952 ) ;
  assign n1954 = n1953 ^ n1909 ^ x66 ;
  assign n1955 = ~n184 & n1950 ;
  assign n1956 = ( x66 & n1953 ) | ( x66 & n1954 ) | ( n1953 & n1954 ) ;
  assign n1957 = ( x67 & ~n1907 ) | ( x67 & n1956 ) | ( ~n1907 & n1956 ) ;
  assign n1958 = ( x68 & ~n1905 ) | ( x68 & n1957 ) | ( ~n1905 & n1957 ) ;
  assign n1959 = ( x69 & ~n1903 ) | ( x69 & n1958 ) | ( ~n1903 & n1958 ) ;
  assign n1960 = ( x70 & ~n1901 ) | ( x70 & n1959 ) | ( ~n1901 & n1959 ) ;
  assign n1961 = ( x71 & ~n1899 ) | ( x71 & n1960 ) | ( ~n1899 & n1960 ) ;
  assign n1962 = ( x72 & ~n1918 ) | ( x72 & n1961 ) | ( ~n1918 & n1961 ) ;
  assign n1963 = ( x73 & ~n1931 ) | ( x73 & n1962 ) | ( ~n1931 & n1962 ) ;
  assign n1964 = ( x74 & ~n1947 ) | ( x74 & n1963 ) | ( ~n1947 & n1963 ) ;
  assign n1965 = ( x75 & ~n1897 ) | ( x75 & n1964 ) | ( ~n1897 & n1964 ) ;
  assign n1966 = ( x76 & ~n1895 ) | ( x76 & n1965 ) | ( ~n1895 & n1965 ) ;
  assign n1967 = ( x77 & ~n1893 ) | ( x77 & n1966 ) | ( ~n1893 & n1966 ) ;
  assign n1968 = ( x78 & ~n1891 ) | ( x78 & n1967 ) | ( ~n1891 & n1967 ) ;
  assign n1969 = ( x79 & ~n1889 ) | ( x79 & n1968 ) | ( ~n1889 & n1968 ) ;
  assign n1970 = n1969 ^ n1887 ^ x80 ;
  assign n1971 = n1956 ^ n1907 ^ x67 ;
  assign n1972 = ( x80 & ~n1887 ) | ( x80 & n1969 ) | ( ~n1887 & n1969 ) ;
  assign n1973 = ( x81 & ~n1939 ) | ( x81 & n1972 ) | ( ~n1939 & n1972 ) ;
  assign n1974 = n1972 ^ n1939 ^ x81 ;
  assign n1975 = ( x82 & ~n1942 ) | ( x82 & n1973 ) | ( ~n1942 & n1973 ) ;
  assign n1976 = ( x83 & ~n1944 ) | ( x83 & n1975 ) | ( ~n1944 & n1975 ) ;
  assign n1977 = ( x84 & ~n1948 ) | ( x84 & n1976 ) | ( ~n1948 & n1976 ) ;
  assign n1978 = ( x85 & ~n1928 ) | ( x85 & n1977 ) | ( ~n1928 & n1977 ) ;
  assign n1979 = ( x86 & ~n1946 ) | ( x86 & n1978 ) | ( ~n1946 & n1978 ) ;
  assign n1980 = ( x87 & ~n1945 ) | ( x87 & n1979 ) | ( ~n1945 & n1979 ) ;
  assign n1981 = ( x88 & ~n1925 ) | ( x88 & n1980 ) | ( ~n1925 & n1980 ) ;
  assign n1982 = ( x89 & ~n1934 ) | ( x89 & n1981 ) | ( ~n1934 & n1981 ) ;
  assign n1983 = ( x90 & ~n1941 ) | ( x90 & n1982 ) | ( ~n1941 & n1982 ) ;
  assign n1984 = ( x91 & ~n1915 ) | ( x91 & n1983 ) | ( ~n1915 & n1983 ) ;
  assign n1985 = n1520 | n1984 ;
  assign n1986 = n1985 ^ n1887 ^ 1'b0 ;
  assign n1987 = ( n1887 & n1970 ) | ( n1887 & ~n1986 ) | ( n1970 & ~n1986 ) ;
  assign n1988 = n1985 ^ n1939 ^ 1'b0 ;
  assign n1989 = n1985 ^ n1903 ^ 1'b0 ;
  assign n1990 = n1982 ^ n1941 ^ x90 ;
  assign n1991 = ( n1939 & n1974 ) | ( n1939 & ~n1988 ) | ( n1974 & ~n1988 ) ;
  assign n1992 = n1985 ^ n1907 ^ 1'b0 ;
  assign n1993 = ( n1907 & n1971 ) | ( n1907 & ~n1992 ) | ( n1971 & ~n1992 ) ;
  assign n1994 = n1981 ^ n1934 ^ x89 ;
  assign n1995 = n1985 ^ n1891 ^ 1'b0 ;
  assign n1996 = n1985 ^ n1934 ^ 1'b0 ;
  assign n1997 = ( n1934 & n1994 ) | ( n1934 & ~n1996 ) | ( n1994 & ~n1996 ) ;
  assign n1998 = n1967 ^ n1891 ^ x78 ;
  assign n1999 = n1958 ^ n1903 ^ x69 ;
  assign n2000 = ( n1903 & ~n1989 ) | ( n1903 & n1999 ) | ( ~n1989 & n1999 ) ;
  assign n2001 = ( n1891 & ~n1995 ) | ( n1891 & n1998 ) | ( ~n1995 & n1998 ) ;
  assign n2002 = n1990 ^ n1985 ^ 1'b0 ;
  assign n2003 = n1985 ^ n1952 ^ 1'b0 ;
  assign n2004 = ( ~n243 & n1955 ) | ( ~n243 & n1984 ) | ( n1955 & n1984 ) ;
  assign n2005 = ( n1951 & n1952 ) | ( n1951 & n2003 ) | ( n1952 & n2003 ) ;
  assign n2006 = ( n1941 & n1990 ) | ( n1941 & n2002 ) | ( n1990 & n2002 ) ;
  assign n2007 = n1978 ^ n1946 ^ x86 ;
  assign n2008 = ( x36 & n175 ) | ( x36 & n1984 ) | ( n175 & n1984 ) ;
  assign n2009 = ~n1984 & n2004 ;
  assign n2010 = n1985 ^ n1946 ^ 1'b0 ;
  assign n2011 = n1964 ^ n1897 ^ x75 ;
  assign n2012 = ( n1946 & n2007 ) | ( n1946 & ~n2010 ) | ( n2007 & ~n2010 ) ;
  assign n2013 = n1985 ^ n1893 ^ 1'b0 ;
  assign n2014 = n1975 ^ n1944 ^ x83 ;
  assign n2015 = n1980 ^ n1925 ^ x88 ;
  assign n2016 = n1973 ^ n1942 ^ x82 ;
  assign n2017 = n1985 ^ n1925 ^ 1'b0 ;
  assign n2018 = ( n1925 & n2015 ) | ( n1925 & ~n2017 ) | ( n2015 & ~n2017 ) ;
  assign n2019 = n1985 ^ n1947 ^ 1'b0 ;
  assign n2020 = n1961 ^ n1918 ^ x72 ;
  assign n2021 = n1985 ^ n1897 ^ 1'b0 ;
  assign n2022 = n1960 ^ n1899 ^ x71 ;
  assign n2023 = n1966 ^ n1893 ^ x77 ;
  assign n2024 = ( n1893 & ~n2013 ) | ( n1893 & n2023 ) | ( ~n2013 & n2023 ) ;
  assign n2025 = n1957 ^ n1905 ^ x68 ;
  assign n2026 = n1968 ^ n1889 ^ x79 ;
  assign n2027 = n1985 ^ n1889 ^ 1'b0 ;
  assign n2028 = n1985 ^ n1895 ^ 1'b0 ;
  assign n2029 = ( n1889 & n2026 ) | ( n1889 & ~n2027 ) | ( n2026 & ~n2027 ) ;
  assign n2030 = n1962 ^ n1931 ^ x73 ;
  assign n2031 = n1985 ^ n1931 ^ 1'b0 ;
  assign n2032 = n1963 ^ n1947 ^ x74 ;
  assign n2033 = n1985 ^ n1944 ^ 1'b0 ;
  assign n2034 = ( n1944 & n2014 ) | ( n1944 & ~n2033 ) | ( n2014 & ~n2033 ) ;
  assign n2035 = n1985 ^ n1942 ^ 1'b0 ;
  assign n2036 = ( n1942 & n2016 ) | ( n1942 & ~n2035 ) | ( n2016 & ~n2035 ) ;
  assign n2037 = n1979 ^ n1945 ^ x87 ;
  assign n2038 = n1985 ^ n1945 ^ 1'b0 ;
  assign n2039 = ( n1945 & n2037 ) | ( n1945 & ~n2038 ) | ( n2037 & ~n2038 ) ;
  assign n2040 = n1985 ^ n1954 ^ 1'b0 ;
  assign n2041 = n1985 ^ n1905 ^ 1'b0 ;
  assign n2042 = n1985 ^ n1899 ^ 1'b0 ;
  assign n2043 = n1985 ^ n1918 ^ 1'b0 ;
  assign n2044 = n1965 ^ n1895 ^ x76 ;
  assign n2045 = ( n1895 & ~n2028 ) | ( n1895 & n2044 ) | ( ~n2028 & n2044 ) ;
  assign n2046 = n1985 ^ n1948 ^ 1'b0 ;
  assign n2047 = n1976 ^ n1948 ^ x84 ;
  assign n2048 = ( n1897 & n2011 ) | ( n1897 & ~n2021 ) | ( n2011 & ~n2021 ) ;
  assign n2049 = ( n1947 & ~n2019 ) | ( n1947 & n2032 ) | ( ~n2019 & n2032 ) ;
  assign n2050 = ( n1931 & n2030 ) | ( n1931 & ~n2031 ) | ( n2030 & ~n2031 ) ;
  assign n2051 = ( n1918 & n2020 ) | ( n1918 & ~n2043 ) | ( n2020 & ~n2043 ) ;
  assign n2052 = ( n1899 & n2022 ) | ( n1899 & ~n2042 ) | ( n2022 & ~n2042 ) ;
  assign n2053 = ( n1948 & ~n2046 ) | ( n1948 & n2047 ) | ( ~n2046 & n2047 ) ;
  assign n2054 = ( n1905 & n2025 ) | ( n1905 & ~n2041 ) | ( n2025 & ~n2041 ) ;
  assign n2055 = ( n1909 & n1954 ) | ( n1909 & n2040 ) | ( n1954 & n2040 ) ;
  assign n2056 = n1959 ^ n1901 ^ x70 ;
  assign n2057 = n1985 ^ n1901 ^ 1'b0 ;
  assign n2058 = x36 & ~x64 ;
  assign n2059 = ( x36 & x92 ) | ( x36 & n202 ) | ( x92 & n202 ) ;
  assign n2060 = ( x36 & n2008 ) | ( x36 & n2059 ) | ( n2008 & n2059 ) ;
  assign n2061 = n1977 ^ n1928 ^ x85 ;
  assign n2062 = n1985 ^ n1928 ^ 1'b0 ;
  assign n2063 = ( n1901 & n2056 ) | ( n1901 & ~n2057 ) | ( n2056 & ~n2057 ) ;
  assign n2064 = ~x35 & x64 ;
  assign n2065 = ( n322 & n1915 ) | ( n322 & n1985 ) | ( n1915 & n1985 ) ;
  assign n2066 = ( ~x94 & x95 ) | ( ~x94 & n206 ) | ( x95 & n206 ) ;
  assign n2067 = ( x36 & n2058 ) | ( x36 & n2060 ) | ( n2058 & n2060 ) ;
  assign n2068 = n2009 | n2067 ;
  assign n2069 = n2068 ^ n2064 ^ x65 ;
  assign n2070 = ( x65 & n2064 ) | ( x65 & n2069 ) | ( n2064 & n2069 ) ;
  assign n2071 = n2070 ^ n2005 ^ x66 ;
  assign n2072 = ( x66 & n2070 ) | ( x66 & n2071 ) | ( n2070 & n2071 ) ;
  assign n2073 = ( x67 & ~n2055 ) | ( x67 & n2072 ) | ( ~n2055 & n2072 ) ;
  assign n2074 = ( x68 & ~n1993 ) | ( x68 & n2073 ) | ( ~n1993 & n2073 ) ;
  assign n2075 = ( x69 & ~n2054 ) | ( x69 & n2074 ) | ( ~n2054 & n2074 ) ;
  assign n2076 = ( x70 & ~n2000 ) | ( x70 & n2075 ) | ( ~n2000 & n2075 ) ;
  assign n2077 = ( x71 & ~n2063 ) | ( x71 & n2076 ) | ( ~n2063 & n2076 ) ;
  assign n2078 = ( x72 & ~n2052 ) | ( x72 & n2077 ) | ( ~n2052 & n2077 ) ;
  assign n2079 = ( x73 & ~n2051 ) | ( x73 & n2078 ) | ( ~n2051 & n2078 ) ;
  assign n2080 = ( x74 & ~n2050 ) | ( x74 & n2079 ) | ( ~n2050 & n2079 ) ;
  assign n2081 = ( x75 & ~n2049 ) | ( x75 & n2080 ) | ( ~n2049 & n2080 ) ;
  assign n2082 = ( x76 & ~n2048 ) | ( x76 & n2081 ) | ( ~n2048 & n2081 ) ;
  assign n2083 = ( x77 & ~n2045 ) | ( x77 & n2082 ) | ( ~n2045 & n2082 ) ;
  assign n2084 = ( x78 & ~n2024 ) | ( x78 & n2083 ) | ( ~n2024 & n2083 ) ;
  assign n2085 = ( x79 & ~n2001 ) | ( x79 & n2084 ) | ( ~n2001 & n2084 ) ;
  assign n2086 = ( x80 & ~n2029 ) | ( x80 & n2085 ) | ( ~n2029 & n2085 ) ;
  assign n2087 = n2086 ^ n1987 ^ x81 ;
  assign n2088 = n2073 ^ n1993 ^ x68 ;
  assign n2089 = n2072 ^ n2055 ^ x67 ;
  assign n2090 = n2074 ^ n2054 ^ x69 ;
  assign n2091 = n2075 ^ n2000 ^ x70 ;
  assign n2092 = n208 & ~n2066 ;
  assign n2093 = ( x81 & ~n1987 ) | ( x81 & n2086 ) | ( ~n1987 & n2086 ) ;
  assign n2094 = ( n1928 & n2061 ) | ( n1928 & ~n2062 ) | ( n2061 & ~n2062 ) ;
  assign n2095 = ( x82 & ~n1991 ) | ( x82 & n2093 ) | ( ~n1991 & n2093 ) ;
  assign n2096 = ( x83 & ~n2036 ) | ( x83 & n2095 ) | ( ~n2036 & n2095 ) ;
  assign n2097 = ( x84 & ~n2034 ) | ( x84 & n2096 ) | ( ~n2034 & n2096 ) ;
  assign n2098 = ( x85 & ~n2053 ) | ( x85 & n2097 ) | ( ~n2053 & n2097 ) ;
  assign n2099 = ( x86 & ~n2094 ) | ( x86 & n2098 ) | ( ~n2094 & n2098 ) ;
  assign n2100 = ( x87 & ~n2012 ) | ( x87 & n2099 ) | ( ~n2012 & n2099 ) ;
  assign n2101 = ( x88 & ~n2039 ) | ( x88 & n2100 ) | ( ~n2039 & n2100 ) ;
  assign n2102 = ( x89 & ~n2018 ) | ( x89 & n2101 ) | ( ~n2018 & n2101 ) ;
  assign n2103 = ( x90 & ~n1997 ) | ( x90 & n2102 ) | ( ~n1997 & n2102 ) ;
  assign n2104 = ( x91 & ~n2006 ) | ( x91 & n2103 ) | ( ~n2006 & n2103 ) ;
  assign n2105 = ( x92 & ~n2065 ) | ( x92 & n2104 ) | ( ~n2065 & n2104 ) ;
  assign n2106 = n1727 | n2105 ;
  assign n2107 = n2092 & ~n2105 ;
  assign n2108 = n2106 ^ n1987 ^ 1'b0 ;
  assign n2109 = n2098 ^ n2094 ^ x86 ;
  assign n2110 = n2096 ^ n2034 ^ x84 ;
  assign n2111 = n2100 ^ n2039 ^ x88 ;
  assign n2112 = n2064 & ~n2106 ;
  assign n2113 = n2099 ^ n2012 ^ x87 ;
  assign n2114 = n2101 ^ n2018 ^ x89 ;
  assign n2115 = n2097 ^ n2053 ^ x85 ;
  assign n2116 = n2102 ^ n1997 ^ x90 ;
  assign n2117 = ( n1987 & n2087 ) | ( n1987 & ~n2108 ) | ( n2087 & ~n2108 ) ;
  assign n2118 = n2106 ^ n2055 ^ 1'b0 ;
  assign n2119 = ( n2055 & n2089 ) | ( n2055 & ~n2118 ) | ( n2089 & ~n2118 ) ;
  assign n2120 = n2106 ^ n2094 ^ 1'b0 ;
  assign n2121 = n2106 ^ n1997 ^ 1'b0 ;
  assign n2122 = n2106 ^ n2069 ^ 1'b0 ;
  assign n2123 = ( n2094 & n2109 ) | ( n2094 & ~n2120 ) | ( n2109 & ~n2120 ) ;
  assign n2124 = ( n2068 & n2069 ) | ( n2068 & n2122 ) | ( n2069 & n2122 ) ;
  assign n2125 = n2103 ^ n2006 ^ x91 ;
  assign n2126 = n2106 ^ n2053 ^ 1'b0 ;
  assign n2127 = n2106 ^ n2054 ^ 1'b0 ;
  assign n2128 = n2106 ^ n2034 ^ 1'b0 ;
  assign n2129 = ( n2034 & n2110 ) | ( n2034 & ~n2128 ) | ( n2110 & ~n2128 ) ;
  assign n2130 = n2106 ^ n2018 ^ 1'b0 ;
  assign n2131 = ( n2018 & n2114 ) | ( n2018 & ~n2130 ) | ( n2114 & ~n2130 ) ;
  assign n2132 = n2106 ^ n2012 ^ 1'b0 ;
  assign n2133 = ( n2053 & n2115 ) | ( n2053 & ~n2126 ) | ( n2115 & ~n2126 ) ;
  assign n2134 = n2106 ^ n1993 ^ 1'b0 ;
  assign n2135 = n2106 ^ n2000 ^ 1'b0 ;
  assign n2136 = n2106 ^ n2071 ^ 1'b0 ;
  assign n2137 = ( n2005 & n2071 ) | ( n2005 & n2136 ) | ( n2071 & n2136 ) ;
  assign n2138 = n2106 ^ n2039 ^ 1'b0 ;
  assign n2139 = ( n2012 & n2113 ) | ( n2012 & ~n2132 ) | ( n2113 & ~n2132 ) ;
  assign n2140 = n2125 ^ n2106 ^ 1'b0 ;
  assign n2141 = ( n2054 & n2090 ) | ( n2054 & ~n2127 ) | ( n2090 & ~n2127 ) ;
  assign n2142 = ( n2006 & n2125 ) | ( n2006 & n2140 ) | ( n2125 & n2140 ) ;
  assign n2143 = ( n1997 & n2116 ) | ( n1997 & ~n2121 ) | ( n2116 & ~n2121 ) ;
  assign n2144 = ( n2039 & n2111 ) | ( n2039 & ~n2138 ) | ( n2111 & ~n2138 ) ;
  assign n2145 = ( n1993 & n2088 ) | ( n1993 & ~n2134 ) | ( n2088 & ~n2134 ) ;
  assign n2146 = ( n2000 & n2091 ) | ( n2000 & ~n2135 ) | ( n2091 & ~n2135 ) ;
  assign n2147 = n2106 ^ n2048 ^ 1'b0 ;
  assign n2148 = n2084 ^ n2001 ^ x79 ;
  assign n2149 = n2093 ^ n1991 ^ x82 ;
  assign n2150 = n2095 ^ n2036 ^ x83 ;
  assign n2151 = n2106 ^ n1991 ^ 1'b0 ;
  assign n2152 = n2065 & n2106 ;
  assign n2153 = ( n322 & n1727 ) | ( n322 & n2065 ) | ( n1727 & n2065 ) ;
  assign n2154 = n2106 ^ n2001 ^ 1'b0 ;
  assign n2155 = ( n2001 & n2148 ) | ( n2001 & ~n2154 ) | ( n2148 & ~n2154 ) ;
  assign n2156 = n2106 ^ n2036 ^ 1'b0 ;
  assign n2157 = n2083 ^ n2024 ^ x78 ;
  assign n2158 = ~x34 & x64 ;
  assign n2159 = n2081 ^ n2048 ^ x76 ;
  assign n2160 = ( x35 & ~n2107 ) | ( x35 & n2112 ) | ( ~n2107 & n2112 ) ;
  assign n2161 = n2106 ^ n2024 ^ 1'b0 ;
  assign n2162 = ( n1991 & n2149 ) | ( n1991 & ~n2151 ) | ( n2149 & ~n2151 ) ;
  assign n2163 = n2160 ^ n2158 ^ x65 ;
  assign n2164 = ( x65 & n2158 ) | ( x65 & n2163 ) | ( n2158 & n2163 ) ;
  assign n2165 = n2164 ^ n2124 ^ x66 ;
  assign n2166 = ( x66 & n2164 ) | ( x66 & n2165 ) | ( n2164 & n2165 ) ;
  assign n2167 = ( n2036 & n2150 ) | ( n2036 & ~n2156 ) | ( n2150 & ~n2156 ) ;
  assign n2168 = ( x67 & ~n2137 ) | ( x67 & n2166 ) | ( ~n2137 & n2166 ) ;
  assign n2169 = ( x68 & ~n2119 ) | ( x68 & n2168 ) | ( ~n2119 & n2168 ) ;
  assign n2170 = ( n2024 & n2157 ) | ( n2024 & ~n2161 ) | ( n2157 & ~n2161 ) ;
  assign n2171 = n2078 ^ n2051 ^ x73 ;
  assign n2172 = n2169 ^ n2145 ^ x69 ;
  assign n2173 = n2106 ^ n2050 ^ 1'b0 ;
  assign n2174 = n2079 ^ n2050 ^ x74 ;
  assign n2175 = ( n2050 & ~n2173 ) | ( n2050 & n2174 ) | ( ~n2173 & n2174 ) ;
  assign n2176 = n2106 ^ n2063 ^ 1'b0 ;
  assign n2177 = ( x69 & ~n2145 ) | ( x69 & n2169 ) | ( ~n2145 & n2169 ) ;
  assign n2178 = ( n2048 & ~n2147 ) | ( n2048 & n2159 ) | ( ~n2147 & n2159 ) ;
  assign n2179 = ( x70 & ~n2141 ) | ( x70 & n2177 ) | ( ~n2141 & n2177 ) ;
  assign n2180 = n2179 ^ n2146 ^ x71 ;
  assign n2181 = n2106 ^ n2052 ^ 1'b0 ;
  assign n2182 = ( x71 & ~n2146 ) | ( x71 & n2179 ) | ( ~n2146 & n2179 ) ;
  assign n2183 = n2077 ^ n2052 ^ x72 ;
  assign n2184 = ( n2052 & ~n2181 ) | ( n2052 & n2183 ) | ( ~n2181 & n2183 ) ;
  assign n2185 = n2076 ^ n2063 ^ x71 ;
  assign n2186 = ( n2063 & ~n2176 ) | ( n2063 & n2185 ) | ( ~n2176 & n2185 ) ;
  assign n2187 = n2106 ^ n2051 ^ 1'b0 ;
  assign n2188 = n2085 ^ n2029 ^ x80 ;
  assign n2189 = n322 | n2152 ;
  assign n2190 = ( x93 & n199 ) | ( x93 & ~n2152 ) | ( n199 & ~n2152 ) ;
  assign n2191 = ( ~x93 & n199 ) | ( ~x93 & n2189 ) | ( n199 & n2189 ) ;
  assign n2192 = ( n2051 & n2171 ) | ( n2051 & ~n2187 ) | ( n2171 & ~n2187 ) ;
  assign n2193 = ( x72 & n2182 ) | ( x72 & ~n2186 ) | ( n2182 & ~n2186 ) ;
  assign n2194 = n2106 ^ n2029 ^ 1'b0 ;
  assign n2195 = n2106 ^ n2045 ^ 1'b0 ;
  assign n2196 = ( n2029 & n2188 ) | ( n2029 & ~n2194 ) | ( n2188 & ~n2194 ) ;
  assign n2197 = n2080 ^ n2049 ^ x75 ;
  assign n2198 = n2177 ^ n2141 ^ x70 ;
  assign n2199 = n2106 ^ n2049 ^ 1'b0 ;
  assign n2200 = x94 | n2066 ;
  assign n2201 = ( x73 & ~n2184 ) | ( x73 & n2193 ) | ( ~n2184 & n2193 ) ;
  assign n2202 = n2168 ^ n2119 ^ x68 ;
  assign n2203 = n2166 ^ n2137 ^ x67 ;
  assign n2204 = ( n2190 & n2191 ) | ( n2190 & ~n2200 ) | ( n2191 & ~n2200 ) ;
  assign n2205 = n2082 ^ n2045 ^ x77 ;
  assign n2206 = ( n2049 & n2197 ) | ( n2049 & ~n2199 ) | ( n2197 & ~n2199 ) ;
  assign n2207 = ( n2045 & ~n2195 ) | ( n2045 & n2205 ) | ( ~n2195 & n2205 ) ;
  assign n2208 = n2201 ^ n2192 ^ x74 ;
  assign n2209 = ( x74 & ~n2192 ) | ( x74 & n2201 ) | ( ~n2192 & n2201 ) ;
  assign n2210 = ( x75 & ~n2175 ) | ( x75 & n2209 ) | ( ~n2175 & n2209 ) ;
  assign n2211 = ( x76 & ~n2206 ) | ( x76 & n2210 ) | ( ~n2206 & n2210 ) ;
  assign n2212 = ( x77 & ~n2178 ) | ( x77 & n2211 ) | ( ~n2178 & n2211 ) ;
  assign n2213 = n2186 ^ n2182 ^ x72 ;
  assign n2214 = ( x78 & ~n2207 ) | ( x78 & n2212 ) | ( ~n2207 & n2212 ) ;
  assign n2215 = n2193 ^ n2184 ^ x73 ;
  assign n2216 = n2209 ^ n2175 ^ x75 ;
  assign n2217 = n2210 ^ n2206 ^ x76 ;
  assign n2218 = n2211 ^ n2178 ^ x77 ;
  assign n2219 = n2212 ^ n2207 ^ x78 ;
  assign n2220 = n1727 & n2189 ;
  assign n2221 = ( x79 & ~n2170 ) | ( x79 & n2214 ) | ( ~n2170 & n2214 ) ;
  assign n2222 = ( x80 & ~n2155 ) | ( x80 & n2221 ) | ( ~n2155 & n2221 ) ;
  assign n2223 = ( x81 & ~n2196 ) | ( x81 & n2222 ) | ( ~n2196 & n2222 ) ;
  assign n2224 = ( x82 & ~n2117 ) | ( x82 & n2223 ) | ( ~n2117 & n2223 ) ;
  assign n2225 = ( x83 & ~n2162 ) | ( x83 & n2224 ) | ( ~n2162 & n2224 ) ;
  assign n2226 = ( x84 & ~n2167 ) | ( x84 & n2225 ) | ( ~n2167 & n2225 ) ;
  assign n2227 = ( x85 & ~n2129 ) | ( x85 & n2226 ) | ( ~n2129 & n2226 ) ;
  assign n2228 = ( x86 & ~n2133 ) | ( x86 & n2227 ) | ( ~n2133 & n2227 ) ;
  assign n2229 = ( x87 & ~n2123 ) | ( x87 & n2228 ) | ( ~n2123 & n2228 ) ;
  assign n2230 = ( x88 & ~n2139 ) | ( x88 & n2229 ) | ( ~n2139 & n2229 ) ;
  assign n2231 = ( x89 & ~n2144 ) | ( x89 & n2230 ) | ( ~n2144 & n2230 ) ;
  assign n2232 = ( x90 & ~n2131 ) | ( x90 & n2231 ) | ( ~n2131 & n2231 ) ;
  assign n2233 = ( x91 & ~n2143 ) | ( x91 & n2232 ) | ( ~n2143 & n2232 ) ;
  assign n2234 = ( x92 & ~n2142 ) | ( x92 & n2233 ) | ( ~n2142 & n2233 ) ;
  assign n2235 = ( ~n2200 & n2204 ) | ( ~n2200 & n2234 ) | ( n2204 & n2234 ) ;
  assign n2236 = n2200 | n2235 ;
  assign n2237 = ( ~n2189 & n2220 ) | ( ~n2189 & n2236 ) | ( n2220 & n2236 ) ;
  assign n2238 = n2237 ^ n2207 ^ 1'b0 ;
  assign n2239 = ( n2207 & n2219 ) | ( n2207 & ~n2238 ) | ( n2219 & ~n2238 ) ;
  assign n2240 = n2237 ^ n2178 ^ 1'b0 ;
  assign n2241 = ( n2178 & n2218 ) | ( n2178 & ~n2240 ) | ( n2218 & ~n2240 ) ;
  assign n2242 = n2237 ^ n2206 ^ 1'b0 ;
  assign n2243 = ( n2206 & n2217 ) | ( n2206 & ~n2242 ) | ( n2217 & ~n2242 ) ;
  assign n2244 = n2237 ^ n2175 ^ 1'b0 ;
  assign n2245 = ( n2175 & n2216 ) | ( n2175 & ~n2244 ) | ( n2216 & ~n2244 ) ;
  assign n2246 = n2237 ^ n2192 ^ 1'b0 ;
  assign n2247 = ( n2192 & n2208 ) | ( n2192 & ~n2246 ) | ( n2208 & ~n2246 ) ;
  assign n2248 = n2237 ^ n2184 ^ 1'b0 ;
  assign n2249 = ( n2184 & n2215 ) | ( n2184 & ~n2248 ) | ( n2215 & ~n2248 ) ;
  assign n2250 = n2237 ^ n2186 ^ 1'b0 ;
  assign n2251 = ( n2186 & n2213 ) | ( n2186 & ~n2250 ) | ( n2213 & ~n2250 ) ;
  assign n2252 = n2237 ^ n2146 ^ 1'b0 ;
  assign n2253 = ( n2146 & n2180 ) | ( n2146 & ~n2252 ) | ( n2180 & ~n2252 ) ;
  assign n2254 = n2237 ^ n2141 ^ 1'b0 ;
  assign n2255 = ( n2141 & n2198 ) | ( n2141 & ~n2254 ) | ( n2198 & ~n2254 ) ;
  assign n2256 = n2237 ^ n2145 ^ 1'b0 ;
  assign n2257 = ( n2145 & n2172 ) | ( n2145 & ~n2256 ) | ( n2172 & ~n2256 ) ;
  assign n2258 = n2237 ^ n2119 ^ 1'b0 ;
  assign n2259 = ( n2119 & n2202 ) | ( n2119 & ~n2258 ) | ( n2202 & ~n2258 ) ;
  assign n2260 = n2237 ^ n2137 ^ 1'b0 ;
  assign n2261 = ( n2137 & n2203 ) | ( n2137 & ~n2260 ) | ( n2203 & ~n2260 ) ;
  assign n2262 = n2237 ^ n2165 ^ 1'b0 ;
  assign n2263 = ( n2124 & n2165 ) | ( n2124 & n2262 ) | ( n2165 & n2262 ) ;
  assign n2264 = n2237 ^ n2163 ^ 1'b0 ;
  assign n2265 = ( n2160 & n2163 ) | ( n2160 & n2264 ) | ( n2163 & n2264 ) ;
  assign n2266 = n322 | n2236 ;
  assign n2267 = ( n322 & n2153 ) | ( n322 & n2266 ) | ( n2153 & n2266 ) ;
  assign n2268 = n2233 ^ n2142 ^ x92 ;
  assign n2269 = n2237 ^ n2142 ^ 1'b0 ;
  assign n2270 = ( n2142 & n2268 ) | ( n2142 & ~n2269 ) | ( n2268 & ~n2269 ) ;
  assign n2271 = n2232 ^ n2143 ^ x91 ;
  assign n2272 = n2237 ^ n2143 ^ 1'b0 ;
  assign n2273 = ( n2143 & n2271 ) | ( n2143 & ~n2272 ) | ( n2271 & ~n2272 ) ;
  assign n2274 = n2231 ^ n2131 ^ x90 ;
  assign n2275 = n2237 ^ n2131 ^ 1'b0 ;
  assign n2276 = ( n2131 & n2274 ) | ( n2131 & ~n2275 ) | ( n2274 & ~n2275 ) ;
  assign n2277 = n2230 ^ n2144 ^ x89 ;
  assign n2278 = n2237 ^ n2144 ^ 1'b0 ;
  assign n2279 = ( n2144 & n2277 ) | ( n2144 & ~n2278 ) | ( n2277 & ~n2278 ) ;
  assign n2280 = n2229 ^ n2139 ^ x88 ;
  assign n2281 = n2237 ^ n2139 ^ 1'b0 ;
  assign n2282 = ( n2139 & n2280 ) | ( n2139 & ~n2281 ) | ( n2280 & ~n2281 ) ;
  assign n2283 = n2228 ^ n2123 ^ x87 ;
  assign n2284 = n2237 ^ n2123 ^ 1'b0 ;
  assign n2285 = ( n2123 & n2283 ) | ( n2123 & ~n2284 ) | ( n2283 & ~n2284 ) ;
  assign n2286 = n2227 ^ n2133 ^ x86 ;
  assign n2287 = n2237 ^ n2133 ^ 1'b0 ;
  assign n2288 = ( n2133 & n2286 ) | ( n2133 & ~n2287 ) | ( n2286 & ~n2287 ) ;
  assign n2289 = n2226 ^ n2129 ^ x85 ;
  assign n2290 = n2237 ^ n2129 ^ 1'b0 ;
  assign n2291 = ( n2129 & n2289 ) | ( n2129 & ~n2290 ) | ( n2289 & ~n2290 ) ;
  assign n2292 = n2225 ^ n2167 ^ x84 ;
  assign n2293 = n2237 ^ n2167 ^ 1'b0 ;
  assign n2294 = ( n2167 & n2292 ) | ( n2167 & ~n2293 ) | ( n2292 & ~n2293 ) ;
  assign n2295 = n2224 ^ n2162 ^ x83 ;
  assign n2296 = n2237 ^ n2162 ^ 1'b0 ;
  assign n2297 = ( n2162 & n2295 ) | ( n2162 & ~n2296 ) | ( n2295 & ~n2296 ) ;
  assign n2298 = n2223 ^ n2117 ^ x82 ;
  assign n2299 = n2237 ^ n2117 ^ 1'b0 ;
  assign n2300 = ( n2117 & n2298 ) | ( n2117 & ~n2299 ) | ( n2298 & ~n2299 ) ;
  assign n2301 = n2222 ^ n2196 ^ x81 ;
  assign n2302 = n2237 ^ n2196 ^ 1'b0 ;
  assign n2303 = ( n2196 & n2301 ) | ( n2196 & ~n2302 ) | ( n2301 & ~n2302 ) ;
  assign n2304 = n2221 ^ n2155 ^ x80 ;
  assign n2305 = n2237 ^ n2155 ^ 1'b0 ;
  assign n2306 = ( n2155 & n2304 ) | ( n2155 & ~n2305 ) | ( n2304 & ~n2305 ) ;
  assign n2307 = n2214 ^ n2170 ^ x79 ;
  assign n2308 = n2237 ^ n2170 ^ 1'b0 ;
  assign n2309 = ( n2170 & n2307 ) | ( n2170 & ~n2308 ) | ( n2307 & ~n2308 ) ;
  assign n2310 = ~x33 & x64 ;
  assign n2311 = x64 & n2237 ;
  assign n2312 = n2311 ^ x64 ^ x34 ;
  assign n2313 = n2312 ^ n2310 ^ x65 ;
  assign n2314 = ( x65 & n2310 ) | ( x65 & n2313 ) | ( n2310 & n2313 ) ;
  assign n2315 = n2314 ^ n2265 ^ x66 ;
  assign n2316 = ( x66 & n2314 ) | ( x66 & n2315 ) | ( n2314 & n2315 ) ;
  assign n2317 = ( x67 & ~n2263 ) | ( x67 & n2316 ) | ( ~n2263 & n2316 ) ;
  assign n2318 = ( x68 & ~n2261 ) | ( x68 & n2317 ) | ( ~n2261 & n2317 ) ;
  assign n2319 = ( x69 & ~n2259 ) | ( x69 & n2318 ) | ( ~n2259 & n2318 ) ;
  assign n2320 = ( x70 & ~n2257 ) | ( x70 & n2319 ) | ( ~n2257 & n2319 ) ;
  assign n2321 = ( x71 & ~n2255 ) | ( x71 & n2320 ) | ( ~n2255 & n2320 ) ;
  assign n2322 = ( x72 & ~n2253 ) | ( x72 & n2321 ) | ( ~n2253 & n2321 ) ;
  assign n2323 = ( x73 & ~n2251 ) | ( x73 & n2322 ) | ( ~n2251 & n2322 ) ;
  assign n2324 = ( x74 & ~n2249 ) | ( x74 & n2323 ) | ( ~n2249 & n2323 ) ;
  assign n2325 = ( x75 & ~n2247 ) | ( x75 & n2324 ) | ( ~n2247 & n2324 ) ;
  assign n2326 = ( x76 & ~n2245 ) | ( x76 & n2325 ) | ( ~n2245 & n2325 ) ;
  assign n2327 = ( x77 & ~n2243 ) | ( x77 & n2326 ) | ( ~n2243 & n2326 ) ;
  assign n2328 = ( x78 & ~n2241 ) | ( x78 & n2327 ) | ( ~n2241 & n2327 ) ;
  assign n2329 = ( x79 & ~n2239 ) | ( x79 & n2328 ) | ( ~n2239 & n2328 ) ;
  assign n2330 = ( x80 & ~n2309 ) | ( x80 & n2329 ) | ( ~n2309 & n2329 ) ;
  assign n2331 = ( x81 & ~n2306 ) | ( x81 & n2330 ) | ( ~n2306 & n2330 ) ;
  assign n2332 = ( x82 & ~n2303 ) | ( x82 & n2331 ) | ( ~n2303 & n2331 ) ;
  assign n2333 = ( x83 & ~n2300 ) | ( x83 & n2332 ) | ( ~n2300 & n2332 ) ;
  assign n2334 = ( x84 & ~n2297 ) | ( x84 & n2333 ) | ( ~n2297 & n2333 ) ;
  assign n2335 = ( x85 & ~n2294 ) | ( x85 & n2334 ) | ( ~n2294 & n2334 ) ;
  assign n2336 = ( x86 & ~n2291 ) | ( x86 & n2335 ) | ( ~n2291 & n2335 ) ;
  assign n2337 = ( x87 & ~n2288 ) | ( x87 & n2336 ) | ( ~n2288 & n2336 ) ;
  assign n2338 = ( x88 & ~n2285 ) | ( x88 & n2337 ) | ( ~n2285 & n2337 ) ;
  assign n2339 = ( x89 & ~n2282 ) | ( x89 & n2338 ) | ( ~n2282 & n2338 ) ;
  assign n2340 = ( x90 & ~n2279 ) | ( x90 & n2339 ) | ( ~n2279 & n2339 ) ;
  assign n2341 = ( x91 & ~n2276 ) | ( x91 & n2340 ) | ( ~n2276 & n2340 ) ;
  assign n2342 = ( x92 & ~n2273 ) | ( x92 & n2341 ) | ( ~n2273 & n2341 ) ;
  assign n2343 = ( x93 & ~n2270 ) | ( x93 & n2342 ) | ( ~n2270 & n2342 ) ;
  assign n2344 = ( x94 & ~n2267 ) | ( x94 & n2343 ) | ( ~n2267 & n2343 ) ;
  assign n2345 = n1310 | n2344 ;
  assign n2346 = n2333 ^ n2297 ^ x84 ;
  assign n2347 = n2345 ^ n2297 ^ 1'b0 ;
  assign n2348 = ( n2297 & n2346 ) | ( n2297 & ~n2347 ) | ( n2346 & ~n2347 ) ;
  assign n2349 = n2329 ^ n2309 ^ x80 ;
  assign n2350 = n2345 ^ n2309 ^ 1'b0 ;
  assign n2351 = ( n2309 & n2349 ) | ( n2309 & ~n2350 ) | ( n2349 & ~n2350 ) ;
  assign n2352 = n2327 ^ n2241 ^ x78 ;
  assign n2353 = n2345 ^ n2241 ^ 1'b0 ;
  assign n2354 = ( n2241 & n2352 ) | ( n2241 & ~n2353 ) | ( n2352 & ~n2353 ) ;
  assign n2355 = n2326 ^ n2243 ^ x77 ;
  assign n2356 = n2345 ^ n2243 ^ 1'b0 ;
  assign n2357 = ( n2243 & n2355 ) | ( n2243 & ~n2356 ) | ( n2355 & ~n2356 ) ;
  assign n2358 = n2322 ^ n2251 ^ x73 ;
  assign n2359 = n2345 ^ n2251 ^ 1'b0 ;
  assign n2360 = ( n2251 & n2358 ) | ( n2251 & ~n2359 ) | ( n2358 & ~n2359 ) ;
  assign n2361 = n2320 ^ n2255 ^ x71 ;
  assign n2362 = n2345 ^ n2255 ^ 1'b0 ;
  assign n2363 = ( n2255 & n2361 ) | ( n2255 & ~n2362 ) | ( n2361 & ~n2362 ) ;
  assign n2364 = n2317 ^ n2261 ^ x68 ;
  assign n2365 = n2345 ^ n2261 ^ 1'b0 ;
  assign n2366 = ( n2261 & n2364 ) | ( n2261 & ~n2365 ) | ( n2364 & ~n2365 ) ;
  assign n2367 = n2316 ^ n2263 ^ x67 ;
  assign n2368 = n2345 ^ n2263 ^ 1'b0 ;
  assign n2369 = ( n2263 & n2367 ) | ( n2263 & ~n2368 ) | ( n2367 & ~n2368 ) ;
  assign n2370 = n2345 ^ n2315 ^ 1'b0 ;
  assign n2371 = ( n2265 & n2315 ) | ( n2265 & n2370 ) | ( n2315 & n2370 ) ;
  assign n2372 = n2345 ^ n2313 ^ 1'b0 ;
  assign n2373 = ( n2312 & n2313 ) | ( n2312 & n2372 ) | ( n2313 & n2372 ) ;
  assign n2374 = n2342 ^ n2270 ^ x93 ;
  assign n2375 = n2374 ^ n2345 ^ 1'b0 ;
  assign n2376 = ( n2270 & n2374 ) | ( n2270 & n2375 ) | ( n2374 & n2375 ) ;
  assign n2377 = n2341 ^ n2273 ^ x92 ;
  assign n2378 = n2345 ^ n2273 ^ 1'b0 ;
  assign n2379 = ( n2273 & n2377 ) | ( n2273 & ~n2378 ) | ( n2377 & ~n2378 ) ;
  assign n2380 = n2340 ^ n2276 ^ x91 ;
  assign n2381 = n2345 ^ n2276 ^ 1'b0 ;
  assign n2382 = ( n2276 & n2380 ) | ( n2276 & ~n2381 ) | ( n2380 & ~n2381 ) ;
  assign n2383 = n2339 ^ n2279 ^ x90 ;
  assign n2384 = n2345 ^ n2279 ^ 1'b0 ;
  assign n2385 = ( n2279 & n2383 ) | ( n2279 & ~n2384 ) | ( n2383 & ~n2384 ) ;
  assign n2386 = n2338 ^ n2282 ^ x89 ;
  assign n2387 = n2345 ^ n2282 ^ 1'b0 ;
  assign n2388 = ( n2282 & n2386 ) | ( n2282 & ~n2387 ) | ( n2386 & ~n2387 ) ;
  assign n2389 = n2337 ^ n2285 ^ x88 ;
  assign n2390 = n2345 ^ n2285 ^ 1'b0 ;
  assign n2391 = ( n2285 & n2389 ) | ( n2285 & ~n2390 ) | ( n2389 & ~n2390 ) ;
  assign n2392 = n2336 ^ n2288 ^ x87 ;
  assign n2393 = n2345 ^ n2288 ^ 1'b0 ;
  assign n2394 = ( n2288 & n2392 ) | ( n2288 & ~n2393 ) | ( n2392 & ~n2393 ) ;
  assign n2395 = n2335 ^ n2291 ^ x86 ;
  assign n2396 = n2345 ^ n2291 ^ 1'b0 ;
  assign n2397 = ( n2291 & n2395 ) | ( n2291 & ~n2396 ) | ( n2395 & ~n2396 ) ;
  assign n2398 = n2334 ^ n2294 ^ x85 ;
  assign n2399 = n2345 ^ n2294 ^ 1'b0 ;
  assign n2400 = ( n2294 & n2398 ) | ( n2294 & ~n2399 ) | ( n2398 & ~n2399 ) ;
  assign n2401 = n2332 ^ n2300 ^ x83 ;
  assign n2402 = n2345 ^ n2300 ^ 1'b0 ;
  assign n2403 = ( n2300 & n2401 ) | ( n2300 & ~n2402 ) | ( n2401 & ~n2402 ) ;
  assign n2404 = n2331 ^ n2303 ^ x82 ;
  assign n2405 = n2345 ^ n2303 ^ 1'b0 ;
  assign n2406 = ( n2303 & n2404 ) | ( n2303 & ~n2405 ) | ( n2404 & ~n2405 ) ;
  assign n2407 = n2330 ^ n2306 ^ x81 ;
  assign n2408 = n2345 ^ n2306 ^ 1'b0 ;
  assign n2409 = ( n2306 & n2407 ) | ( n2306 & ~n2408 ) | ( n2407 & ~n2408 ) ;
  assign n2410 = n2328 ^ n2239 ^ x79 ;
  assign n2411 = n2345 ^ n2239 ^ 1'b0 ;
  assign n2412 = ( n2239 & n2410 ) | ( n2239 & ~n2411 ) | ( n2410 & ~n2411 ) ;
  assign n2413 = n2325 ^ n2245 ^ x76 ;
  assign n2414 = n2345 ^ n2245 ^ 1'b0 ;
  assign n2415 = ( n2245 & n2413 ) | ( n2245 & ~n2414 ) | ( n2413 & ~n2414 ) ;
  assign n2416 = n2323 ^ n2249 ^ x74 ;
  assign n2417 = n2345 ^ n2249 ^ 1'b0 ;
  assign n2418 = ( n2249 & n2416 ) | ( n2249 & ~n2417 ) | ( n2416 & ~n2417 ) ;
  assign n2419 = n2321 ^ n2253 ^ x72 ;
  assign n2420 = n2345 ^ n2253 ^ 1'b0 ;
  assign n2421 = ( n2253 & n2419 ) | ( n2253 & ~n2420 ) | ( n2419 & ~n2420 ) ;
  assign n2422 = n2319 ^ n2257 ^ x70 ;
  assign n2423 = n2345 ^ n2257 ^ 1'b0 ;
  assign n2424 = ( n2257 & n2422 ) | ( n2257 & ~n2423 ) | ( n2422 & ~n2423 ) ;
  assign n2425 = n2318 ^ n2259 ^ x69 ;
  assign n2426 = n2345 ^ n2259 ^ 1'b0 ;
  assign n2427 = ( n2259 & n2425 ) | ( n2259 & ~n2426 ) | ( n2425 & ~n2426 ) ;
  assign n2428 = n2310 & ~n2345 ;
  assign n2429 = ~x32 & x64 ;
  assign n2430 = ( ~x33 & x64 ) | ( ~x33 & n2344 ) | ( x64 & n2344 ) ;
  assign n2431 = x64 & ~n2430 ;
  assign n2432 = ( ~x95 & n243 ) | ( ~x95 & n2431 ) | ( n243 & n2431 ) ;
  assign n2433 = ~n243 & n2432 ;
  assign n2434 = ( x33 & n2428 ) | ( x33 & ~n2433 ) | ( n2428 & ~n2433 ) ;
  assign n2435 = n2345 ^ n2247 ^ 1'b0 ;
  assign n2436 = n2434 ^ n2429 ^ x65 ;
  assign n2437 = ( x65 & n2429 ) | ( x65 & n2436 ) | ( n2429 & n2436 ) ;
  assign n2438 = n2437 ^ n2373 ^ x66 ;
  assign n2439 = ( x66 & n2437 ) | ( x66 & n2438 ) | ( n2437 & n2438 ) ;
  assign n2440 = ( x67 & ~n2371 ) | ( x67 & n2439 ) | ( ~n2371 & n2439 ) ;
  assign n2441 = ( x68 & ~n2369 ) | ( x68 & n2440 ) | ( ~n2369 & n2440 ) ;
  assign n2442 = ( x69 & ~n2366 ) | ( x69 & n2441 ) | ( ~n2366 & n2441 ) ;
  assign n2443 = ( x70 & ~n2427 ) | ( x70 & n2442 ) | ( ~n2427 & n2442 ) ;
  assign n2444 = n2324 ^ n2247 ^ x75 ;
  assign n2445 = ( n2247 & ~n2435 ) | ( n2247 & n2444 ) | ( ~n2435 & n2444 ) ;
  assign n2446 = n2440 ^ n2369 ^ x68 ;
  assign n2447 = ( x71 & ~n2424 ) | ( x71 & n2443 ) | ( ~n2424 & n2443 ) ;
  assign n2448 = ( x72 & ~n2363 ) | ( x72 & n2447 ) | ( ~n2363 & n2447 ) ;
  assign n2449 = ( x73 & ~n2421 ) | ( x73 & n2448 ) | ( ~n2421 & n2448 ) ;
  assign n2450 = ( x74 & ~n2360 ) | ( x74 & n2449 ) | ( ~n2360 & n2449 ) ;
  assign n2451 = ( x75 & ~n2418 ) | ( x75 & n2450 ) | ( ~n2418 & n2450 ) ;
  assign n2452 = ( x76 & ~n2445 ) | ( x76 & n2451 ) | ( ~n2445 & n2451 ) ;
  assign n2453 = ( x77 & ~n2415 ) | ( x77 & n2452 ) | ( ~n2415 & n2452 ) ;
  assign n2454 = ( x78 & ~n2357 ) | ( x78 & n2453 ) | ( ~n2357 & n2453 ) ;
  assign n2455 = ( x79 & ~n2354 ) | ( x79 & n2454 ) | ( ~n2354 & n2454 ) ;
  assign n2456 = ( x80 & ~n2412 ) | ( x80 & n2455 ) | ( ~n2412 & n2455 ) ;
  assign n2457 = ( x81 & ~n2351 ) | ( x81 & n2456 ) | ( ~n2351 & n2456 ) ;
  assign n2458 = n2448 ^ n2421 ^ x73 ;
  assign n2459 = n2449 ^ n2360 ^ x74 ;
  assign n2460 = n2457 ^ n2409 ^ x82 ;
  assign n2461 = ( x82 & ~n2409 ) | ( x82 & n2457 ) | ( ~n2409 & n2457 ) ;
  assign n2462 = ( x83 & ~n2406 ) | ( x83 & n2461 ) | ( ~n2406 & n2461 ) ;
  assign n2463 = ( x84 & ~n2403 ) | ( x84 & n2462 ) | ( ~n2403 & n2462 ) ;
  assign n2464 = ( x85 & ~n2348 ) | ( x85 & n2463 ) | ( ~n2348 & n2463 ) ;
  assign n2465 = n2463 ^ n2348 ^ x85 ;
  assign n2466 = n2442 ^ n2427 ^ x70 ;
  assign n2467 = n2447 ^ n2363 ^ x72 ;
  assign n2468 = n2451 ^ n2445 ^ x76 ;
  assign n2469 = ( n322 & n2267 ) | ( n322 & n2345 ) | ( n2267 & n2345 ) ;
  assign n2470 = n2453 ^ n2357 ^ x78 ;
  assign n2471 = n2452 ^ n2415 ^ x77 ;
  assign n2472 = ( x86 & ~n2400 ) | ( x86 & n2464 ) | ( ~n2400 & n2464 ) ;
  assign n2473 = ( x87 & ~n2397 ) | ( x87 & n2472 ) | ( ~n2397 & n2472 ) ;
  assign n2474 = ( x88 & ~n2394 ) | ( x88 & n2473 ) | ( ~n2394 & n2473 ) ;
  assign n2475 = ( x89 & ~n2391 ) | ( x89 & n2474 ) | ( ~n2391 & n2474 ) ;
  assign n2476 = ( x90 & ~n2388 ) | ( x90 & n2475 ) | ( ~n2388 & n2475 ) ;
  assign n2477 = ( x91 & ~n2385 ) | ( x91 & n2476 ) | ( ~n2385 & n2476 ) ;
  assign n2478 = ( x92 & ~n2382 ) | ( x92 & n2477 ) | ( ~n2382 & n2477 ) ;
  assign n2479 = ( x93 & ~n2379 ) | ( x93 & n2478 ) | ( ~n2379 & n2478 ) ;
  assign n2480 = ( x94 & ~n2376 ) | ( x94 & n2479 ) | ( ~n2376 & n2479 ) ;
  assign n2481 = ( x95 & ~n2469 ) | ( x95 & n2480 ) | ( ~n2469 & n2480 ) ;
  assign n2482 = n243 | n2481 ;
  assign n2483 = n2477 ^ n2382 ^ x92 ;
  assign n2484 = n2482 ^ n2382 ^ 1'b0 ;
  assign n2485 = ( n2382 & n2483 ) | ( n2382 & ~n2484 ) | ( n2483 & ~n2484 ) ;
  assign n2486 = n2476 ^ n2385 ^ x91 ;
  assign n2487 = n2482 ^ n2385 ^ 1'b0 ;
  assign n2488 = ( n2385 & n2486 ) | ( n2385 & ~n2487 ) | ( n2486 & ~n2487 ) ;
  assign n2489 = n2475 ^ n2388 ^ x90 ;
  assign n2490 = n2482 ^ n2388 ^ 1'b0 ;
  assign n2491 = ( n2388 & n2489 ) | ( n2388 & ~n2490 ) | ( n2489 & ~n2490 ) ;
  assign n2492 = n2474 ^ n2391 ^ x89 ;
  assign n2493 = n2482 ^ n2391 ^ 1'b0 ;
  assign n2494 = ( n2391 & n2492 ) | ( n2391 & ~n2493 ) | ( n2492 & ~n2493 ) ;
  assign n2495 = n2473 ^ n2394 ^ x88 ;
  assign n2496 = n2482 ^ n2394 ^ 1'b0 ;
  assign n2497 = ( n2394 & n2495 ) | ( n2394 & ~n2496 ) | ( n2495 & ~n2496 ) ;
  assign n2498 = n2482 ^ n2348 ^ 1'b0 ;
  assign n2499 = ( n2348 & n2465 ) | ( n2348 & ~n2498 ) | ( n2465 & ~n2498 ) ;
  assign n2500 = n2462 ^ n2403 ^ x84 ;
  assign n2501 = n2482 ^ n2403 ^ 1'b0 ;
  assign n2502 = n2482 ^ n2409 ^ 1'b0 ;
  assign n2503 = ( n2409 & n2460 ) | ( n2409 & ~n2502 ) | ( n2460 & ~n2502 ) ;
  assign n2504 = n2482 ^ n2357 ^ 1'b0 ;
  assign n2505 = ( n2357 & n2470 ) | ( n2357 & ~n2504 ) | ( n2470 & ~n2504 ) ;
  assign n2506 = n2482 ^ n2415 ^ 1'b0 ;
  assign n2507 = ( n2415 & n2471 ) | ( n2415 & ~n2506 ) | ( n2471 & ~n2506 ) ;
  assign n2508 = n2482 ^ n2445 ^ 1'b0 ;
  assign n2509 = ( n2445 & n2468 ) | ( n2445 & ~n2508 ) | ( n2468 & ~n2508 ) ;
  assign n2510 = ( n2403 & n2500 ) | ( n2403 & ~n2501 ) | ( n2500 & ~n2501 ) ;
  assign n2511 = n2482 ^ n2360 ^ 1'b0 ;
  assign n2512 = ( n2360 & n2459 ) | ( n2360 & ~n2511 ) | ( n2459 & ~n2511 ) ;
  assign n2513 = n2482 ^ n2421 ^ 1'b0 ;
  assign n2514 = ( n2421 & n2458 ) | ( n2421 & ~n2513 ) | ( n2458 & ~n2513 ) ;
  assign n2515 = n2482 ^ n2363 ^ 1'b0 ;
  assign n2516 = ( n2363 & n2467 ) | ( n2363 & ~n2515 ) | ( n2467 & ~n2515 ) ;
  assign n2517 = n2482 ^ n2427 ^ 1'b0 ;
  assign n2518 = ( n2427 & n2466 ) | ( n2427 & ~n2517 ) | ( n2466 & ~n2517 ) ;
  assign n2519 = n2482 ^ n2369 ^ 1'b0 ;
  assign n2520 = ( n2369 & n2446 ) | ( n2369 & ~n2519 ) | ( n2446 & ~n2519 ) ;
  assign n2521 = n2482 ^ n2438 ^ 1'b0 ;
  assign n2522 = ( n2373 & n2438 ) | ( n2373 & n2521 ) | ( n2438 & n2521 ) ;
  assign n2523 = n2482 ^ n2436 ^ 1'b0 ;
  assign n2524 = ( n2434 & n2436 ) | ( n2434 & n2523 ) | ( n2436 & n2523 ) ;
  assign n2525 = n2479 ^ n2376 ^ x94 ;
  assign n2526 = n2482 ^ n2376 ^ 1'b0 ;
  assign n2527 = ( n2376 & n2525 ) | ( n2376 & ~n2526 ) | ( n2525 & ~n2526 ) ;
  assign n2528 = n2478 ^ n2379 ^ x93 ;
  assign n2529 = n2482 ^ n2379 ^ 1'b0 ;
  assign n2530 = ( n2379 & n2528 ) | ( n2379 & ~n2529 ) | ( n2528 & ~n2529 ) ;
  assign n2531 = n2472 ^ n2397 ^ x87 ;
  assign n2532 = n2482 ^ n2397 ^ 1'b0 ;
  assign n2533 = ( n2397 & n2531 ) | ( n2397 & ~n2532 ) | ( n2531 & ~n2532 ) ;
  assign n2534 = n2464 ^ n2400 ^ x86 ;
  assign n2535 = n2482 ^ n2400 ^ 1'b0 ;
  assign n2536 = ( n2400 & n2534 ) | ( n2400 & ~n2535 ) | ( n2534 & ~n2535 ) ;
  assign n2537 = n2461 ^ n2406 ^ x83 ;
  assign n2538 = n2482 ^ n2406 ^ 1'b0 ;
  assign n2539 = ( n2406 & n2537 ) | ( n2406 & ~n2538 ) | ( n2537 & ~n2538 ) ;
  assign n2540 = n2456 ^ n2351 ^ x81 ;
  assign n2541 = n2482 ^ n2351 ^ 1'b0 ;
  assign n2542 = ( n2351 & n2540 ) | ( n2351 & ~n2541 ) | ( n2540 & ~n2541 ) ;
  assign n2543 = n2455 ^ n2412 ^ x80 ;
  assign n2544 = n2482 ^ n2412 ^ 1'b0 ;
  assign n2545 = ( n2412 & n2543 ) | ( n2412 & ~n2544 ) | ( n2543 & ~n2544 ) ;
  assign n2546 = n2454 ^ n2354 ^ x79 ;
  assign n2547 = n2482 ^ n2354 ^ 1'b0 ;
  assign n2548 = ( n2354 & n2546 ) | ( n2354 & ~n2547 ) | ( n2546 & ~n2547 ) ;
  assign n2549 = n2450 ^ n2418 ^ x75 ;
  assign n2550 = n2482 ^ n2418 ^ 1'b0 ;
  assign n2551 = ( n2418 & n2549 ) | ( n2418 & ~n2550 ) | ( n2549 & ~n2550 ) ;
  assign n2552 = n2443 ^ n2424 ^ x71 ;
  assign n2553 = n2482 ^ n2424 ^ 1'b0 ;
  assign n2554 = ( n2424 & n2552 ) | ( n2424 & ~n2553 ) | ( n2552 & ~n2553 ) ;
  assign n2555 = n2441 ^ n2366 ^ x69 ;
  assign n2556 = n2482 ^ n2366 ^ 1'b0 ;
  assign n2557 = ( n2366 & n2555 ) | ( n2366 & ~n2556 ) | ( n2555 & ~n2556 ) ;
  assign n2558 = n2439 ^ n2371 ^ x67 ;
  assign n2559 = n2482 ^ n2371 ^ 1'b0 ;
  assign n2560 = ( n2371 & n2558 ) | ( n2371 & ~n2559 ) | ( n2558 & ~n2559 ) ;
  assign n2561 = n2429 & ~n2482 ;
  assign n2562 = x32 & x64 ;
  assign n2563 = ( ~x96 & n168 ) | ( ~x96 & n2562 ) | ( n168 & n2562 ) ;
  assign n2564 = ~n168 & n2563 ;
  assign n2565 = ( ~n197 & n2481 ) | ( ~n197 & n2564 ) | ( n2481 & n2564 ) ;
  assign n2566 = ~n2481 & n2565 ;
  assign n2567 = ( x32 & n2561 ) | ( x32 & ~n2566 ) | ( n2561 & ~n2566 ) ;
  assign n2568 = ~x31 & x64 ;
  assign n2569 = n2469 & n2482 ;
  assign n2570 = n322 | n2569 ;
  assign n2571 = ( ~x96 & n202 ) | ( ~x96 & n2570 ) | ( n202 & n2570 ) ;
  assign n2572 = n243 & n2570 ;
  assign n2573 = ( n243 & n322 ) | ( n243 & n2469 ) | ( n322 & n2469 ) ;
  assign n2574 = n2568 ^ n2567 ^ x65 ;
  assign n2575 = ( x65 & n2568 ) | ( x65 & n2574 ) | ( n2568 & n2574 ) ;
  assign n2576 = n2575 ^ n2524 ^ x66 ;
  assign n2577 = ( x66 & n2575 ) | ( x66 & n2576 ) | ( n2575 & n2576 ) ;
  assign n2578 = ( x67 & ~n2522 ) | ( x67 & n2577 ) | ( ~n2522 & n2577 ) ;
  assign n2579 = ( x68 & ~n2560 ) | ( x68 & n2578 ) | ( ~n2560 & n2578 ) ;
  assign n2580 = ( x69 & ~n2520 ) | ( x69 & n2579 ) | ( ~n2520 & n2579 ) ;
  assign n2581 = ( x70 & ~n2557 ) | ( x70 & n2580 ) | ( ~n2557 & n2580 ) ;
  assign n2582 = ( x71 & ~n2518 ) | ( x71 & n2581 ) | ( ~n2518 & n2581 ) ;
  assign n2583 = ( x72 & ~n2554 ) | ( x72 & n2582 ) | ( ~n2554 & n2582 ) ;
  assign n2584 = ( x73 & ~n2516 ) | ( x73 & n2583 ) | ( ~n2516 & n2583 ) ;
  assign n2585 = ( x74 & ~n2514 ) | ( x74 & n2584 ) | ( ~n2514 & n2584 ) ;
  assign n2586 = ( x75 & ~n2512 ) | ( x75 & n2585 ) | ( ~n2512 & n2585 ) ;
  assign n2587 = ( x76 & ~n2551 ) | ( x76 & n2586 ) | ( ~n2551 & n2586 ) ;
  assign n2588 = ( x77 & ~n2509 ) | ( x77 & n2587 ) | ( ~n2509 & n2587 ) ;
  assign n2589 = ( x78 & ~n2507 ) | ( x78 & n2588 ) | ( ~n2507 & n2588 ) ;
  assign n2590 = ( x79 & ~n2505 ) | ( x79 & n2589 ) | ( ~n2505 & n2589 ) ;
  assign n2591 = n2577 ^ n2522 ^ x67 ;
  assign n2592 = n2578 ^ n2560 ^ x68 ;
  assign n2593 = n2579 ^ n2520 ^ x69 ;
  assign n2594 = n2580 ^ n2557 ^ x70 ;
  assign n2595 = n2581 ^ n2518 ^ x71 ;
  assign n2596 = n2582 ^ n2554 ^ x72 ;
  assign n2597 = n2583 ^ n2516 ^ x73 ;
  assign n2598 = n2584 ^ n2514 ^ x74 ;
  assign n2599 = n2585 ^ n2512 ^ x75 ;
  assign n2600 = n2586 ^ n2551 ^ x76 ;
  assign n2601 = n2587 ^ n2509 ^ x77 ;
  assign n2602 = ( x96 & n202 ) | ( x96 & ~n2569 ) | ( n202 & ~n2569 ) ;
  assign n2603 = n2589 ^ n2505 ^ x79 ;
  assign n2604 = ( x80 & ~n2548 ) | ( x80 & n2590 ) | ( ~n2548 & n2590 ) ;
  assign n2605 = n2588 ^ n2507 ^ x78 ;
  assign n2606 = ( x81 & ~n2545 ) | ( x81 & n2604 ) | ( ~n2545 & n2604 ) ;
  assign n2607 = ( x82 & ~n2542 ) | ( x82 & n2606 ) | ( ~n2542 & n2606 ) ;
  assign n2608 = ( x83 & ~n2503 ) | ( x83 & n2607 ) | ( ~n2503 & n2607 ) ;
  assign n2609 = ( x84 & ~n2539 ) | ( x84 & n2608 ) | ( ~n2539 & n2608 ) ;
  assign n2610 = ( x85 & ~n2510 ) | ( x85 & n2609 ) | ( ~n2510 & n2609 ) ;
  assign n2611 = ( x86 & ~n2499 ) | ( x86 & n2610 ) | ( ~n2499 & n2610 ) ;
  assign n2612 = ( x87 & ~n2536 ) | ( x87 & n2611 ) | ( ~n2536 & n2611 ) ;
  assign n2613 = ( x88 & ~n2533 ) | ( x88 & n2612 ) | ( ~n2533 & n2612 ) ;
  assign n2614 = ( x89 & ~n2497 ) | ( x89 & n2613 ) | ( ~n2497 & n2613 ) ;
  assign n2615 = ( x90 & ~n2494 ) | ( x90 & n2614 ) | ( ~n2494 & n2614 ) ;
  assign n2616 = ( x91 & ~n2491 ) | ( x91 & n2615 ) | ( ~n2491 & n2615 ) ;
  assign n2617 = ( x92 & ~n2488 ) | ( x92 & n2616 ) | ( ~n2488 & n2616 ) ;
  assign n2618 = ( x93 & ~n2485 ) | ( x93 & n2617 ) | ( ~n2485 & n2617 ) ;
  assign n2619 = ( x94 & ~n2530 ) | ( x94 & n2618 ) | ( ~n2530 & n2618 ) ;
  assign n2620 = ( x95 & ~n2527 ) | ( x95 & n2619 ) | ( ~n2527 & n2619 ) ;
  assign n2621 = ( n2571 & n2602 ) | ( n2571 & ~n2620 ) | ( n2602 & ~n2620 ) ;
  assign n2622 = n2620 | n2621 ;
  assign n2623 = ( ~n2570 & n2572 ) | ( ~n2570 & n2622 ) | ( n2572 & n2622 ) ;
  assign n2624 = n2618 ^ n2530 ^ x94 ;
  assign n2625 = n2623 ^ n2530 ^ 1'b0 ;
  assign n2626 = ( n2530 & n2624 ) | ( n2530 & ~n2625 ) | ( n2624 & ~n2625 ) ;
  assign n2627 = n2623 ^ n2505 ^ 1'b0 ;
  assign n2628 = ( n2505 & n2603 ) | ( n2505 & ~n2627 ) | ( n2603 & ~n2627 ) ;
  assign n2629 = n2623 ^ n2507 ^ 1'b0 ;
  assign n2630 = ( n2507 & n2605 ) | ( n2507 & ~n2629 ) | ( n2605 & ~n2629 ) ;
  assign n2631 = n2623 ^ n2509 ^ 1'b0 ;
  assign n2632 = ( n2509 & n2601 ) | ( n2509 & ~n2631 ) | ( n2601 & ~n2631 ) ;
  assign n2633 = n2623 ^ n2551 ^ 1'b0 ;
  assign n2634 = ( n2551 & n2600 ) | ( n2551 & ~n2633 ) | ( n2600 & ~n2633 ) ;
  assign n2635 = n2623 ^ n2512 ^ 1'b0 ;
  assign n2636 = ( n2512 & n2599 ) | ( n2512 & ~n2635 ) | ( n2599 & ~n2635 ) ;
  assign n2637 = n2623 ^ n2514 ^ 1'b0 ;
  assign n2638 = ( n2514 & n2598 ) | ( n2514 & ~n2637 ) | ( n2598 & ~n2637 ) ;
  assign n2639 = n2623 ^ n2516 ^ 1'b0 ;
  assign n2640 = ( n2516 & n2597 ) | ( n2516 & ~n2639 ) | ( n2597 & ~n2639 ) ;
  assign n2641 = n2623 ^ n2554 ^ 1'b0 ;
  assign n2642 = ( n2554 & n2596 ) | ( n2554 & ~n2641 ) | ( n2596 & ~n2641 ) ;
  assign n2643 = n2623 ^ n2518 ^ 1'b0 ;
  assign n2644 = ( n2518 & n2595 ) | ( n2518 & ~n2643 ) | ( n2595 & ~n2643 ) ;
  assign n2645 = n2623 ^ n2557 ^ 1'b0 ;
  assign n2646 = ( n2557 & n2594 ) | ( n2557 & ~n2645 ) | ( n2594 & ~n2645 ) ;
  assign n2647 = n2623 ^ n2520 ^ 1'b0 ;
  assign n2648 = ( n2520 & n2593 ) | ( n2520 & ~n2647 ) | ( n2593 & ~n2647 ) ;
  assign n2649 = n2623 ^ n2560 ^ 1'b0 ;
  assign n2650 = ( n2560 & n2592 ) | ( n2560 & ~n2649 ) | ( n2592 & ~n2649 ) ;
  assign n2651 = n2623 ^ n2522 ^ 1'b0 ;
  assign n2652 = ( n2522 & n2591 ) | ( n2522 & ~n2651 ) | ( n2591 & ~n2651 ) ;
  assign n2653 = n2623 ^ n2576 ^ 1'b0 ;
  assign n2654 = ( n2524 & n2576 ) | ( n2524 & n2653 ) | ( n2576 & n2653 ) ;
  assign n2655 = n2623 ^ n2574 ^ 1'b0 ;
  assign n2656 = ( n2567 & n2574 ) | ( n2567 & n2655 ) | ( n2574 & n2655 ) ;
  assign n2657 = n322 | n2622 ;
  assign n2658 = ( n322 & n2573 ) | ( n322 & n2657 ) | ( n2573 & n2657 ) ;
  assign n2659 = n2619 ^ n2527 ^ x95 ;
  assign n2660 = n2623 ^ n2527 ^ 1'b0 ;
  assign n2661 = ( n2527 & n2659 ) | ( n2527 & ~n2660 ) | ( n2659 & ~n2660 ) ;
  assign n2662 = n2617 ^ n2485 ^ x93 ;
  assign n2663 = n2623 ^ n2485 ^ 1'b0 ;
  assign n2664 = ( n2485 & n2662 ) | ( n2485 & ~n2663 ) | ( n2662 & ~n2663 ) ;
  assign n2665 = n2616 ^ n2488 ^ x92 ;
  assign n2666 = n2623 ^ n2488 ^ 1'b0 ;
  assign n2667 = ( n2488 & n2665 ) | ( n2488 & ~n2666 ) | ( n2665 & ~n2666 ) ;
  assign n2668 = n2615 ^ n2491 ^ x91 ;
  assign n2669 = n2623 ^ n2491 ^ 1'b0 ;
  assign n2670 = ( n2491 & n2668 ) | ( n2491 & ~n2669 ) | ( n2668 & ~n2669 ) ;
  assign n2671 = n2614 ^ n2494 ^ x90 ;
  assign n2672 = n2623 ^ n2494 ^ 1'b0 ;
  assign n2673 = ( n2494 & n2671 ) | ( n2494 & ~n2672 ) | ( n2671 & ~n2672 ) ;
  assign n2674 = n2613 ^ n2497 ^ x89 ;
  assign n2675 = n2623 ^ n2497 ^ 1'b0 ;
  assign n2676 = ( n2497 & n2674 ) | ( n2497 & ~n2675 ) | ( n2674 & ~n2675 ) ;
  assign n2677 = n2612 ^ n2533 ^ x88 ;
  assign n2678 = n2623 ^ n2533 ^ 1'b0 ;
  assign n2679 = ( n2533 & n2677 ) | ( n2533 & ~n2678 ) | ( n2677 & ~n2678 ) ;
  assign n2680 = n2611 ^ n2536 ^ x87 ;
  assign n2681 = n2623 ^ n2536 ^ 1'b0 ;
  assign n2682 = ( n2536 & n2680 ) | ( n2536 & ~n2681 ) | ( n2680 & ~n2681 ) ;
  assign n2683 = n2610 ^ n2499 ^ x86 ;
  assign n2684 = n2623 ^ n2499 ^ 1'b0 ;
  assign n2685 = ( n2499 & n2683 ) | ( n2499 & ~n2684 ) | ( n2683 & ~n2684 ) ;
  assign n2686 = n2609 ^ n2510 ^ x85 ;
  assign n2687 = n2623 ^ n2510 ^ 1'b0 ;
  assign n2688 = ( n2510 & n2686 ) | ( n2510 & ~n2687 ) | ( n2686 & ~n2687 ) ;
  assign n2689 = n2608 ^ n2539 ^ x84 ;
  assign n2690 = n2623 ^ n2539 ^ 1'b0 ;
  assign n2691 = ( n2539 & n2689 ) | ( n2539 & ~n2690 ) | ( n2689 & ~n2690 ) ;
  assign n2692 = n2607 ^ n2503 ^ x83 ;
  assign n2693 = n2623 ^ n2503 ^ 1'b0 ;
  assign n2694 = ( n2503 & n2692 ) | ( n2503 & ~n2693 ) | ( n2692 & ~n2693 ) ;
  assign n2695 = n2606 ^ n2542 ^ x82 ;
  assign n2696 = n2623 ^ n2542 ^ 1'b0 ;
  assign n2697 = ( n2542 & n2695 ) | ( n2542 & ~n2696 ) | ( n2695 & ~n2696 ) ;
  assign n2698 = n2604 ^ n2545 ^ x81 ;
  assign n2699 = n2623 ^ n2545 ^ 1'b0 ;
  assign n2700 = ( n2545 & n2698 ) | ( n2545 & ~n2699 ) | ( n2698 & ~n2699 ) ;
  assign n2701 = n2590 ^ n2548 ^ x80 ;
  assign n2702 = n2623 ^ n2548 ^ 1'b0 ;
  assign n2703 = ( n2548 & n2701 ) | ( n2548 & ~n2702 ) | ( n2701 & ~n2702 ) ;
  assign n2704 = ~x30 & x64 ;
  assign n2705 = x64 & n2623 ;
  assign n2706 = n2705 ^ x64 ^ x31 ;
  assign n2707 = n2706 ^ n2704 ^ x65 ;
  assign n2708 = ( x65 & n2704 ) | ( x65 & n2707 ) | ( n2704 & n2707 ) ;
  assign n2709 = n2708 ^ n2656 ^ x66 ;
  assign n2710 = ( x66 & n2708 ) | ( x66 & n2709 ) | ( n2708 & n2709 ) ;
  assign n2711 = ( x67 & ~n2654 ) | ( x67 & n2710 ) | ( ~n2654 & n2710 ) ;
  assign n2712 = ( x68 & ~n2652 ) | ( x68 & n2711 ) | ( ~n2652 & n2711 ) ;
  assign n2713 = ( x69 & ~n2650 ) | ( x69 & n2712 ) | ( ~n2650 & n2712 ) ;
  assign n2714 = ( x70 & ~n2648 ) | ( x70 & n2713 ) | ( ~n2648 & n2713 ) ;
  assign n2715 = ( x71 & ~n2646 ) | ( x71 & n2714 ) | ( ~n2646 & n2714 ) ;
  assign n2716 = ( x72 & ~n2644 ) | ( x72 & n2715 ) | ( ~n2644 & n2715 ) ;
  assign n2717 = ( x73 & ~n2642 ) | ( x73 & n2716 ) | ( ~n2642 & n2716 ) ;
  assign n2718 = ( x74 & ~n2640 ) | ( x74 & n2717 ) | ( ~n2640 & n2717 ) ;
  assign n2719 = ( x75 & ~n2638 ) | ( x75 & n2718 ) | ( ~n2638 & n2718 ) ;
  assign n2720 = ( x76 & ~n2636 ) | ( x76 & n2719 ) | ( ~n2636 & n2719 ) ;
  assign n2721 = ( x77 & ~n2634 ) | ( x77 & n2720 ) | ( ~n2634 & n2720 ) ;
  assign n2722 = ( x78 & ~n2632 ) | ( x78 & n2721 ) | ( ~n2632 & n2721 ) ;
  assign n2723 = ( x79 & ~n2630 ) | ( x79 & n2722 ) | ( ~n2630 & n2722 ) ;
  assign n2724 = ( x80 & ~n2628 ) | ( x80 & n2723 ) | ( ~n2628 & n2723 ) ;
  assign n2725 = ( x81 & ~n2703 ) | ( x81 & n2724 ) | ( ~n2703 & n2724 ) ;
  assign n2726 = ( x82 & ~n2700 ) | ( x82 & n2725 ) | ( ~n2700 & n2725 ) ;
  assign n2727 = ( x83 & ~n2697 ) | ( x83 & n2726 ) | ( ~n2697 & n2726 ) ;
  assign n2728 = ( x84 & ~n2694 ) | ( x84 & n2727 ) | ( ~n2694 & n2727 ) ;
  assign n2729 = ( x85 & ~n2691 ) | ( x85 & n2728 ) | ( ~n2691 & n2728 ) ;
  assign n2730 = ( x86 & ~n2688 ) | ( x86 & n2729 ) | ( ~n2688 & n2729 ) ;
  assign n2731 = ( x87 & ~n2685 ) | ( x87 & n2730 ) | ( ~n2685 & n2730 ) ;
  assign n2732 = ( x88 & ~n2682 ) | ( x88 & n2731 ) | ( ~n2682 & n2731 ) ;
  assign n2733 = ( x89 & ~n2679 ) | ( x89 & n2732 ) | ( ~n2679 & n2732 ) ;
  assign n2734 = ( x90 & ~n2676 ) | ( x90 & n2733 ) | ( ~n2676 & n2733 ) ;
  assign n2735 = ( x91 & ~n2673 ) | ( x91 & n2734 ) | ( ~n2673 & n2734 ) ;
  assign n2736 = ( x92 & ~n2670 ) | ( x92 & n2735 ) | ( ~n2670 & n2735 ) ;
  assign n2737 = ( x93 & ~n2667 ) | ( x93 & n2736 ) | ( ~n2667 & n2736 ) ;
  assign n2738 = ( x94 & ~n2664 ) | ( x94 & n2737 ) | ( ~n2664 & n2737 ) ;
  assign n2739 = ( x95 & ~n2626 ) | ( x95 & n2738 ) | ( ~n2626 & n2738 ) ;
  assign n2740 = ( ~x98 & x99 ) | ( ~x98 & n188 ) | ( x99 & n188 ) ;
  assign n2741 = x98 | n2740 ;
  assign n2742 = ( x96 & ~n2661 ) | ( x96 & n2739 ) | ( ~n2661 & n2739 ) ;
  assign n2743 = ( x97 & ~n2658 ) | ( x97 & n2742 ) | ( ~n2658 & n2742 ) ;
  assign n2744 = n183 | n194 ;
  assign n2745 = ( ~n2741 & n2743 ) | ( ~n2741 & n2744 ) | ( n2743 & n2744 ) ;
  assign n2746 = n2741 | n2745 ;
  assign n2747 = n2724 ^ n2703 ^ x81 ;
  assign n2748 = n2746 ^ n2703 ^ 1'b0 ;
  assign n2749 = ( n2703 & n2747 ) | ( n2703 & ~n2748 ) | ( n2747 & ~n2748 ) ;
  assign n2750 = n2723 ^ n2628 ^ x80 ;
  assign n2751 = n2746 ^ n2628 ^ 1'b0 ;
  assign n2752 = ( n2628 & n2750 ) | ( n2628 & ~n2751 ) | ( n2750 & ~n2751 ) ;
  assign n2753 = n2720 ^ n2634 ^ x77 ;
  assign n2754 = n2746 ^ n2634 ^ 1'b0 ;
  assign n2755 = ( n2634 & n2753 ) | ( n2634 & ~n2754 ) | ( n2753 & ~n2754 ) ;
  assign n2756 = n2718 ^ n2638 ^ x75 ;
  assign n2757 = n2746 ^ n2638 ^ 1'b0 ;
  assign n2758 = ( n2638 & n2756 ) | ( n2638 & ~n2757 ) | ( n2756 & ~n2757 ) ;
  assign n2759 = n2715 ^ n2644 ^ x72 ;
  assign n2760 = n2746 ^ n2644 ^ 1'b0 ;
  assign n2761 = ( n2644 & n2759 ) | ( n2644 & ~n2760 ) | ( n2759 & ~n2760 ) ;
  assign n2762 = n2712 ^ n2650 ^ x69 ;
  assign n2763 = n2746 ^ n2650 ^ 1'b0 ;
  assign n2764 = ( n2650 & n2762 ) | ( n2650 & ~n2763 ) | ( n2762 & ~n2763 ) ;
  assign n2765 = n2711 ^ n2652 ^ x68 ;
  assign n2766 = n2746 ^ n2652 ^ 1'b0 ;
  assign n2767 = ( n2652 & n2765 ) | ( n2652 & ~n2766 ) | ( n2765 & ~n2766 ) ;
  assign n2768 = n2710 ^ n2654 ^ x67 ;
  assign n2769 = n2746 ^ n2654 ^ 1'b0 ;
  assign n2770 = ( n2654 & n2768 ) | ( n2654 & ~n2769 ) | ( n2768 & ~n2769 ) ;
  assign n2771 = n2746 ^ n2709 ^ 1'b0 ;
  assign n2772 = ( n2656 & n2709 ) | ( n2656 & n2771 ) | ( n2709 & n2771 ) ;
  assign n2773 = n2746 ^ n2707 ^ 1'b0 ;
  assign n2774 = ( n2706 & n2707 ) | ( n2706 & n2773 ) | ( n2707 & n2773 ) ;
  assign n2775 = n2739 ^ n2661 ^ x96 ;
  assign n2776 = n2775 ^ n2746 ^ 1'b0 ;
  assign n2777 = ( n2661 & n2775 ) | ( n2661 & n2776 ) | ( n2775 & n2776 ) ;
  assign n2778 = n2738 ^ n2626 ^ x95 ;
  assign n2779 = n2746 ^ n2626 ^ 1'b0 ;
  assign n2780 = ( n2626 & n2778 ) | ( n2626 & ~n2779 ) | ( n2778 & ~n2779 ) ;
  assign n2781 = n2737 ^ n2664 ^ x94 ;
  assign n2782 = n2746 ^ n2664 ^ 1'b0 ;
  assign n2783 = ( n2664 & n2781 ) | ( n2664 & ~n2782 ) | ( n2781 & ~n2782 ) ;
  assign n2784 = n2735 ^ n2670 ^ x92 ;
  assign n2785 = n2746 ^ n2670 ^ 1'b0 ;
  assign n2786 = ( n2670 & n2784 ) | ( n2670 & ~n2785 ) | ( n2784 & ~n2785 ) ;
  assign n2787 = n2734 ^ n2673 ^ x91 ;
  assign n2788 = n2746 ^ n2673 ^ 1'b0 ;
  assign n2789 = ( n2673 & n2787 ) | ( n2673 & ~n2788 ) | ( n2787 & ~n2788 ) ;
  assign n2790 = n2733 ^ n2676 ^ x90 ;
  assign n2791 = n2746 ^ n2676 ^ 1'b0 ;
  assign n2792 = ( n2676 & n2790 ) | ( n2676 & ~n2791 ) | ( n2790 & ~n2791 ) ;
  assign n2793 = n2732 ^ n2679 ^ x89 ;
  assign n2794 = n2746 ^ n2679 ^ 1'b0 ;
  assign n2795 = ( n2679 & n2793 ) | ( n2679 & ~n2794 ) | ( n2793 & ~n2794 ) ;
  assign n2796 = n2731 ^ n2682 ^ x88 ;
  assign n2797 = n2746 ^ n2682 ^ 1'b0 ;
  assign n2798 = ( n2682 & n2796 ) | ( n2682 & ~n2797 ) | ( n2796 & ~n2797 ) ;
  assign n2799 = n2730 ^ n2685 ^ x87 ;
  assign n2800 = n2746 ^ n2685 ^ 1'b0 ;
  assign n2801 = ( n2685 & n2799 ) | ( n2685 & ~n2800 ) | ( n2799 & ~n2800 ) ;
  assign n2802 = n2729 ^ n2688 ^ x86 ;
  assign n2803 = n2746 ^ n2688 ^ 1'b0 ;
  assign n2804 = ( n2688 & n2802 ) | ( n2688 & ~n2803 ) | ( n2802 & ~n2803 ) ;
  assign n2805 = n2728 ^ n2691 ^ x85 ;
  assign n2806 = n2746 ^ n2691 ^ 1'b0 ;
  assign n2807 = ( n2691 & n2805 ) | ( n2691 & ~n2806 ) | ( n2805 & ~n2806 ) ;
  assign n2808 = n2727 ^ n2694 ^ x84 ;
  assign n2809 = n2746 ^ n2694 ^ 1'b0 ;
  assign n2810 = ( n2694 & n2808 ) | ( n2694 & ~n2809 ) | ( n2808 & ~n2809 ) ;
  assign n2811 = n2726 ^ n2697 ^ x83 ;
  assign n2812 = n2746 ^ n2697 ^ 1'b0 ;
  assign n2813 = ( n2697 & n2811 ) | ( n2697 & ~n2812 ) | ( n2811 & ~n2812 ) ;
  assign n2814 = n2725 ^ n2700 ^ x82 ;
  assign n2815 = n2746 ^ n2700 ^ 1'b0 ;
  assign n2816 = ( n2700 & n2814 ) | ( n2700 & ~n2815 ) | ( n2814 & ~n2815 ) ;
  assign n2817 = n2721 ^ n2632 ^ x78 ;
  assign n2818 = n2746 ^ n2632 ^ 1'b0 ;
  assign n2819 = ( n2632 & n2817 ) | ( n2632 & ~n2818 ) | ( n2817 & ~n2818 ) ;
  assign n2820 = n2719 ^ n2636 ^ x76 ;
  assign n2821 = n2746 ^ n2636 ^ 1'b0 ;
  assign n2822 = ( n2636 & n2820 ) | ( n2636 & ~n2821 ) | ( n2820 & ~n2821 ) ;
  assign n2823 = n2717 ^ n2640 ^ x74 ;
  assign n2824 = n2746 ^ n2640 ^ 1'b0 ;
  assign n2825 = ( n2640 & n2823 ) | ( n2640 & ~n2824 ) | ( n2823 & ~n2824 ) ;
  assign n2826 = n2716 ^ n2642 ^ x73 ;
  assign n2827 = n2746 ^ n2642 ^ 1'b0 ;
  assign n2828 = ( n2642 & n2826 ) | ( n2642 & ~n2827 ) | ( n2826 & ~n2827 ) ;
  assign n2829 = n2714 ^ n2646 ^ x71 ;
  assign n2830 = n2746 ^ n2646 ^ 1'b0 ;
  assign n2831 = ( n2646 & n2829 ) | ( n2646 & ~n2830 ) | ( n2829 & ~n2830 ) ;
  assign n2832 = n2713 ^ n2648 ^ x70 ;
  assign n2833 = n2746 ^ n2648 ^ 1'b0 ;
  assign n2834 = ( n2648 & n2832 ) | ( n2648 & ~n2833 ) | ( n2832 & ~n2833 ) ;
  assign n2835 = n2704 | n2746 ;
  assign n2836 = ~x29 & x64 ;
  assign n2837 = ( x30 & x98 ) | ( x30 & n162 ) | ( x98 & n162 ) ;
  assign n2838 = n2722 ^ n2630 ^ x79 ;
  assign n2839 = n2746 ^ n2630 ^ 1'b0 ;
  assign n2840 = ( x30 & n191 ) | ( x30 & n2743 ) | ( n191 & n2743 ) ;
  assign n2841 = n2746 ^ n2667 ^ 1'b0 ;
  assign n2842 = n162 | n191 ;
  assign n2843 = ( x30 & n2837 ) | ( x30 & n2840 ) | ( n2837 & n2840 ) ;
  assign n2844 = x30 & ~x64 ;
  assign n2845 = ( x30 & n2843 ) | ( x30 & n2844 ) | ( n2843 & n2844 ) ;
  assign n2846 = ( ~n2746 & n2835 ) | ( ~n2746 & n2845 ) | ( n2835 & n2845 ) ;
  assign n2847 = n2846 ^ n2836 ^ x65 ;
  assign n2848 = ( x65 & n2836 ) | ( x65 & n2847 ) | ( n2836 & n2847 ) ;
  assign n2849 = ( n2630 & n2838 ) | ( n2630 & ~n2839 ) | ( n2838 & ~n2839 ) ;
  assign n2850 = n2848 ^ n2774 ^ x66 ;
  assign n2851 = ( x66 & n2848 ) | ( x66 & n2850 ) | ( n2848 & n2850 ) ;
  assign n2852 = ( x67 & ~n2772 ) | ( x67 & n2851 ) | ( ~n2772 & n2851 ) ;
  assign n2853 = ( x68 & ~n2770 ) | ( x68 & n2852 ) | ( ~n2770 & n2852 ) ;
  assign n2854 = ( x69 & ~n2767 ) | ( x69 & n2853 ) | ( ~n2767 & n2853 ) ;
  assign n2855 = ( x70 & ~n2764 ) | ( x70 & n2854 ) | ( ~n2764 & n2854 ) ;
  assign n2856 = ( x71 & ~n2834 ) | ( x71 & n2855 ) | ( ~n2834 & n2855 ) ;
  assign n2857 = ( x72 & ~n2831 ) | ( x72 & n2856 ) | ( ~n2831 & n2856 ) ;
  assign n2858 = ( x73 & ~n2761 ) | ( x73 & n2857 ) | ( ~n2761 & n2857 ) ;
  assign n2859 = ( x74 & ~n2828 ) | ( x74 & n2858 ) | ( ~n2828 & n2858 ) ;
  assign n2860 = ( x75 & ~n2825 ) | ( x75 & n2859 ) | ( ~n2825 & n2859 ) ;
  assign n2861 = ( x76 & ~n2758 ) | ( x76 & n2860 ) | ( ~n2758 & n2860 ) ;
  assign n2862 = ( x77 & ~n2822 ) | ( x77 & n2861 ) | ( ~n2822 & n2861 ) ;
  assign n2863 = ( x78 & ~n2755 ) | ( x78 & n2862 ) | ( ~n2755 & n2862 ) ;
  assign n2864 = ( x79 & ~n2819 ) | ( x79 & n2863 ) | ( ~n2819 & n2863 ) ;
  assign n2865 = ( x80 & ~n2849 ) | ( x80 & n2864 ) | ( ~n2849 & n2864 ) ;
  assign n2866 = ( x81 & ~n2752 ) | ( x81 & n2865 ) | ( ~n2752 & n2865 ) ;
  assign n2867 = n2736 ^ n2667 ^ x93 ;
  assign n2868 = ( x82 & ~n2749 ) | ( x82 & n2866 ) | ( ~n2749 & n2866 ) ;
  assign n2869 = ( x83 & ~n2816 ) | ( x83 & n2868 ) | ( ~n2816 & n2868 ) ;
  assign n2870 = n2856 ^ n2831 ^ x72 ;
  assign n2871 = n2854 ^ n2764 ^ x70 ;
  assign n2872 = n2861 ^ n2822 ^ x77 ;
  assign n2873 = n2862 ^ n2755 ^ x78 ;
  assign n2874 = n2863 ^ n2819 ^ x79 ;
  assign n2875 = n2857 ^ n2761 ^ x73 ;
  assign n2876 = n2858 ^ n2828 ^ x74 ;
  assign n2877 = ( x84 & ~n2813 ) | ( x84 & n2869 ) | ( ~n2813 & n2869 ) ;
  assign n2878 = ( n322 & n2658 ) | ( n322 & n2746 ) | ( n2658 & n2746 ) ;
  assign n2879 = n2869 ^ n2813 ^ x84 ;
  assign n2880 = ( n2667 & ~n2841 ) | ( n2667 & n2867 ) | ( ~n2841 & n2867 ) ;
  assign n2881 = ( x85 & ~n2810 ) | ( x85 & n2877 ) | ( ~n2810 & n2877 ) ;
  assign n2882 = ( x86 & ~n2807 ) | ( x86 & n2881 ) | ( ~n2807 & n2881 ) ;
  assign n2883 = ( x87 & ~n2804 ) | ( x87 & n2882 ) | ( ~n2804 & n2882 ) ;
  assign n2884 = ( x88 & ~n2801 ) | ( x88 & n2883 ) | ( ~n2801 & n2883 ) ;
  assign n2885 = ( x89 & ~n2798 ) | ( x89 & n2884 ) | ( ~n2798 & n2884 ) ;
  assign n2886 = ( x90 & ~n2795 ) | ( x90 & n2885 ) | ( ~n2795 & n2885 ) ;
  assign n2887 = ( x91 & ~n2792 ) | ( x91 & n2886 ) | ( ~n2792 & n2886 ) ;
  assign n2888 = ( x92 & ~n2789 ) | ( x92 & n2887 ) | ( ~n2789 & n2887 ) ;
  assign n2889 = n2887 ^ n2789 ^ x92 ;
  assign n2890 = ( x93 & ~n2786 ) | ( x93 & n2888 ) | ( ~n2786 & n2888 ) ;
  assign n2891 = ( x94 & ~n2880 ) | ( x94 & n2890 ) | ( ~n2880 & n2890 ) ;
  assign n2892 = n2888 ^ n2786 ^ x93 ;
  assign n2893 = ( x95 & ~n2783 ) | ( x95 & n2891 ) | ( ~n2783 & n2891 ) ;
  assign n2894 = ( x96 & ~n2780 ) | ( x96 & n2893 ) | ( ~n2780 & n2893 ) ;
  assign n2895 = ( x97 & ~n2777 ) | ( x97 & n2894 ) | ( ~n2777 & n2894 ) ;
  assign n2896 = ( x98 & ~n2878 ) | ( x98 & n2895 ) | ( ~n2878 & n2895 ) ;
  assign n2897 = ( x64 & ~x99 ) | ( x64 & n2896 ) | ( ~x99 & n2896 ) ;
  assign n2898 = n2891 ^ n2783 ^ x95 ;
  assign n2899 = ( ~n188 & n194 ) | ( ~n188 & n2897 ) | ( n194 & n2897 ) ;
  assign n2900 = n2842 | n2896 ;
  assign n2901 = n2900 ^ n2789 ^ 1'b0 ;
  assign n2902 = ( n2789 & n2889 ) | ( n2789 & ~n2901 ) | ( n2889 & ~n2901 ) ;
  assign n2903 = n2900 ^ n2831 ^ 1'b0 ;
  assign n2904 = n2900 ^ n2783 ^ 1'b0 ;
  assign n2905 = ( n2783 & n2898 ) | ( n2783 & ~n2904 ) | ( n2898 & ~n2904 ) ;
  assign n2906 = n2900 ^ n2828 ^ 1'b0 ;
  assign n2907 = n2900 ^ n2786 ^ 1'b0 ;
  assign n2908 = n2836 | n2900 ;
  assign n2909 = ( n2786 & n2892 ) | ( n2786 & ~n2907 ) | ( n2892 & ~n2907 ) ;
  assign n2910 = n2900 ^ n2847 ^ 1'b0 ;
  assign n2911 = n2900 ^ n2795 ^ 1'b0 ;
  assign n2912 = n2885 ^ n2795 ^ x90 ;
  assign n2913 = ( n2846 & n2847 ) | ( n2846 & n2910 ) | ( n2847 & n2910 ) ;
  assign n2914 = n2900 ^ n2780 ^ 1'b0 ;
  assign n2915 = n2900 ^ n2761 ^ 1'b0 ;
  assign n2916 = ( n2795 & ~n2911 ) | ( n2795 & n2912 ) | ( ~n2911 & n2912 ) ;
  assign n2917 = n2893 ^ n2780 ^ x96 ;
  assign n2918 = n2900 ^ n2880 ^ 1'b0 ;
  assign n2919 = n2884 ^ n2798 ^ x89 ;
  assign n2920 = n2886 ^ n2792 ^ x91 ;
  assign n2921 = n2900 ^ n2798 ^ 1'b0 ;
  assign n2922 = ( n2798 & n2919 ) | ( n2798 & ~n2921 ) | ( n2919 & ~n2921 ) ;
  assign n2923 = n2900 ^ n2822 ^ 1'b0 ;
  assign n2924 = ( n2822 & n2872 ) | ( n2822 & ~n2923 ) | ( n2872 & ~n2923 ) ;
  assign n2925 = n2900 ^ n2764 ^ 1'b0 ;
  assign n2926 = ( n2828 & n2876 ) | ( n2828 & ~n2906 ) | ( n2876 & ~n2906 ) ;
  assign n2927 = n2900 ^ n2819 ^ 1'b0 ;
  assign n2928 = ( n2831 & n2870 ) | ( n2831 & ~n2903 ) | ( n2870 & ~n2903 ) ;
  assign n2929 = n2900 ^ n2813 ^ 1'b0 ;
  assign n2930 = n2900 ^ n2755 ^ 1'b0 ;
  assign n2931 = ( n2780 & ~n2914 ) | ( n2780 & n2917 ) | ( ~n2914 & n2917 ) ;
  assign n2932 = n2890 ^ n2880 ^ x94 ;
  assign n2933 = ( n2755 & n2873 ) | ( n2755 & ~n2930 ) | ( n2873 & ~n2930 ) ;
  assign n2934 = ( n2813 & n2879 ) | ( n2813 & ~n2929 ) | ( n2879 & ~n2929 ) ;
  assign n2935 = n2744 & ~n2896 ;
  assign n2936 = ( n2880 & ~n2918 ) | ( n2880 & n2932 ) | ( ~n2918 & n2932 ) ;
  assign n2937 = ( n2761 & n2875 ) | ( n2761 & ~n2915 ) | ( n2875 & ~n2915 ) ;
  assign n2938 = ( n2896 & n2899 ) | ( n2896 & ~n2935 ) | ( n2899 & ~n2935 ) ;
  assign n2939 = ( n2819 & n2874 ) | ( n2819 & ~n2927 ) | ( n2874 & ~n2927 ) ;
  assign n2940 = ( x29 & n2896 ) | ( x29 & ~n2938 ) | ( n2896 & ~n2938 ) ;
  assign n2941 = ( ~n2900 & n2908 ) | ( ~n2900 & n2940 ) | ( n2908 & n2940 ) ;
  assign n2942 = ( n2764 & n2871 ) | ( n2764 & ~n2925 ) | ( n2871 & ~n2925 ) ;
  assign n2943 = n2894 ^ n2777 ^ x97 ;
  assign n2944 = n2943 ^ n2900 ^ 1'b0 ;
  assign n2945 = ( n2777 & n2943 ) | ( n2777 & n2944 ) | ( n2943 & n2944 ) ;
  assign n2946 = n2900 ^ n2792 ^ 1'b0 ;
  assign n2947 = n2883 ^ n2801 ^ x88 ;
  assign n2948 = n2900 ^ n2801 ^ 1'b0 ;
  assign n2949 = ( n2801 & n2947 ) | ( n2801 & ~n2948 ) | ( n2947 & ~n2948 ) ;
  assign n2950 = n2882 ^ n2804 ^ x87 ;
  assign n2951 = n2900 ^ n2804 ^ 1'b0 ;
  assign n2952 = ( n2804 & n2950 ) | ( n2804 & ~n2951 ) | ( n2950 & ~n2951 ) ;
  assign n2953 = n2881 ^ n2807 ^ x86 ;
  assign n2954 = n2900 ^ n2807 ^ 1'b0 ;
  assign n2955 = ( n2807 & n2953 ) | ( n2807 & ~n2954 ) | ( n2953 & ~n2954 ) ;
  assign n2956 = n2877 ^ n2810 ^ x85 ;
  assign n2957 = n2900 ^ n2810 ^ 1'b0 ;
  assign n2958 = ( n2810 & n2956 ) | ( n2810 & ~n2957 ) | ( n2956 & ~n2957 ) ;
  assign n2959 = ( n2792 & n2920 ) | ( n2792 & ~n2946 ) | ( n2920 & ~n2946 ) ;
  assign n2960 = n2868 ^ n2816 ^ x83 ;
  assign n2961 = n2900 ^ n2816 ^ 1'b0 ;
  assign n2962 = ( n2816 & n2960 ) | ( n2816 & ~n2961 ) | ( n2960 & ~n2961 ) ;
  assign n2963 = n2866 ^ n2749 ^ x82 ;
  assign n2964 = n2900 ^ n2749 ^ 1'b0 ;
  assign n2965 = ( n2749 & n2963 ) | ( n2749 & ~n2964 ) | ( n2963 & ~n2964 ) ;
  assign n2966 = n2865 ^ n2752 ^ x81 ;
  assign n2967 = n2900 ^ n2752 ^ 1'b0 ;
  assign n2968 = ( n2752 & n2966 ) | ( n2752 & ~n2967 ) | ( n2966 & ~n2967 ) ;
  assign n2969 = n2864 ^ n2849 ^ x80 ;
  assign n2970 = n2900 ^ n2849 ^ 1'b0 ;
  assign n2971 = ( n2849 & n2969 ) | ( n2849 & ~n2970 ) | ( n2969 & ~n2970 ) ;
  assign n2972 = n2860 ^ n2758 ^ x76 ;
  assign n2973 = n2900 ^ n2758 ^ 1'b0 ;
  assign n2974 = ( n2758 & n2972 ) | ( n2758 & ~n2973 ) | ( n2972 & ~n2973 ) ;
  assign n2975 = n2859 ^ n2825 ^ x75 ;
  assign n2976 = n2900 ^ n2825 ^ 1'b0 ;
  assign n2977 = ( n2825 & n2975 ) | ( n2825 & ~n2976 ) | ( n2975 & ~n2976 ) ;
  assign n2978 = n2855 ^ n2834 ^ x71 ;
  assign n2979 = n2900 ^ n2834 ^ 1'b0 ;
  assign n2980 = ( n2834 & n2978 ) | ( n2834 & ~n2979 ) | ( n2978 & ~n2979 ) ;
  assign n2981 = n2853 ^ n2767 ^ x69 ;
  assign n2982 = n2900 ^ n2767 ^ 1'b0 ;
  assign n2983 = ( n2767 & n2981 ) | ( n2767 & ~n2982 ) | ( n2981 & ~n2982 ) ;
  assign n2984 = n2852 ^ n2770 ^ x68 ;
  assign n2985 = n2900 ^ n2770 ^ 1'b0 ;
  assign n2986 = ( n2770 & n2984 ) | ( n2770 & ~n2985 ) | ( n2984 & ~n2985 ) ;
  assign n2987 = n2851 ^ n2772 ^ x67 ;
  assign n2988 = n2900 ^ n2772 ^ 1'b0 ;
  assign n2989 = ( n2772 & n2987 ) | ( n2772 & ~n2988 ) | ( n2987 & ~n2988 ) ;
  assign n2990 = n2878 & n2900 ;
  assign n2991 = ~x28 & x64 ;
  assign n2992 = n322 | n2990 ;
  assign n2993 = n2991 ^ n2941 ^ x65 ;
  assign n2994 = ( x65 & n2991 ) | ( x65 & n2993 ) | ( n2991 & n2993 ) ;
  assign n2995 = n2994 ^ n2913 ^ x66 ;
  assign n2996 = n2900 ^ n2850 ^ 1'b0 ;
  assign n2997 = ( n2774 & n2850 ) | ( n2774 & n2996 ) | ( n2850 & n2996 ) ;
  assign n2998 = ( x66 & n2994 ) | ( x66 & n2995 ) | ( n2994 & n2995 ) ;
  assign n2999 = ( x67 & ~n2997 ) | ( x67 & n2998 ) | ( ~n2997 & n2998 ) ;
  assign n3000 = ( x68 & ~n2989 ) | ( x68 & n2999 ) | ( ~n2989 & n2999 ) ;
  assign n3001 = ( x69 & ~n2986 ) | ( x69 & n3000 ) | ( ~n2986 & n3000 ) ;
  assign n3002 = ( x70 & ~n2983 ) | ( x70 & n3001 ) | ( ~n2983 & n3001 ) ;
  assign n3003 = ( x71 & ~n2942 ) | ( x71 & n3002 ) | ( ~n2942 & n3002 ) ;
  assign n3004 = ( x72 & ~n2980 ) | ( x72 & n3003 ) | ( ~n2980 & n3003 ) ;
  assign n3005 = ( x73 & ~n2928 ) | ( x73 & n3004 ) | ( ~n2928 & n3004 ) ;
  assign n3006 = ( x74 & ~n2937 ) | ( x74 & n3005 ) | ( ~n2937 & n3005 ) ;
  assign n3007 = ( x75 & ~n2926 ) | ( x75 & n3006 ) | ( ~n2926 & n3006 ) ;
  assign n3008 = ( x76 & ~n2977 ) | ( x76 & n3007 ) | ( ~n2977 & n3007 ) ;
  assign n3009 = ( x77 & ~n2974 ) | ( x77 & n3008 ) | ( ~n2974 & n3008 ) ;
  assign n3010 = n2842 & n2992 ;
  assign n3011 = ( n322 & n2842 ) | ( n322 & n2878 ) | ( n2842 & n2878 ) ;
  assign n3012 = ( x78 & ~n2924 ) | ( x78 & n3009 ) | ( ~n2924 & n3009 ) ;
  assign n3013 = ( x79 & ~n2933 ) | ( x79 & n3012 ) | ( ~n2933 & n3012 ) ;
  assign n3014 = ( x80 & ~n2939 ) | ( x80 & n3013 ) | ( ~n2939 & n3013 ) ;
  assign n3015 = ( ~x99 & n199 ) | ( ~x99 & n2992 ) | ( n199 & n2992 ) ;
  assign n3016 = n2998 ^ n2997 ^ x67 ;
  assign n3017 = n2999 ^ n2989 ^ x68 ;
  assign n3018 = n3000 ^ n2986 ^ x69 ;
  assign n3019 = n3001 ^ n2983 ^ x70 ;
  assign n3020 = n3002 ^ n2942 ^ x71 ;
  assign n3021 = n3003 ^ n2980 ^ x72 ;
  assign n3022 = n3004 ^ n2928 ^ x73 ;
  assign n3023 = n3005 ^ n2937 ^ x74 ;
  assign n3024 = n3006 ^ n2926 ^ x75 ;
  assign n3025 = n3007 ^ n2977 ^ x76 ;
  assign n3026 = n3008 ^ n2974 ^ x77 ;
  assign n3027 = n3009 ^ n2924 ^ x78 ;
  assign n3028 = ( x99 & n199 ) | ( x99 & ~n2990 ) | ( n199 & ~n2990 ) ;
  assign n3029 = n3013 ^ n2939 ^ x80 ;
  assign n3030 = ( x81 & ~n2971 ) | ( x81 & n3014 ) | ( ~n2971 & n3014 ) ;
  assign n3031 = n3012 ^ n2933 ^ x79 ;
  assign n3032 = ( x82 & ~n2968 ) | ( x82 & n3030 ) | ( ~n2968 & n3030 ) ;
  assign n3033 = ( x83 & ~n2965 ) | ( x83 & n3032 ) | ( ~n2965 & n3032 ) ;
  assign n3034 = ( x84 & ~n2962 ) | ( x84 & n3033 ) | ( ~n2962 & n3033 ) ;
  assign n3035 = ( x85 & ~n2934 ) | ( x85 & n3034 ) | ( ~n2934 & n3034 ) ;
  assign n3036 = ( x86 & ~n2958 ) | ( x86 & n3035 ) | ( ~n2958 & n3035 ) ;
  assign n3037 = ( x87 & ~n2955 ) | ( x87 & n3036 ) | ( ~n2955 & n3036 ) ;
  assign n3038 = ( x88 & ~n2952 ) | ( x88 & n3037 ) | ( ~n2952 & n3037 ) ;
  assign n3039 = ( x89 & ~n2949 ) | ( x89 & n3038 ) | ( ~n2949 & n3038 ) ;
  assign n3040 = ( x90 & ~n2922 ) | ( x90 & n3039 ) | ( ~n2922 & n3039 ) ;
  assign n3041 = ( x91 & ~n2916 ) | ( x91 & n3040 ) | ( ~n2916 & n3040 ) ;
  assign n3042 = ( x92 & ~n2959 ) | ( x92 & n3041 ) | ( ~n2959 & n3041 ) ;
  assign n3043 = ( x93 & ~n2902 ) | ( x93 & n3042 ) | ( ~n2902 & n3042 ) ;
  assign n3044 = ( x94 & ~n2909 ) | ( x94 & n3043 ) | ( ~n2909 & n3043 ) ;
  assign n3045 = ( x95 & ~n2936 ) | ( x95 & n3044 ) | ( ~n2936 & n3044 ) ;
  assign n3046 = ( x96 & ~n2905 ) | ( x96 & n3045 ) | ( ~n2905 & n3045 ) ;
  assign n3047 = ( x97 & ~n2931 ) | ( x97 & n3046 ) | ( ~n2931 & n3046 ) ;
  assign n3048 = ( x98 & ~n2945 ) | ( x98 & n3047 ) | ( ~n2945 & n3047 ) ;
  assign n3049 = ( n3015 & n3028 ) | ( n3015 & ~n3048 ) | ( n3028 & ~n3048 ) ;
  assign n3050 = n3048 | n3049 ;
  assign n3051 = ( ~n2992 & n3010 ) | ( ~n2992 & n3050 ) | ( n3010 & n3050 ) ;
  assign n3052 = n3046 ^ n2931 ^ x97 ;
  assign n3053 = n3051 ^ n2931 ^ 1'b0 ;
  assign n3054 = ( n2931 & n3052 ) | ( n2931 & ~n3053 ) | ( n3052 & ~n3053 ) ;
  assign n3055 = n3030 ^ n2968 ^ x82 ;
  assign n3056 = n3051 ^ n2968 ^ 1'b0 ;
  assign n3057 = ( n2968 & n3055 ) | ( n2968 & ~n3056 ) | ( n3055 & ~n3056 ) ;
  assign n3058 = n3051 ^ n2939 ^ 1'b0 ;
  assign n3059 = ( n2939 & n3029 ) | ( n2939 & ~n3058 ) | ( n3029 & ~n3058 ) ;
  assign n3060 = n3051 ^ n2933 ^ 1'b0 ;
  assign n3061 = ( n2933 & n3031 ) | ( n2933 & ~n3060 ) | ( n3031 & ~n3060 ) ;
  assign n3062 = n3051 ^ n2924 ^ 1'b0 ;
  assign n3063 = ( n2924 & n3027 ) | ( n2924 & ~n3062 ) | ( n3027 & ~n3062 ) ;
  assign n3064 = n3051 ^ n2977 ^ 1'b0 ;
  assign n3065 = ( n2977 & n3025 ) | ( n2977 & ~n3064 ) | ( n3025 & ~n3064 ) ;
  assign n3066 = n3051 ^ n2926 ^ 1'b0 ;
  assign n3067 = ( n2926 & n3024 ) | ( n2926 & ~n3066 ) | ( n3024 & ~n3066 ) ;
  assign n3068 = n3051 ^ n2937 ^ 1'b0 ;
  assign n3069 = ( n2937 & n3023 ) | ( n2937 & ~n3068 ) | ( n3023 & ~n3068 ) ;
  assign n3070 = n3051 ^ n2928 ^ 1'b0 ;
  assign n3071 = ( n2928 & n3022 ) | ( n2928 & ~n3070 ) | ( n3022 & ~n3070 ) ;
  assign n3072 = n3051 ^ n2980 ^ 1'b0 ;
  assign n3073 = ( n2980 & n3021 ) | ( n2980 & ~n3072 ) | ( n3021 & ~n3072 ) ;
  assign n3074 = n3051 ^ n2942 ^ 1'b0 ;
  assign n3075 = ( n2942 & n3020 ) | ( n2942 & ~n3074 ) | ( n3020 & ~n3074 ) ;
  assign n3076 = n3051 ^ n2983 ^ 1'b0 ;
  assign n3077 = ( n2983 & n3019 ) | ( n2983 & ~n3076 ) | ( n3019 & ~n3076 ) ;
  assign n3078 = n3051 ^ n2986 ^ 1'b0 ;
  assign n3079 = ( n2986 & n3018 ) | ( n2986 & ~n3078 ) | ( n3018 & ~n3078 ) ;
  assign n3080 = n3051 ^ n2989 ^ 1'b0 ;
  assign n3081 = ( n2989 & n3017 ) | ( n2989 & ~n3080 ) | ( n3017 & ~n3080 ) ;
  assign n3082 = n3051 ^ n2997 ^ 1'b0 ;
  assign n3083 = ( n2997 & n3016 ) | ( n2997 & ~n3082 ) | ( n3016 & ~n3082 ) ;
  assign n3084 = n3051 ^ n2995 ^ 1'b0 ;
  assign n3085 = ( n2913 & n2995 ) | ( n2913 & n3084 ) | ( n2995 & n3084 ) ;
  assign n3086 = n3051 ^ n2993 ^ 1'b0 ;
  assign n3087 = ( n2941 & n2993 ) | ( n2941 & n3086 ) | ( n2993 & n3086 ) ;
  assign n3088 = n322 | n3050 ;
  assign n3089 = ( n322 & n3011 ) | ( n322 & n3088 ) | ( n3011 & n3088 ) ;
  assign n3090 = n3047 ^ n2945 ^ x98 ;
  assign n3091 = n3051 ^ n2945 ^ 1'b0 ;
  assign n3092 = ( n2945 & n3090 ) | ( n2945 & ~n3091 ) | ( n3090 & ~n3091 ) ;
  assign n3093 = n3045 ^ n2905 ^ x96 ;
  assign n3094 = n3051 ^ n2905 ^ 1'b0 ;
  assign n3095 = ( n2905 & n3093 ) | ( n2905 & ~n3094 ) | ( n3093 & ~n3094 ) ;
  assign n3096 = n3044 ^ n2936 ^ x95 ;
  assign n3097 = n3051 ^ n2936 ^ 1'b0 ;
  assign n3098 = ( n2936 & n3096 ) | ( n2936 & ~n3097 ) | ( n3096 & ~n3097 ) ;
  assign n3099 = n3043 ^ n2909 ^ x94 ;
  assign n3100 = n3051 ^ n2909 ^ 1'b0 ;
  assign n3101 = ( n2909 & n3099 ) | ( n2909 & ~n3100 ) | ( n3099 & ~n3100 ) ;
  assign n3102 = n3042 ^ n2902 ^ x93 ;
  assign n3103 = n3051 ^ n2902 ^ 1'b0 ;
  assign n3104 = ( n2902 & n3102 ) | ( n2902 & ~n3103 ) | ( n3102 & ~n3103 ) ;
  assign n3105 = n3041 ^ n2959 ^ x92 ;
  assign n3106 = n3051 ^ n2959 ^ 1'b0 ;
  assign n3107 = ( n2959 & n3105 ) | ( n2959 & ~n3106 ) | ( n3105 & ~n3106 ) ;
  assign n3108 = n3040 ^ n2916 ^ x91 ;
  assign n3109 = n3051 ^ n2916 ^ 1'b0 ;
  assign n3110 = ( n2916 & n3108 ) | ( n2916 & ~n3109 ) | ( n3108 & ~n3109 ) ;
  assign n3111 = n3039 ^ n2922 ^ x90 ;
  assign n3112 = n3051 ^ n2922 ^ 1'b0 ;
  assign n3113 = ( n2922 & n3111 ) | ( n2922 & ~n3112 ) | ( n3111 & ~n3112 ) ;
  assign n3114 = n3038 ^ n2949 ^ x89 ;
  assign n3115 = n3051 ^ n2949 ^ 1'b0 ;
  assign n3116 = ( n2949 & n3114 ) | ( n2949 & ~n3115 ) | ( n3114 & ~n3115 ) ;
  assign n3117 = n3051 ^ n2952 ^ 1'b0 ;
  assign n3118 = n3036 ^ n2955 ^ x87 ;
  assign n3119 = n3051 ^ n2955 ^ 1'b0 ;
  assign n3120 = ( n2955 & n3118 ) | ( n2955 & ~n3119 ) | ( n3118 & ~n3119 ) ;
  assign n3121 = n3035 ^ n2958 ^ x86 ;
  assign n3122 = n3051 ^ n2958 ^ 1'b0 ;
  assign n3123 = ( n2958 & n3121 ) | ( n2958 & ~n3122 ) | ( n3121 & ~n3122 ) ;
  assign n3124 = n3034 ^ n2934 ^ x85 ;
  assign n3125 = n3051 ^ n2934 ^ 1'b0 ;
  assign n3126 = ( n2934 & n3124 ) | ( n2934 & ~n3125 ) | ( n3124 & ~n3125 ) ;
  assign n3127 = n3037 ^ n2952 ^ x88 ;
  assign n3128 = ( n2952 & ~n3117 ) | ( n2952 & n3127 ) | ( ~n3117 & n3127 ) ;
  assign n3129 = n3033 ^ n2962 ^ x84 ;
  assign n3130 = n3051 ^ n2962 ^ 1'b0 ;
  assign n3131 = ( n2962 & n3129 ) | ( n2962 & ~n3130 ) | ( n3129 & ~n3130 ) ;
  assign n3132 = n3032 ^ n2965 ^ x83 ;
  assign n3133 = n3051 ^ n2965 ^ 1'b0 ;
  assign n3134 = ( n2965 & n3132 ) | ( n2965 & ~n3133 ) | ( n3132 & ~n3133 ) ;
  assign n3135 = n3014 ^ n2971 ^ x81 ;
  assign n3136 = n3051 ^ n2971 ^ 1'b0 ;
  assign n3137 = ( n2971 & n3135 ) | ( n2971 & ~n3136 ) | ( n3135 & ~n3136 ) ;
  assign n3138 = n3051 ^ n2974 ^ 1'b0 ;
  assign n3139 = ( n2974 & n3026 ) | ( n2974 & ~n3138 ) | ( n3026 & ~n3138 ) ;
  assign n3140 = ~x27 & x64 ;
  assign n3141 = x64 & n3051 ;
  assign n3142 = n3141 ^ x64 ^ x28 ;
  assign n3143 = n3142 ^ n3140 ^ x65 ;
  assign n3144 = ( x65 & n3140 ) | ( x65 & n3143 ) | ( n3140 & n3143 ) ;
  assign n3145 = n3144 ^ n3087 ^ x66 ;
  assign n3146 = ( x66 & n3144 ) | ( x66 & n3145 ) | ( n3144 & n3145 ) ;
  assign n3147 = ( x67 & ~n3085 ) | ( x67 & n3146 ) | ( ~n3085 & n3146 ) ;
  assign n3148 = ( x68 & ~n3083 ) | ( x68 & n3147 ) | ( ~n3083 & n3147 ) ;
  assign n3149 = ( x69 & ~n3081 ) | ( x69 & n3148 ) | ( ~n3081 & n3148 ) ;
  assign n3150 = ( x70 & ~n3079 ) | ( x70 & n3149 ) | ( ~n3079 & n3149 ) ;
  assign n3151 = ( x71 & ~n3077 ) | ( x71 & n3150 ) | ( ~n3077 & n3150 ) ;
  assign n3152 = ( x72 & ~n3075 ) | ( x72 & n3151 ) | ( ~n3075 & n3151 ) ;
  assign n3153 = ( x73 & ~n3073 ) | ( x73 & n3152 ) | ( ~n3073 & n3152 ) ;
  assign n3154 = ( x74 & ~n3071 ) | ( x74 & n3153 ) | ( ~n3071 & n3153 ) ;
  assign n3155 = ( x75 & ~n3069 ) | ( x75 & n3154 ) | ( ~n3069 & n3154 ) ;
  assign n3156 = ( x76 & ~n3067 ) | ( x76 & n3155 ) | ( ~n3067 & n3155 ) ;
  assign n3157 = ( x77 & ~n3065 ) | ( x77 & n3156 ) | ( ~n3065 & n3156 ) ;
  assign n3158 = ( x78 & ~n3139 ) | ( x78 & n3157 ) | ( ~n3139 & n3157 ) ;
  assign n3159 = ( x79 & ~n3063 ) | ( x79 & n3158 ) | ( ~n3063 & n3158 ) ;
  assign n3160 = ( x80 & ~n3061 ) | ( x80 & n3159 ) | ( ~n3061 & n3159 ) ;
  assign n3161 = ( x81 & ~n3059 ) | ( x81 & n3160 ) | ( ~n3059 & n3160 ) ;
  assign n3162 = ( x82 & ~n3137 ) | ( x82 & n3161 ) | ( ~n3137 & n3161 ) ;
  assign n3163 = ( x83 & ~n3057 ) | ( x83 & n3162 ) | ( ~n3057 & n3162 ) ;
  assign n3164 = ( x84 & ~n3134 ) | ( x84 & n3163 ) | ( ~n3134 & n3163 ) ;
  assign n3165 = ( x85 & ~n3131 ) | ( x85 & n3164 ) | ( ~n3131 & n3164 ) ;
  assign n3166 = ( x86 & ~n3126 ) | ( x86 & n3165 ) | ( ~n3126 & n3165 ) ;
  assign n3167 = ( x87 & ~n3123 ) | ( x87 & n3166 ) | ( ~n3123 & n3166 ) ;
  assign n3168 = ( x88 & ~n3120 ) | ( x88 & n3167 ) | ( ~n3120 & n3167 ) ;
  assign n3169 = ( x89 & ~n3128 ) | ( x89 & n3168 ) | ( ~n3128 & n3168 ) ;
  assign n3170 = ( x90 & ~n3116 ) | ( x90 & n3169 ) | ( ~n3116 & n3169 ) ;
  assign n3171 = ( x91 & ~n3113 ) | ( x91 & n3170 ) | ( ~n3113 & n3170 ) ;
  assign n3172 = ( x92 & ~n3110 ) | ( x92 & n3171 ) | ( ~n3110 & n3171 ) ;
  assign n3173 = ( x93 & ~n3107 ) | ( x93 & n3172 ) | ( ~n3107 & n3172 ) ;
  assign n3174 = ( x94 & ~n3104 ) | ( x94 & n3173 ) | ( ~n3104 & n3173 ) ;
  assign n3175 = ( x95 & ~n3101 ) | ( x95 & n3174 ) | ( ~n3101 & n3174 ) ;
  assign n3176 = ( x96 & ~n3098 ) | ( x96 & n3175 ) | ( ~n3098 & n3175 ) ;
  assign n3177 = ( x97 & ~n3095 ) | ( x97 & n3176 ) | ( ~n3095 & n3176 ) ;
  assign n3178 = ( x98 & ~n3054 ) | ( x98 & n3177 ) | ( ~n3054 & n3177 ) ;
  assign n3179 = n3178 ^ n3092 ^ x99 ;
  assign n3180 = ( x99 & ~n3092 ) | ( x99 & n3178 ) | ( ~n3092 & n3178 ) ;
  assign n3181 = ( x100 & ~n3089 ) | ( x100 & n3180 ) | ( ~n3089 & n3180 ) ;
  assign n3182 = n168 | n3181 ;
  assign n3183 = n3182 ^ n3092 ^ 1'b0 ;
  assign n3184 = ( n3092 & n3179 ) | ( n3092 & ~n3183 ) | ( n3179 & ~n3183 ) ;
  assign n3185 = n3177 ^ n3054 ^ x98 ;
  assign n3186 = n3182 ^ n3054 ^ 1'b0 ;
  assign n3187 = ( n3054 & n3185 ) | ( n3054 & ~n3186 ) | ( n3185 & ~n3186 ) ;
  assign n3188 = n3176 ^ n3095 ^ x97 ;
  assign n3189 = n3182 ^ n3095 ^ 1'b0 ;
  assign n3190 = ( n3095 & n3188 ) | ( n3095 & ~n3189 ) | ( n3188 & ~n3189 ) ;
  assign n3191 = n3175 ^ n3098 ^ x96 ;
  assign n3192 = n3182 ^ n3098 ^ 1'b0 ;
  assign n3193 = ( n3098 & n3191 ) | ( n3098 & ~n3192 ) | ( n3191 & ~n3192 ) ;
  assign n3194 = n3172 ^ n3107 ^ x93 ;
  assign n3195 = n3182 ^ n3107 ^ 1'b0 ;
  assign n3196 = ( n3107 & n3194 ) | ( n3107 & ~n3195 ) | ( n3194 & ~n3195 ) ;
  assign n3197 = n3153 ^ n3071 ^ x74 ;
  assign n3198 = n3182 ^ n3071 ^ 1'b0 ;
  assign n3199 = ( n3071 & n3197 ) | ( n3071 & ~n3198 ) | ( n3197 & ~n3198 ) ;
  assign n3200 = n3151 ^ n3075 ^ x72 ;
  assign n3201 = n3182 ^ n3075 ^ 1'b0 ;
  assign n3202 = ( n3075 & n3200 ) | ( n3075 & ~n3201 ) | ( n3200 & ~n3201 ) ;
  assign n3203 = n3149 ^ n3079 ^ x70 ;
  assign n3204 = n3182 ^ n3079 ^ 1'b0 ;
  assign n3205 = ( n3079 & n3203 ) | ( n3079 & ~n3204 ) | ( n3203 & ~n3204 ) ;
  assign n3206 = n3146 ^ n3085 ^ x67 ;
  assign n3207 = n3182 ^ n3085 ^ 1'b0 ;
  assign n3208 = ( n3085 & n3206 ) | ( n3085 & ~n3207 ) | ( n3206 & ~n3207 ) ;
  assign n3209 = n3182 ^ n3145 ^ 1'b0 ;
  assign n3210 = ( n3087 & n3145 ) | ( n3087 & n3209 ) | ( n3145 & n3209 ) ;
  assign n3211 = n3182 ^ n3143 ^ 1'b0 ;
  assign n3212 = ( n3142 & n3143 ) | ( n3142 & n3211 ) | ( n3143 & n3211 ) ;
  assign n3213 = n3174 ^ n3101 ^ x95 ;
  assign n3214 = n3182 ^ n3101 ^ 1'b0 ;
  assign n3215 = ( n3101 & n3213 ) | ( n3101 & ~n3214 ) | ( n3213 & ~n3214 ) ;
  assign n3216 = n3173 ^ n3104 ^ x94 ;
  assign n3217 = n3182 ^ n3104 ^ 1'b0 ;
  assign n3218 = ( n3104 & n3216 ) | ( n3104 & ~n3217 ) | ( n3216 & ~n3217 ) ;
  assign n3219 = n3171 ^ n3110 ^ x92 ;
  assign n3220 = n3182 ^ n3110 ^ 1'b0 ;
  assign n3221 = ( n3110 & n3219 ) | ( n3110 & ~n3220 ) | ( n3219 & ~n3220 ) ;
  assign n3222 = n3169 ^ n3116 ^ x90 ;
  assign n3223 = n3182 ^ n3116 ^ 1'b0 ;
  assign n3224 = ( n3116 & n3222 ) | ( n3116 & ~n3223 ) | ( n3222 & ~n3223 ) ;
  assign n3225 = n3168 ^ n3128 ^ x89 ;
  assign n3226 = n3182 ^ n3128 ^ 1'b0 ;
  assign n3227 = ( n3128 & n3225 ) | ( n3128 & ~n3226 ) | ( n3225 & ~n3226 ) ;
  assign n3228 = n3167 ^ n3120 ^ x88 ;
  assign n3229 = n3182 ^ n3120 ^ 1'b0 ;
  assign n3230 = ( n3120 & n3228 ) | ( n3120 & ~n3229 ) | ( n3228 & ~n3229 ) ;
  assign n3231 = n3166 ^ n3123 ^ x87 ;
  assign n3232 = n3182 ^ n3123 ^ 1'b0 ;
  assign n3233 = ( n3123 & n3231 ) | ( n3123 & ~n3232 ) | ( n3231 & ~n3232 ) ;
  assign n3234 = n3165 ^ n3126 ^ x86 ;
  assign n3235 = n3182 ^ n3126 ^ 1'b0 ;
  assign n3236 = ( n3126 & n3234 ) | ( n3126 & ~n3235 ) | ( n3234 & ~n3235 ) ;
  assign n3237 = n3164 ^ n3131 ^ x85 ;
  assign n3238 = n3182 ^ n3131 ^ 1'b0 ;
  assign n3239 = ( n3131 & n3237 ) | ( n3131 & ~n3238 ) | ( n3237 & ~n3238 ) ;
  assign n3240 = n3163 ^ n3134 ^ x84 ;
  assign n3241 = n3182 ^ n3134 ^ 1'b0 ;
  assign n3242 = ( n3134 & n3240 ) | ( n3134 & ~n3241 ) | ( n3240 & ~n3241 ) ;
  assign n3243 = n3161 ^ n3137 ^ x82 ;
  assign n3244 = n3182 ^ n3137 ^ 1'b0 ;
  assign n3245 = ( n3137 & n3243 ) | ( n3137 & ~n3244 ) | ( n3243 & ~n3244 ) ;
  assign n3246 = n3160 ^ n3059 ^ x81 ;
  assign n3247 = n3182 ^ n3059 ^ 1'b0 ;
  assign n3248 = ( n3059 & n3246 ) | ( n3059 & ~n3247 ) | ( n3246 & ~n3247 ) ;
  assign n3249 = n3159 ^ n3061 ^ x80 ;
  assign n3250 = n3182 ^ n3061 ^ 1'b0 ;
  assign n3251 = ( n3061 & n3249 ) | ( n3061 & ~n3250 ) | ( n3249 & ~n3250 ) ;
  assign n3252 = n3156 ^ n3065 ^ x77 ;
  assign n3253 = n3182 ^ n3065 ^ 1'b0 ;
  assign n3254 = ( n3065 & n3252 ) | ( n3065 & ~n3253 ) | ( n3252 & ~n3253 ) ;
  assign n3255 = n3155 ^ n3067 ^ x76 ;
  assign n3256 = n3182 ^ n3067 ^ 1'b0 ;
  assign n3257 = ( n3067 & n3255 ) | ( n3067 & ~n3256 ) | ( n3255 & ~n3256 ) ;
  assign n3258 = n3154 ^ n3069 ^ x75 ;
  assign n3259 = n3182 ^ n3069 ^ 1'b0 ;
  assign n3260 = ( n3069 & n3258 ) | ( n3069 & ~n3259 ) | ( n3258 & ~n3259 ) ;
  assign n3261 = n3152 ^ n3073 ^ x73 ;
  assign n3262 = n3182 ^ n3073 ^ 1'b0 ;
  assign n3263 = ( n3073 & n3261 ) | ( n3073 & ~n3262 ) | ( n3261 & ~n3262 ) ;
  assign n3264 = n3150 ^ n3077 ^ x71 ;
  assign n3265 = n3182 ^ n3077 ^ 1'b0 ;
  assign n3266 = ( n3077 & n3264 ) | ( n3077 & ~n3265 ) | ( n3264 & ~n3265 ) ;
  assign n3267 = n3148 ^ n3081 ^ x69 ;
  assign n3268 = n3182 ^ n3081 ^ 1'b0 ;
  assign n3269 = ( n3081 & n3267 ) | ( n3081 & ~n3268 ) | ( n3267 & ~n3268 ) ;
  assign n3270 = n3147 ^ n3083 ^ x68 ;
  assign n3271 = n3182 ^ n3083 ^ 1'b0 ;
  assign n3272 = ( n3083 & n3270 ) | ( n3083 & ~n3271 ) | ( n3270 & ~n3271 ) ;
  assign n3273 = n183 | n193 ;
  assign n3274 = ( ~x102 & x103 ) | ( ~x102 & n189 ) | ( x103 & n189 ) ;
  assign n3275 = x102 | n3274 ;
  assign n3276 = n3170 ^ n3113 ^ x91 ;
  assign n3277 = n3273 | n3275 ;
  assign n3278 = x27 & x64 ;
  assign n3279 = x101 | n3181 ;
  assign n3280 = ( n3277 & n3278 ) | ( n3277 & ~n3279 ) | ( n3278 & ~n3279 ) ;
  assign n3281 = n3182 ^ n3057 ^ 1'b0 ;
  assign n3282 = n3157 ^ n3139 ^ x78 ;
  assign n3283 = n3182 ^ n3113 ^ 1'b0 ;
  assign n3284 = ~n3277 & n3280 ;
  assign n3285 = n3140 & ~n3182 ;
  assign n3286 = ( x27 & ~n3284 ) | ( x27 & n3285 ) | ( ~n3284 & n3285 ) ;
  assign n3287 = n3158 ^ n3063 ^ x79 ;
  assign n3288 = ~x26 & x64 ;
  assign n3289 = n3288 ^ n3286 ^ x65 ;
  assign n3290 = ( x65 & n3288 ) | ( x65 & n3289 ) | ( n3288 & n3289 ) ;
  assign n3291 = n3290 ^ n3212 ^ x66 ;
  assign n3292 = ( x66 & n3290 ) | ( x66 & n3291 ) | ( n3290 & n3291 ) ;
  assign n3293 = ( x67 & ~n3210 ) | ( x67 & n3292 ) | ( ~n3210 & n3292 ) ;
  assign n3294 = ( x68 & ~n3208 ) | ( x68 & n3293 ) | ( ~n3208 & n3293 ) ;
  assign n3295 = n3162 ^ n3057 ^ x83 ;
  assign n3296 = n3182 ^ n3139 ^ 1'b0 ;
  assign n3297 = ( x69 & ~n3272 ) | ( x69 & n3294 ) | ( ~n3272 & n3294 ) ;
  assign n3298 = ( x70 & ~n3269 ) | ( x70 & n3297 ) | ( ~n3269 & n3297 ) ;
  assign n3299 = ~n3273 & n3288 ;
  assign n3300 = ( x71 & ~n3205 ) | ( x71 & n3298 ) | ( ~n3205 & n3298 ) ;
  assign n3301 = ( x72 & ~n3266 ) | ( x72 & n3300 ) | ( ~n3266 & n3300 ) ;
  assign n3302 = ( x73 & ~n3202 ) | ( x73 & n3301 ) | ( ~n3202 & n3301 ) ;
  assign n3303 = ( x74 & ~n3263 ) | ( x74 & n3302 ) | ( ~n3263 & n3302 ) ;
  assign n3304 = n3293 ^ n3208 ^ x68 ;
  assign n3305 = n3294 ^ n3272 ^ x69 ;
  assign n3306 = ( x75 & ~n3199 ) | ( x75 & n3303 ) | ( ~n3199 & n3303 ) ;
  assign n3307 = ( x76 & ~n3260 ) | ( x76 & n3306 ) | ( ~n3260 & n3306 ) ;
  assign n3308 = ( x77 & ~n3257 ) | ( x77 & n3307 ) | ( ~n3257 & n3307 ) ;
  assign n3309 = ( n3139 & n3282 ) | ( n3139 & ~n3296 ) | ( n3282 & ~n3296 ) ;
  assign n3310 = ( x78 & ~n3254 ) | ( x78 & n3308 ) | ( ~n3254 & n3308 ) ;
  assign n3311 = ( x79 & ~n3309 ) | ( x79 & n3310 ) | ( ~n3309 & n3310 ) ;
  assign n3312 = n3182 ^ n3063 ^ 1'b0 ;
  assign n3313 = ( n322 & n3089 ) | ( n322 & n3182 ) | ( n3089 & n3182 ) ;
  assign n3314 = ( n3063 & n3287 ) | ( n3063 & ~n3312 ) | ( n3287 & ~n3312 ) ;
  assign n3315 = ( x80 & n3311 ) | ( x80 & ~n3314 ) | ( n3311 & ~n3314 ) ;
  assign n3316 = ( x81 & ~n3251 ) | ( x81 & n3315 ) | ( ~n3251 & n3315 ) ;
  assign n3317 = ( n3057 & ~n3281 ) | ( n3057 & n3295 ) | ( ~n3281 & n3295 ) ;
  assign n3318 = ( x82 & ~n3248 ) | ( x82 & n3316 ) | ( ~n3248 & n3316 ) ;
  assign n3319 = ( x83 & ~n3245 ) | ( x83 & n3318 ) | ( ~n3245 & n3318 ) ;
  assign n3320 = ( n3113 & n3276 ) | ( n3113 & ~n3283 ) | ( n3276 & ~n3283 ) ;
  assign n3321 = ( x84 & ~n3317 ) | ( x84 & n3319 ) | ( ~n3317 & n3319 ) ;
  assign n3322 = ( x85 & ~n3242 ) | ( x85 & n3321 ) | ( ~n3242 & n3321 ) ;
  assign n3323 = ( x86 & ~n3239 ) | ( x86 & n3322 ) | ( ~n3239 & n3322 ) ;
  assign n3324 = ( x87 & ~n3236 ) | ( x87 & n3323 ) | ( ~n3236 & n3323 ) ;
  assign n3325 = ( x88 & ~n3233 ) | ( x88 & n3324 ) | ( ~n3233 & n3324 ) ;
  assign n3326 = ( x89 & ~n3230 ) | ( x89 & n3325 ) | ( ~n3230 & n3325 ) ;
  assign n3327 = ( x90 & ~n3227 ) | ( x90 & n3326 ) | ( ~n3227 & n3326 ) ;
  assign n3328 = ( x91 & ~n3224 ) | ( x91 & n3327 ) | ( ~n3224 & n3327 ) ;
  assign n3329 = ( x92 & ~n3320 ) | ( x92 & n3328 ) | ( ~n3320 & n3328 ) ;
  assign n3330 = ( x93 & ~n3221 ) | ( x93 & n3329 ) | ( ~n3221 & n3329 ) ;
  assign n3331 = ( x94 & ~n3196 ) | ( x94 & n3330 ) | ( ~n3196 & n3330 ) ;
  assign n3332 = ( x95 & ~n3218 ) | ( x95 & n3331 ) | ( ~n3218 & n3331 ) ;
  assign n3333 = ( x96 & ~n3215 ) | ( x96 & n3332 ) | ( ~n3215 & n3332 ) ;
  assign n3334 = ( x97 & ~n3193 ) | ( x97 & n3333 ) | ( ~n3193 & n3333 ) ;
  assign n3335 = n3326 ^ n3227 ^ x90 ;
  assign n3336 = ( x98 & ~n3190 ) | ( x98 & n3334 ) | ( ~n3190 & n3334 ) ;
  assign n3337 = ( x99 & ~n3187 ) | ( x99 & n3336 ) | ( ~n3187 & n3336 ) ;
  assign n3338 = ( x100 & ~n3184 ) | ( x100 & n3337 ) | ( ~n3184 & n3337 ) ;
  assign n3339 = ( x101 & ~n3313 ) | ( x101 & n3338 ) | ( ~n3313 & n3338 ) ;
  assign n3340 = n3277 | n3339 ;
  assign n3341 = n3327 ^ n3224 ^ x91 ;
  assign n3342 = n3333 ^ n3193 ^ x97 ;
  assign n3343 = ( ~n3275 & n3299 ) | ( ~n3275 & n3339 ) | ( n3299 & n3339 ) ;
  assign n3344 = n3340 ^ n3291 ^ 1'b0 ;
  assign n3345 = n3337 ^ n3184 ^ x100 ;
  assign n3346 = n3328 ^ n3320 ^ x92 ;
  assign n3347 = n3330 ^ n3196 ^ x94 ;
  assign n3348 = ( n3212 & n3291 ) | ( n3212 & n3344 ) | ( n3291 & n3344 ) ;
  assign n3349 = n3340 ^ n3218 ^ 1'b0 ;
  assign n3350 = n3340 ^ n3196 ^ 1'b0 ;
  assign n3351 = ( n3196 & n3347 ) | ( n3196 & ~n3350 ) | ( n3347 & ~n3350 ) ;
  assign n3352 = n3345 ^ n3340 ^ 1'b0 ;
  assign n3353 = n3340 ^ n3227 ^ 1'b0 ;
  assign n3354 = n3332 ^ n3215 ^ x96 ;
  assign n3355 = ( n3227 & n3335 ) | ( n3227 & ~n3353 ) | ( n3335 & ~n3353 ) ;
  assign n3356 = n3340 ^ n3193 ^ 1'b0 ;
  assign n3357 = n3340 ^ n3208 ^ 1'b0 ;
  assign n3358 = ( n3208 & n3304 ) | ( n3208 & ~n3357 ) | ( n3304 & ~n3357 ) ;
  assign n3359 = n3340 ^ n3224 ^ 1'b0 ;
  assign n3360 = n3329 ^ n3221 ^ x93 ;
  assign n3361 = n3331 ^ n3218 ^ x95 ;
  assign n3362 = n3336 ^ n3187 ^ x99 ;
  assign n3363 = n3340 ^ n3187 ^ 1'b0 ;
  assign n3364 = ( n3224 & n3341 ) | ( n3224 & ~n3359 ) | ( n3341 & ~n3359 ) ;
  assign n3365 = n3340 ^ n3215 ^ 1'b0 ;
  assign n3366 = n3340 ^ n3190 ^ 1'b0 ;
  assign n3367 = ( n3218 & ~n3349 ) | ( n3218 & n3361 ) | ( ~n3349 & n3361 ) ;
  assign n3368 = n3340 ^ n3272 ^ 1'b0 ;
  assign n3369 = n3340 ^ n3221 ^ 1'b0 ;
  assign n3370 = n3334 ^ n3190 ^ x98 ;
  assign n3371 = ( n3193 & n3342 ) | ( n3193 & ~n3356 ) | ( n3342 & ~n3356 ) ;
  assign n3372 = ( n3187 & n3362 ) | ( n3187 & ~n3363 ) | ( n3362 & ~n3363 ) ;
  assign n3373 = ( n3221 & n3360 ) | ( n3221 & ~n3369 ) | ( n3360 & ~n3369 ) ;
  assign n3374 = n3340 ^ n3289 ^ 1'b0 ;
  assign n3375 = ( n3286 & n3289 ) | ( n3286 & n3374 ) | ( n3289 & n3374 ) ;
  assign n3376 = ( n3272 & n3305 ) | ( n3272 & ~n3368 ) | ( n3305 & ~n3368 ) ;
  assign n3377 = ( n3190 & ~n3366 ) | ( n3190 & n3370 ) | ( ~n3366 & n3370 ) ;
  assign n3378 = n3340 ^ n3320 ^ 1'b0 ;
  assign n3379 = ( n3215 & n3354 ) | ( n3215 & ~n3365 ) | ( n3354 & ~n3365 ) ;
  assign n3380 = ( n3320 & n3346 ) | ( n3320 & ~n3378 ) | ( n3346 & ~n3378 ) ;
  assign n3381 = ( n3184 & n3345 ) | ( n3184 & n3352 ) | ( n3345 & n3352 ) ;
  assign n3382 = n3325 ^ n3230 ^ x89 ;
  assign n3383 = n3340 ^ n3230 ^ 1'b0 ;
  assign n3384 = ( n3230 & n3382 ) | ( n3230 & ~n3383 ) | ( n3382 & ~n3383 ) ;
  assign n3385 = n3324 ^ n3233 ^ x88 ;
  assign n3386 = n3340 ^ n3233 ^ 1'b0 ;
  assign n3387 = ( n3233 & n3385 ) | ( n3233 & ~n3386 ) | ( n3385 & ~n3386 ) ;
  assign n3388 = n3316 ^ n3248 ^ x82 ;
  assign n3389 = n3340 ^ n3248 ^ 1'b0 ;
  assign n3390 = ( n3248 & n3388 ) | ( n3248 & ~n3389 ) | ( n3388 & ~n3389 ) ;
  assign n3391 = n3315 ^ n3251 ^ x81 ;
  assign n3392 = n3340 ^ n3251 ^ 1'b0 ;
  assign n3393 = ( n3251 & n3391 ) | ( n3251 & ~n3392 ) | ( n3391 & ~n3392 ) ;
  assign n3394 = n3314 ^ n3311 ^ x80 ;
  assign n3395 = n3340 ^ n3314 ^ 1'b0 ;
  assign n3396 = ( n3314 & n3394 ) | ( n3314 & ~n3395 ) | ( n3394 & ~n3395 ) ;
  assign n3397 = n3310 ^ n3309 ^ x79 ;
  assign n3398 = n3340 ^ n3309 ^ 1'b0 ;
  assign n3399 = ( n3309 & n3397 ) | ( n3309 & ~n3398 ) | ( n3397 & ~n3398 ) ;
  assign n3400 = n3340 ^ n3254 ^ 1'b0 ;
  assign n3401 = n3307 ^ n3257 ^ x77 ;
  assign n3402 = n3340 ^ n3257 ^ 1'b0 ;
  assign n3403 = ( n3257 & n3401 ) | ( n3257 & ~n3402 ) | ( n3401 & ~n3402 ) ;
  assign n3404 = n3306 ^ n3260 ^ x76 ;
  assign n3405 = n3340 ^ n3260 ^ 1'b0 ;
  assign n3406 = n3308 ^ n3254 ^ x78 ;
  assign n3407 = ( n3254 & ~n3400 ) | ( n3254 & n3406 ) | ( ~n3400 & n3406 ) ;
  assign n3408 = ( n3260 & n3404 ) | ( n3260 & ~n3405 ) | ( n3404 & ~n3405 ) ;
  assign n3409 = n3303 ^ n3199 ^ x75 ;
  assign n3410 = n3340 ^ n3199 ^ 1'b0 ;
  assign n3411 = ( n3199 & n3409 ) | ( n3199 & ~n3410 ) | ( n3409 & ~n3410 ) ;
  assign n3412 = n3302 ^ n3263 ^ x74 ;
  assign n3413 = n3340 ^ n3263 ^ 1'b0 ;
  assign n3414 = ( n3263 & n3412 ) | ( n3263 & ~n3413 ) | ( n3412 & ~n3413 ) ;
  assign n3415 = n3301 ^ n3202 ^ x73 ;
  assign n3416 = n3340 ^ n3202 ^ 1'b0 ;
  assign n3417 = ( n3202 & n3415 ) | ( n3202 & ~n3416 ) | ( n3415 & ~n3416 ) ;
  assign n3418 = n3300 ^ n3266 ^ x72 ;
  assign n3419 = n3340 ^ n3266 ^ 1'b0 ;
  assign n3420 = ( n3266 & n3418 ) | ( n3266 & ~n3419 ) | ( n3418 & ~n3419 ) ;
  assign n3421 = n3298 ^ n3205 ^ x71 ;
  assign n3422 = n3340 ^ n3205 ^ 1'b0 ;
  assign n3423 = ( n3205 & n3421 ) | ( n3205 & ~n3422 ) | ( n3421 & ~n3422 ) ;
  assign n3424 = n3297 ^ n3269 ^ x70 ;
  assign n3425 = n3340 ^ n3269 ^ 1'b0 ;
  assign n3426 = ( n3269 & n3424 ) | ( n3269 & ~n3425 ) | ( n3424 & ~n3425 ) ;
  assign n3427 = n3292 ^ n3210 ^ x67 ;
  assign n3428 = n3340 ^ n3210 ^ 1'b0 ;
  assign n3429 = ( n3210 & n3427 ) | ( n3210 & ~n3428 ) | ( n3427 & ~n3428 ) ;
  assign n3430 = x26 & x64 ;
  assign n3431 = ( ~x102 & n3339 ) | ( ~x102 & n3430 ) | ( n3339 & n3430 ) ;
  assign n3432 = ~n3339 & n3431 ;
  assign n3433 = ~n3339 & n3343 ;
  assign n3434 = ~x25 & x64 ;
  assign n3435 = ( ~n176 & n1297 ) | ( ~n176 & n3432 ) | ( n1297 & n3432 ) ;
  assign n3436 = n3313 & n3340 ;
  assign n3437 = n322 | n3436 ;
  assign n3438 = ~n1297 & n3435 ;
  assign n3439 = n3321 ^ n3242 ^ x85 ;
  assign n3440 = ( x26 & n3433 ) | ( x26 & ~n3438 ) | ( n3433 & ~n3438 ) ;
  assign n3441 = n3340 ^ n3242 ^ 1'b0 ;
  assign n3442 = ( n3242 & n3439 ) | ( n3242 & ~n3441 ) | ( n3439 & ~n3441 ) ;
  assign n3443 = n3340 ^ n3245 ^ 1'b0 ;
  assign n3444 = n3318 ^ n3245 ^ x83 ;
  assign n3445 = ( n3245 & ~n3443 ) | ( n3245 & n3444 ) | ( ~n3443 & n3444 ) ;
  assign n3446 = n3440 ^ n3434 ^ x65 ;
  assign n3447 = ( n322 & n3277 ) | ( n322 & n3313 ) | ( n3277 & n3313 ) ;
  assign n3448 = ( ~x102 & n1297 ) | ( ~x102 & n3437 ) | ( n1297 & n3437 ) ;
  assign n3449 = ( x65 & n3434 ) | ( x65 & n3446 ) | ( n3434 & n3446 ) ;
  assign n3450 = ( x102 & n1297 ) | ( x102 & ~n3436 ) | ( n1297 & ~n3436 ) ;
  assign n3451 = n3449 ^ n3375 ^ x66 ;
  assign n3452 = ( x66 & n3449 ) | ( x66 & n3451 ) | ( n3449 & n3451 ) ;
  assign n3453 = ( ~n176 & n3448 ) | ( ~n176 & n3450 ) | ( n3448 & n3450 ) ;
  assign n3454 = n3322 ^ n3239 ^ x86 ;
  assign n3455 = ( x67 & ~n3348 ) | ( x67 & n3452 ) | ( ~n3348 & n3452 ) ;
  assign n3456 = n3277 & n3437 ;
  assign n3457 = n3452 ^ n3348 ^ x67 ;
  assign n3458 = n3340 ^ n3317 ^ 1'b0 ;
  assign n3459 = n3323 ^ n3236 ^ x87 ;
  assign n3460 = n3319 ^ n3317 ^ x84 ;
  assign n3461 = ( n3317 & ~n3458 ) | ( n3317 & n3460 ) | ( ~n3458 & n3460 ) ;
  assign n3462 = n3340 ^ n3239 ^ 1'b0 ;
  assign n3463 = ( x68 & ~n3429 ) | ( x68 & n3455 ) | ( ~n3429 & n3455 ) ;
  assign n3464 = n3455 ^ n3429 ^ x68 ;
  assign n3465 = ( n3239 & n3454 ) | ( n3239 & ~n3462 ) | ( n3454 & ~n3462 ) ;
  assign n3466 = n3463 ^ n3358 ^ x69 ;
  assign n3467 = n3340 ^ n3236 ^ 1'b0 ;
  assign n3468 = ( x69 & ~n3358 ) | ( x69 & n3463 ) | ( ~n3358 & n3463 ) ;
  assign n3469 = ( n3236 & n3459 ) | ( n3236 & ~n3467 ) | ( n3459 & ~n3467 ) ;
  assign n3470 = n3468 ^ n3376 ^ x70 ;
  assign n3471 = ( x70 & ~n3376 ) | ( x70 & n3468 ) | ( ~n3376 & n3468 ) ;
  assign n3472 = ( x71 & ~n3426 ) | ( x71 & n3471 ) | ( ~n3426 & n3471 ) ;
  assign n3473 = n3471 ^ n3426 ^ x71 ;
  assign n3474 = ( x72 & ~n3423 ) | ( x72 & n3472 ) | ( ~n3423 & n3472 ) ;
  assign n3475 = ( x73 & ~n3420 ) | ( x73 & n3474 ) | ( ~n3420 & n3474 ) ;
  assign n3476 = ( x74 & ~n3417 ) | ( x74 & n3475 ) | ( ~n3417 & n3475 ) ;
  assign n3477 = ( x75 & ~n3414 ) | ( x75 & n3476 ) | ( ~n3414 & n3476 ) ;
  assign n3478 = ( x76 & ~n3411 ) | ( x76 & n3477 ) | ( ~n3411 & n3477 ) ;
  assign n3479 = ( x77 & ~n3408 ) | ( x77 & n3478 ) | ( ~n3408 & n3478 ) ;
  assign n3480 = ( x78 & ~n3403 ) | ( x78 & n3479 ) | ( ~n3403 & n3479 ) ;
  assign n3481 = ( x79 & ~n3407 ) | ( x79 & n3480 ) | ( ~n3407 & n3480 ) ;
  assign n3482 = ( x80 & ~n3399 ) | ( x80 & n3481 ) | ( ~n3399 & n3481 ) ;
  assign n3483 = ( x81 & ~n3396 ) | ( x81 & n3482 ) | ( ~n3396 & n3482 ) ;
  assign n3484 = ( x82 & ~n3393 ) | ( x82 & n3483 ) | ( ~n3393 & n3483 ) ;
  assign n3485 = ( x83 & ~n3390 ) | ( x83 & n3484 ) | ( ~n3390 & n3484 ) ;
  assign n3486 = ( x84 & ~n3445 ) | ( x84 & n3485 ) | ( ~n3445 & n3485 ) ;
  assign n3487 = ( x85 & ~n3461 ) | ( x85 & n3486 ) | ( ~n3461 & n3486 ) ;
  assign n3488 = ( x86 & ~n3442 ) | ( x86 & n3487 ) | ( ~n3442 & n3487 ) ;
  assign n3489 = ( x87 & ~n3465 ) | ( x87 & n3488 ) | ( ~n3465 & n3488 ) ;
  assign n3490 = ( x88 & ~n3469 ) | ( x88 & n3489 ) | ( ~n3469 & n3489 ) ;
  assign n3491 = ( x89 & ~n3387 ) | ( x89 & n3490 ) | ( ~n3387 & n3490 ) ;
  assign n3492 = ( x90 & ~n3384 ) | ( x90 & n3491 ) | ( ~n3384 & n3491 ) ;
  assign n3493 = ( x91 & ~n3355 ) | ( x91 & n3492 ) | ( ~n3355 & n3492 ) ;
  assign n3494 = ( x92 & ~n3364 ) | ( x92 & n3493 ) | ( ~n3364 & n3493 ) ;
  assign n3495 = ( x93 & ~n3380 ) | ( x93 & n3494 ) | ( ~n3380 & n3494 ) ;
  assign n3496 = ( x94 & ~n3373 ) | ( x94 & n3495 ) | ( ~n3373 & n3495 ) ;
  assign n3497 = ( x95 & ~n3351 ) | ( x95 & n3496 ) | ( ~n3351 & n3496 ) ;
  assign n3498 = ( x96 & ~n3367 ) | ( x96 & n3497 ) | ( ~n3367 & n3497 ) ;
  assign n3499 = ( x97 & ~n3379 ) | ( x97 & n3498 ) | ( ~n3379 & n3498 ) ;
  assign n3500 = ( x98 & ~n3371 ) | ( x98 & n3499 ) | ( ~n3371 & n3499 ) ;
  assign n3501 = ( x99 & ~n3377 ) | ( x99 & n3500 ) | ( ~n3377 & n3500 ) ;
  assign n3502 = ( x100 & ~n3372 ) | ( x100 & n3501 ) | ( ~n3372 & n3501 ) ;
  assign n3503 = ( x101 & ~n3381 ) | ( x101 & n3502 ) | ( ~n3381 & n3502 ) ;
  assign n3504 = ( ~n176 & n3453 ) | ( ~n176 & n3503 ) | ( n3453 & n3503 ) ;
  assign n3505 = n176 | n3504 ;
  assign n3506 = ( ~n3437 & n3456 ) | ( ~n3437 & n3505 ) | ( n3456 & n3505 ) ;
  assign n3507 = n3493 ^ n3364 ^ x92 ;
  assign n3508 = n3506 ^ n3364 ^ 1'b0 ;
  assign n3509 = ( n3364 & n3507 ) | ( n3364 & ~n3508 ) | ( n3507 & ~n3508 ) ;
  assign n3510 = n3490 ^ n3387 ^ x89 ;
  assign n3511 = n3484 ^ n3390 ^ x83 ;
  assign n3512 = n3506 ^ n3390 ^ 1'b0 ;
  assign n3513 = ( n3390 & n3511 ) | ( n3390 & ~n3512 ) | ( n3511 & ~n3512 ) ;
  assign n3514 = n3479 ^ n3403 ^ x78 ;
  assign n3515 = n3506 ^ n3403 ^ 1'b0 ;
  assign n3516 = ( n3403 & n3514 ) | ( n3403 & ~n3515 ) | ( n3514 & ~n3515 ) ;
  assign n3517 = n3478 ^ n3408 ^ x77 ;
  assign n3518 = n3506 ^ n3408 ^ 1'b0 ;
  assign n3519 = ( n3408 & n3517 ) | ( n3408 & ~n3518 ) | ( n3517 & ~n3518 ) ;
  assign n3520 = n3476 ^ n3414 ^ x75 ;
  assign n3521 = n3506 ^ n3414 ^ 1'b0 ;
  assign n3522 = ( n3414 & n3520 ) | ( n3414 & ~n3521 ) | ( n3520 & ~n3521 ) ;
  assign n3523 = n3506 ^ n3426 ^ 1'b0 ;
  assign n3524 = ( n3426 & n3473 ) | ( n3426 & ~n3523 ) | ( n3473 & ~n3523 ) ;
  assign n3525 = n3506 ^ n3376 ^ 1'b0 ;
  assign n3526 = ( n3376 & n3470 ) | ( n3376 & ~n3525 ) | ( n3470 & ~n3525 ) ;
  assign n3527 = n3506 ^ n3358 ^ 1'b0 ;
  assign n3528 = ( n3358 & n3466 ) | ( n3358 & ~n3527 ) | ( n3466 & ~n3527 ) ;
  assign n3529 = n3506 ^ n3429 ^ 1'b0 ;
  assign n3530 = ( n3429 & n3464 ) | ( n3429 & ~n3529 ) | ( n3464 & ~n3529 ) ;
  assign n3531 = n3506 ^ n3348 ^ 1'b0 ;
  assign n3532 = ( n3348 & n3457 ) | ( n3348 & ~n3531 ) | ( n3457 & ~n3531 ) ;
  assign n3533 = n322 | n3505 ;
  assign n3534 = ( n322 & n3447 ) | ( n322 & n3533 ) | ( n3447 & n3533 ) ;
  assign n3535 = n3497 ^ n3367 ^ x96 ;
  assign n3536 = n3506 ^ n3367 ^ 1'b0 ;
  assign n3537 = ( n3367 & n3535 ) | ( n3367 & ~n3536 ) | ( n3535 & ~n3536 ) ;
  assign n3538 = n3496 ^ n3351 ^ x95 ;
  assign n3539 = n3506 ^ n3351 ^ 1'b0 ;
  assign n3540 = ( n3351 & n3538 ) | ( n3351 & ~n3539 ) | ( n3538 & ~n3539 ) ;
  assign n3541 = n3495 ^ n3373 ^ x94 ;
  assign n3542 = n3506 ^ n3373 ^ 1'b0 ;
  assign n3543 = ( n3373 & n3541 ) | ( n3373 & ~n3542 ) | ( n3541 & ~n3542 ) ;
  assign n3544 = n3494 ^ n3380 ^ x93 ;
  assign n3545 = n3506 ^ n3380 ^ 1'b0 ;
  assign n3546 = ( n3380 & n3544 ) | ( n3380 & ~n3545 ) | ( n3544 & ~n3545 ) ;
  assign n3547 = n3492 ^ n3355 ^ x91 ;
  assign n3548 = n3506 ^ n3355 ^ 1'b0 ;
  assign n3549 = ( n3355 & n3547 ) | ( n3355 & ~n3548 ) | ( n3547 & ~n3548 ) ;
  assign n3550 = n3491 ^ n3384 ^ x90 ;
  assign n3551 = n3506 ^ n3384 ^ 1'b0 ;
  assign n3552 = ( n3384 & n3550 ) | ( n3384 & ~n3551 ) | ( n3550 & ~n3551 ) ;
  assign n3553 = n3506 ^ n3387 ^ 1'b0 ;
  assign n3554 = n3489 ^ n3469 ^ x88 ;
  assign n3555 = n3506 ^ n3469 ^ 1'b0 ;
  assign n3556 = ( n3469 & n3554 ) | ( n3469 & ~n3555 ) | ( n3554 & ~n3555 ) ;
  assign n3557 = n3488 ^ n3465 ^ x87 ;
  assign n3558 = n3487 ^ n3442 ^ x86 ;
  assign n3559 = n3506 ^ n3442 ^ 1'b0 ;
  assign n3560 = ( n3442 & n3558 ) | ( n3442 & ~n3559 ) | ( n3558 & ~n3559 ) ;
  assign n3561 = n3506 ^ n3461 ^ 1'b0 ;
  assign n3562 = n3486 ^ n3461 ^ x85 ;
  assign n3563 = ( n3461 & ~n3561 ) | ( n3461 & n3562 ) | ( ~n3561 & n3562 ) ;
  assign n3564 = n3485 ^ n3445 ^ x84 ;
  assign n3565 = n3506 ^ n3445 ^ 1'b0 ;
  assign n3566 = ( n3445 & n3564 ) | ( n3445 & ~n3565 ) | ( n3564 & ~n3565 ) ;
  assign n3567 = n3483 ^ n3393 ^ x82 ;
  assign n3568 = n3506 ^ n3393 ^ 1'b0 ;
  assign n3569 = ( n3393 & n3567 ) | ( n3393 & ~n3568 ) | ( n3567 & ~n3568 ) ;
  assign n3570 = n3480 ^ n3407 ^ x79 ;
  assign n3571 = n3506 ^ n3407 ^ 1'b0 ;
  assign n3572 = ( n3407 & n3570 ) | ( n3407 & ~n3571 ) | ( n3570 & ~n3571 ) ;
  assign n3573 = n3477 ^ n3411 ^ x76 ;
  assign n3574 = ( n3387 & n3510 ) | ( n3387 & ~n3553 ) | ( n3510 & ~n3553 ) ;
  assign n3575 = n3506 ^ n3411 ^ 1'b0 ;
  assign n3576 = ( n3411 & n3573 ) | ( n3411 & ~n3575 ) | ( n3573 & ~n3575 ) ;
  assign n3577 = n3475 ^ n3417 ^ x74 ;
  assign n3578 = n3506 ^ n3417 ^ 1'b0 ;
  assign n3579 = ( n3417 & n3577 ) | ( n3417 & ~n3578 ) | ( n3577 & ~n3578 ) ;
  assign n3580 = n3472 ^ n3423 ^ x72 ;
  assign n3581 = n3506 ^ n3423 ^ 1'b0 ;
  assign n3582 = ( n3423 & n3580 ) | ( n3423 & ~n3581 ) | ( n3580 & ~n3581 ) ;
  assign n3583 = n3506 ^ n3451 ^ 1'b0 ;
  assign n3584 = ( n3375 & n3451 ) | ( n3375 & n3583 ) | ( n3451 & n3583 ) ;
  assign n3585 = n3506 ^ n3377 ^ 1'b0 ;
  assign n3586 = x64 & n3506 ;
  assign n3587 = n3586 ^ x64 ^ x25 ;
  assign n3588 = n3506 ^ n3446 ^ 1'b0 ;
  assign n3589 = ( n3440 & n3446 ) | ( n3440 & n3588 ) | ( n3446 & n3588 ) ;
  assign n3590 = n3506 ^ n3372 ^ 1'b0 ;
  assign n3591 = n3506 ^ n3465 ^ 1'b0 ;
  assign n3592 = n3506 ^ n3399 ^ 1'b0 ;
  assign n3593 = ~x24 & x64 ;
  assign n3594 = n3506 ^ n3371 ^ 1'b0 ;
  assign n3595 = ~n3273 & n3593 ;
  assign n3596 = ( n3465 & n3557 ) | ( n3465 & ~n3591 ) | ( n3557 & ~n3591 ) ;
  assign n3597 = n3593 ^ n3587 ^ x65 ;
  assign n3598 = ( x65 & n3593 ) | ( x65 & n3597 ) | ( n3593 & n3597 ) ;
  assign n3599 = n3501 ^ n3372 ^ x100 ;
  assign n3600 = n3598 ^ n3589 ^ x66 ;
  assign n3601 = ( x66 & n3598 ) | ( x66 & n3600 ) | ( n3598 & n3600 ) ;
  assign n3602 = n3481 ^ n3399 ^ x80 ;
  assign n3603 = ( n3399 & ~n3592 ) | ( n3399 & n3602 ) | ( ~n3592 & n3602 ) ;
  assign n3604 = n3482 ^ n3396 ^ x81 ;
  assign n3605 = n3506 ^ n3396 ^ 1'b0 ;
  assign n3606 = ( n3396 & n3604 ) | ( n3396 & ~n3605 ) | ( n3604 & ~n3605 ) ;
  assign n3607 = n3500 ^ n3377 ^ x99 ;
  assign n3608 = n3474 ^ n3420 ^ x73 ;
  assign n3609 = n3498 ^ n3379 ^ x97 ;
  assign n3610 = n3506 ^ n3379 ^ 1'b0 ;
  assign n3611 = n3506 ^ n3381 ^ 1'b0 ;
  assign n3612 = ( x67 & ~n3584 ) | ( x67 & n3601 ) | ( ~n3584 & n3601 ) ;
  assign n3613 = n3499 ^ n3371 ^ x98 ;
  assign n3614 = ( n3371 & ~n3594 ) | ( n3371 & n3613 ) | ( ~n3594 & n3613 ) ;
  assign n3615 = ( n3372 & ~n3590 ) | ( n3372 & n3599 ) | ( ~n3590 & n3599 ) ;
  assign n3616 = n3502 ^ n3381 ^ x101 ;
  assign n3617 = n3506 ^ n3420 ^ 1'b0 ;
  assign n3618 = ( n3379 & n3609 ) | ( n3379 & ~n3610 ) | ( n3609 & ~n3610 ) ;
  assign n3619 = ( x68 & ~n3532 ) | ( x68 & n3612 ) | ( ~n3532 & n3612 ) ;
  assign n3620 = ( n3377 & ~n3585 ) | ( n3377 & n3607 ) | ( ~n3585 & n3607 ) ;
  assign n3621 = ( x69 & ~n3530 ) | ( x69 & n3619 ) | ( ~n3530 & n3619 ) ;
  assign n3622 = ( x70 & ~n3528 ) | ( x70 & n3621 ) | ( ~n3528 & n3621 ) ;
  assign n3623 = ( x71 & ~n3526 ) | ( x71 & n3622 ) | ( ~n3526 & n3622 ) ;
  assign n3624 = ( x72 & ~n3524 ) | ( x72 & n3623 ) | ( ~n3524 & n3623 ) ;
  assign n3625 = ( x73 & ~n3582 ) | ( x73 & n3624 ) | ( ~n3582 & n3624 ) ;
  assign n3626 = ( n3420 & n3608 ) | ( n3420 & ~n3617 ) | ( n3608 & ~n3617 ) ;
  assign n3627 = ( x74 & n3625 ) | ( x74 & ~n3626 ) | ( n3625 & ~n3626 ) ;
  assign n3628 = ( x75 & ~n3579 ) | ( x75 & n3627 ) | ( ~n3579 & n3627 ) ;
  assign n3629 = ( x76 & ~n3522 ) | ( x76 & n3628 ) | ( ~n3522 & n3628 ) ;
  assign n3630 = ( n3381 & ~n3611 ) | ( n3381 & n3616 ) | ( ~n3611 & n3616 ) ;
  assign n3631 = ( x77 & ~n3576 ) | ( x77 & n3629 ) | ( ~n3576 & n3629 ) ;
  assign n3632 = ( x78 & ~n3519 ) | ( x78 & n3631 ) | ( ~n3519 & n3631 ) ;
  assign n3633 = ( x79 & ~n3516 ) | ( x79 & n3632 ) | ( ~n3516 & n3632 ) ;
  assign n3634 = ( x80 & ~n3572 ) | ( x80 & n3633 ) | ( ~n3572 & n3633 ) ;
  assign n3635 = ( x81 & ~n3603 ) | ( x81 & n3634 ) | ( ~n3603 & n3634 ) ;
  assign n3636 = ( x82 & ~n3606 ) | ( x82 & n3635 ) | ( ~n3606 & n3635 ) ;
  assign n3637 = ( x83 & ~n3569 ) | ( x83 & n3636 ) | ( ~n3569 & n3636 ) ;
  assign n3638 = ( x84 & ~n3513 ) | ( x84 & n3637 ) | ( ~n3513 & n3637 ) ;
  assign n3639 = ( x85 & ~n3566 ) | ( x85 & n3638 ) | ( ~n3566 & n3638 ) ;
  assign n3640 = ( x86 & ~n3563 ) | ( x86 & n3639 ) | ( ~n3563 & n3639 ) ;
  assign n3641 = ( x87 & ~n3560 ) | ( x87 & n3640 ) | ( ~n3560 & n3640 ) ;
  assign n3642 = ( x88 & ~n3596 ) | ( x88 & n3641 ) | ( ~n3596 & n3641 ) ;
  assign n3643 = ( x89 & ~n3556 ) | ( x89 & n3642 ) | ( ~n3556 & n3642 ) ;
  assign n3644 = ( x90 & ~n3574 ) | ( x90 & n3643 ) | ( ~n3574 & n3643 ) ;
  assign n3645 = ( x91 & ~n3552 ) | ( x91 & n3644 ) | ( ~n3552 & n3644 ) ;
  assign n3646 = ( x92 & ~n3549 ) | ( x92 & n3645 ) | ( ~n3549 & n3645 ) ;
  assign n3647 = ( x93 & ~n3509 ) | ( x93 & n3646 ) | ( ~n3509 & n3646 ) ;
  assign n3648 = ( x94 & ~n3546 ) | ( x94 & n3647 ) | ( ~n3546 & n3647 ) ;
  assign n3649 = ( x95 & ~n3543 ) | ( x95 & n3648 ) | ( ~n3543 & n3648 ) ;
  assign n3650 = n3649 ^ n3540 ^ x96 ;
  assign n3651 = n3646 ^ n3509 ^ x93 ;
  assign n3652 = n3647 ^ n3546 ^ x94 ;
  assign n3653 = ( x96 & ~n3540 ) | ( x96 & n3649 ) | ( ~n3540 & n3649 ) ;
  assign n3654 = ( x97 & ~n3537 ) | ( x97 & n3653 ) | ( ~n3537 & n3653 ) ;
  assign n3655 = ( x98 & ~n3618 ) | ( x98 & n3654 ) | ( ~n3618 & n3654 ) ;
  assign n3656 = ( x99 & ~n3614 ) | ( x99 & n3655 ) | ( ~n3614 & n3655 ) ;
  assign n3657 = ( x100 & ~n3620 ) | ( x100 & n3656 ) | ( ~n3620 & n3656 ) ;
  assign n3658 = ( x101 & ~n3615 ) | ( x101 & n3657 ) | ( ~n3615 & n3657 ) ;
  assign n3659 = ( x102 & ~n3630 ) | ( x102 & n3658 ) | ( ~n3630 & n3658 ) ;
  assign n3660 = ( x103 & ~n3534 ) | ( x103 & n3659 ) | ( ~n3534 & n3659 ) ;
  assign n3661 = ( ~n189 & n3595 ) | ( ~n189 & n3660 ) | ( n3595 & n3660 ) ;
  assign n3662 = n2744 | n3660 ;
  assign n3663 = n3656 ^ n3620 ^ x100 ;
  assign n3664 = n3662 ^ n3546 ^ 1'b0 ;
  assign n3665 = n3658 ^ n3630 ^ x102 ;
  assign n3666 = n3653 ^ n3537 ^ x97 ;
  assign n3667 = ( n3546 & n3652 ) | ( n3546 & ~n3664 ) | ( n3652 & ~n3664 ) ;
  assign n3668 = n3662 ^ n3597 ^ 1'b0 ;
  assign n3669 = n3662 ^ n3509 ^ 1'b0 ;
  assign n3670 = ( n3509 & n3651 ) | ( n3509 & ~n3669 ) | ( n3651 & ~n3669 ) ;
  assign n3671 = n3655 ^ n3614 ^ x99 ;
  assign n3672 = n3662 ^ n3614 ^ 1'b0 ;
  assign n3673 = n3648 ^ n3543 ^ x95 ;
  assign n3674 = n3662 ^ n3543 ^ 1'b0 ;
  assign n3675 = ( n3543 & n3673 ) | ( n3543 & ~n3674 ) | ( n3673 & ~n3674 ) ;
  assign n3676 = ( n3614 & n3671 ) | ( n3614 & ~n3672 ) | ( n3671 & ~n3672 ) ;
  assign n3677 = n3662 ^ n3600 ^ 1'b0 ;
  assign n3678 = n3662 ^ n3537 ^ 1'b0 ;
  assign n3679 = ( n3589 & n3600 ) | ( n3589 & n3677 ) | ( n3600 & n3677 ) ;
  assign n3680 = n3662 ^ n3615 ^ 1'b0 ;
  assign n3681 = ( n3587 & n3597 ) | ( n3587 & n3668 ) | ( n3597 & n3668 ) ;
  assign n3682 = n3657 ^ n3615 ^ x101 ;
  assign n3683 = n3662 ^ n3540 ^ 1'b0 ;
  assign n3684 = n3662 ^ n3620 ^ 1'b0 ;
  assign n3685 = ( n3537 & n3666 ) | ( n3537 & ~n3678 ) | ( n3666 & ~n3678 ) ;
  assign n3686 = n3665 ^ n3662 ^ 1'b0 ;
  assign n3687 = ( n3630 & n3665 ) | ( n3630 & n3686 ) | ( n3665 & n3686 ) ;
  assign n3688 = ( n3540 & n3650 ) | ( n3540 & ~n3683 ) | ( n3650 & ~n3683 ) ;
  assign n3689 = ( n3620 & n3663 ) | ( n3620 & ~n3684 ) | ( n3663 & ~n3684 ) ;
  assign n3690 = ( n3615 & ~n3680 ) | ( n3615 & n3682 ) | ( ~n3680 & n3682 ) ;
  assign n3691 = n3644 ^ n3552 ^ x91 ;
  assign n3692 = n3662 ^ n3552 ^ 1'b0 ;
  assign n3693 = ( n3552 & n3691 ) | ( n3552 & ~n3692 ) | ( n3691 & ~n3692 ) ;
  assign n3694 = n3640 ^ n3560 ^ x87 ;
  assign n3695 = n3662 ^ n3560 ^ 1'b0 ;
  assign n3696 = ( n3560 & n3694 ) | ( n3560 & ~n3695 ) | ( n3694 & ~n3695 ) ;
  assign n3697 = n3638 ^ n3566 ^ x85 ;
  assign n3698 = n3662 ^ n3566 ^ 1'b0 ;
  assign n3699 = ( n3566 & n3697 ) | ( n3566 & ~n3698 ) | ( n3697 & ~n3698 ) ;
  assign n3700 = n3637 ^ n3513 ^ x84 ;
  assign n3701 = n3662 ^ n3513 ^ 1'b0 ;
  assign n3702 = ( n3513 & n3700 ) | ( n3513 & ~n3701 ) | ( n3700 & ~n3701 ) ;
  assign n3703 = n3636 ^ n3569 ^ x83 ;
  assign n3704 = n3662 ^ n3569 ^ 1'b0 ;
  assign n3705 = ( n3569 & n3703 ) | ( n3569 & ~n3704 ) | ( n3703 & ~n3704 ) ;
  assign n3706 = n3635 ^ n3606 ^ x82 ;
  assign n3707 = n3662 ^ n3606 ^ 1'b0 ;
  assign n3708 = ( n3606 & n3706 ) | ( n3606 & ~n3707 ) | ( n3706 & ~n3707 ) ;
  assign n3709 = n3662 ^ n3603 ^ 1'b0 ;
  assign n3710 = n3632 ^ n3516 ^ x79 ;
  assign n3711 = n3662 ^ n3516 ^ 1'b0 ;
  assign n3712 = ( n3516 & n3710 ) | ( n3516 & ~n3711 ) | ( n3710 & ~n3711 ) ;
  assign n3713 = n3631 ^ n3519 ^ x78 ;
  assign n3714 = n3662 ^ n3519 ^ 1'b0 ;
  assign n3715 = n3634 ^ n3603 ^ x81 ;
  assign n3716 = ( n3603 & ~n3709 ) | ( n3603 & n3715 ) | ( ~n3709 & n3715 ) ;
  assign n3717 = ( n3519 & n3713 ) | ( n3519 & ~n3714 ) | ( n3713 & ~n3714 ) ;
  assign n3718 = n3627 ^ n3579 ^ x75 ;
  assign n3719 = n3662 ^ n3579 ^ 1'b0 ;
  assign n3720 = ( n3579 & n3718 ) | ( n3579 & ~n3719 ) | ( n3718 & ~n3719 ) ;
  assign n3721 = n3624 ^ n3582 ^ x73 ;
  assign n3722 = n3662 ^ n3582 ^ 1'b0 ;
  assign n3723 = ( n3582 & n3721 ) | ( n3582 & ~n3722 ) | ( n3721 & ~n3722 ) ;
  assign n3724 = n3623 ^ n3524 ^ x72 ;
  assign n3725 = n3662 ^ n3524 ^ 1'b0 ;
  assign n3726 = ( n3524 & n3724 ) | ( n3524 & ~n3725 ) | ( n3724 & ~n3725 ) ;
  assign n3727 = n3622 ^ n3526 ^ x71 ;
  assign n3728 = n3662 ^ n3526 ^ 1'b0 ;
  assign n3729 = ( n3526 & n3727 ) | ( n3526 & ~n3728 ) | ( n3727 & ~n3728 ) ;
  assign n3730 = n3619 ^ n3530 ^ x69 ;
  assign n3731 = n3662 ^ n3530 ^ 1'b0 ;
  assign n3732 = ( n3530 & n3730 ) | ( n3530 & ~n3731 ) | ( n3730 & ~n3731 ) ;
  assign n3733 = n3612 ^ n3532 ^ x68 ;
  assign n3734 = n3662 ^ n3532 ^ 1'b0 ;
  assign n3735 = ( n3532 & n3733 ) | ( n3532 & ~n3734 ) | ( n3733 & ~n3734 ) ;
  assign n3736 = n3601 ^ n3584 ^ x67 ;
  assign n3737 = n3662 ^ n3584 ^ 1'b0 ;
  assign n3738 = ( n3584 & n3736 ) | ( n3584 & ~n3737 ) | ( n3736 & ~n3737 ) ;
  assign n3739 = n3654 ^ n3618 ^ x98 ;
  assign n3740 = n3662 ^ n3618 ^ 1'b0 ;
  assign n3741 = ( n3618 & n3739 ) | ( n3618 & ~n3740 ) | ( n3739 & ~n3740 ) ;
  assign n3742 = n3645 ^ n3549 ^ x92 ;
  assign n3743 = n3662 ^ n3549 ^ 1'b0 ;
  assign n3744 = ( n3549 & n3742 ) | ( n3549 & ~n3743 ) | ( n3742 & ~n3743 ) ;
  assign n3745 = n3643 ^ n3574 ^ x90 ;
  assign n3746 = n3662 ^ n3574 ^ 1'b0 ;
  assign n3747 = ( n3574 & n3745 ) | ( n3574 & ~n3746 ) | ( n3745 & ~n3746 ) ;
  assign n3748 = n3642 ^ n3556 ^ x89 ;
  assign n3749 = n3662 ^ n3556 ^ 1'b0 ;
  assign n3750 = ( n3556 & n3748 ) | ( n3556 & ~n3749 ) | ( n3748 & ~n3749 ) ;
  assign n3751 = n3641 ^ n3596 ^ x88 ;
  assign n3752 = n3662 ^ n3596 ^ 1'b0 ;
  assign n3753 = ( n3596 & n3751 ) | ( n3596 & ~n3752 ) | ( n3751 & ~n3752 ) ;
  assign n3754 = n3662 ^ n3563 ^ 1'b0 ;
  assign n3755 = n3633 ^ n3572 ^ x80 ;
  assign n3756 = n3662 ^ n3572 ^ 1'b0 ;
  assign n3757 = ( n3572 & n3755 ) | ( n3572 & ~n3756 ) | ( n3755 & ~n3756 ) ;
  assign n3758 = n3629 ^ n3576 ^ x77 ;
  assign n3759 = n3662 ^ n3576 ^ 1'b0 ;
  assign n3760 = ( n3576 & n3758 ) | ( n3576 & ~n3759 ) | ( n3758 & ~n3759 ) ;
  assign n3761 = n3628 ^ n3522 ^ x76 ;
  assign n3762 = n3662 ^ n3522 ^ 1'b0 ;
  assign n3763 = ( n3522 & n3761 ) | ( n3522 & ~n3762 ) | ( n3761 & ~n3762 ) ;
  assign n3764 = n3626 ^ n3625 ^ x74 ;
  assign n3765 = n3662 ^ n3626 ^ 1'b0 ;
  assign n3766 = ( n3626 & n3764 ) | ( n3626 & ~n3765 ) | ( n3764 & ~n3765 ) ;
  assign n3767 = n3621 ^ n3528 ^ x70 ;
  assign n3768 = n3639 ^ n3563 ^ x86 ;
  assign n3769 = ( n3563 & ~n3754 ) | ( n3563 & n3768 ) | ( ~n3754 & n3768 ) ;
  assign n3770 = n3662 ^ n3528 ^ 1'b0 ;
  assign n3771 = ( n3528 & n3767 ) | ( n3528 & ~n3770 ) | ( n3767 & ~n3770 ) ;
  assign n3772 = ~n3660 & n3661 ;
  assign n3773 = x104 | n151 ;
  assign n3774 = ( ~x24 & x64 ) | ( ~x24 & n3773 ) | ( x64 & n3773 ) ;
  assign n3775 = x64 & ~n3774 ;
  assign n3776 = ( ~n176 & n3660 ) | ( ~n176 & n3775 ) | ( n3660 & n3775 ) ;
  assign n3777 = ~n3660 & n3776 ;
  assign n3778 = ( x24 & n3772 ) | ( x24 & ~n3777 ) | ( n3772 & ~n3777 ) ;
  assign n3779 = ( n322 & n3534 ) | ( n322 & n3662 ) | ( n3534 & n3662 ) ;
  assign n3780 = ( ~x106 & x107 ) | ( ~x106 & n193 ) | ( x107 & n193 ) ;
  assign n3781 = ~x23 & x64 ;
  assign n3782 = n3781 ^ n3778 ^ x65 ;
  assign n3783 = ( x65 & n3781 ) | ( x65 & n3782 ) | ( n3781 & n3782 ) ;
  assign n3784 = n3783 ^ n3681 ^ x66 ;
  assign n3785 = ( x66 & n3783 ) | ( x66 & n3784 ) | ( n3783 & n3784 ) ;
  assign n3786 = ( x67 & ~n3679 ) | ( x67 & n3785 ) | ( ~n3679 & n3785 ) ;
  assign n3787 = ( x68 & ~n3738 ) | ( x68 & n3786 ) | ( ~n3738 & n3786 ) ;
  assign n3788 = ( x69 & ~n3735 ) | ( x69 & n3787 ) | ( ~n3735 & n3787 ) ;
  assign n3789 = ( x70 & ~n3732 ) | ( x70 & n3788 ) | ( ~n3732 & n3788 ) ;
  assign n3790 = ( x71 & ~n3771 ) | ( x71 & n3789 ) | ( ~n3771 & n3789 ) ;
  assign n3791 = ( x72 & ~n3729 ) | ( x72 & n3790 ) | ( ~n3729 & n3790 ) ;
  assign n3792 = ( x73 & ~n3726 ) | ( x73 & n3791 ) | ( ~n3726 & n3791 ) ;
  assign n3793 = ( x74 & ~n3723 ) | ( x74 & n3792 ) | ( ~n3723 & n3792 ) ;
  assign n3794 = ( x75 & ~n3766 ) | ( x75 & n3793 ) | ( ~n3766 & n3793 ) ;
  assign n3795 = ( x76 & ~n3720 ) | ( x76 & n3794 ) | ( ~n3720 & n3794 ) ;
  assign n3796 = ( x77 & ~n3763 ) | ( x77 & n3795 ) | ( ~n3763 & n3795 ) ;
  assign n3797 = ( x78 & ~n3760 ) | ( x78 & n3796 ) | ( ~n3760 & n3796 ) ;
  assign n3798 = ( x79 & ~n3717 ) | ( x79 & n3797 ) | ( ~n3717 & n3797 ) ;
  assign n3799 = ( x80 & ~n3712 ) | ( x80 & n3798 ) | ( ~n3712 & n3798 ) ;
  assign n3800 = ( x81 & ~n3757 ) | ( x81 & n3799 ) | ( ~n3757 & n3799 ) ;
  assign n3801 = ( x82 & ~n3716 ) | ( x82 & n3800 ) | ( ~n3716 & n3800 ) ;
  assign n3802 = ( x83 & ~n3708 ) | ( x83 & n3801 ) | ( ~n3708 & n3801 ) ;
  assign n3803 = ( x84 & ~n3705 ) | ( x84 & n3802 ) | ( ~n3705 & n3802 ) ;
  assign n3804 = n3791 ^ n3726 ^ x73 ;
  assign n3805 = ( x85 & ~n3702 ) | ( x85 & n3803 ) | ( ~n3702 & n3803 ) ;
  assign n3806 = ( x86 & ~n3699 ) | ( x86 & n3805 ) | ( ~n3699 & n3805 ) ;
  assign n3807 = n3794 ^ n3720 ^ x76 ;
  assign n3808 = ( x87 & ~n3769 ) | ( x87 & n3806 ) | ( ~n3769 & n3806 ) ;
  assign n3809 = ( x88 & ~n3696 ) | ( x88 & n3808 ) | ( ~n3696 & n3808 ) ;
  assign n3810 = n3797 ^ n3717 ^ x79 ;
  assign n3811 = n3790 ^ n3729 ^ x72 ;
  assign n3812 = n3789 ^ n3771 ^ x71 ;
  assign n3813 = n3800 ^ n3716 ^ x82 ;
  assign n3814 = n3787 ^ n3735 ^ x69 ;
  assign n3815 = n3802 ^ n3705 ^ x84 ;
  assign n3816 = n3803 ^ n3702 ^ x85 ;
  assign n3817 = n3808 ^ n3696 ^ x88 ;
  assign n3818 = ~n151 & n3781 ;
  assign n3819 = ( x89 & ~n3753 ) | ( x89 & n3809 ) | ( ~n3753 & n3809 ) ;
  assign n3820 = n3785 ^ n3679 ^ x67 ;
  assign n3821 = n3809 ^ n3753 ^ x89 ;
  assign n3822 = ( x90 & ~n3750 ) | ( x90 & n3819 ) | ( ~n3750 & n3819 ) ;
  assign n3823 = ( x91 & ~n3747 ) | ( x91 & n3822 ) | ( ~n3747 & n3822 ) ;
  assign n3824 = ( x92 & ~n3693 ) | ( x92 & n3823 ) | ( ~n3693 & n3823 ) ;
  assign n3825 = ( x93 & ~n3744 ) | ( x93 & n3824 ) | ( ~n3744 & n3824 ) ;
  assign n3826 = ( x94 & ~n3670 ) | ( x94 & n3825 ) | ( ~n3670 & n3825 ) ;
  assign n3827 = ( x95 & ~n3667 ) | ( x95 & n3826 ) | ( ~n3667 & n3826 ) ;
  assign n3828 = ( x96 & ~n3675 ) | ( x96 & n3827 ) | ( ~n3675 & n3827 ) ;
  assign n3829 = ( x97 & ~n3688 ) | ( x97 & n3828 ) | ( ~n3688 & n3828 ) ;
  assign n3830 = ( x98 & ~n3685 ) | ( x98 & n3829 ) | ( ~n3685 & n3829 ) ;
  assign n3831 = ( x99 & ~n3741 ) | ( x99 & n3830 ) | ( ~n3741 & n3830 ) ;
  assign n3832 = ( x100 & ~n3676 ) | ( x100 & n3831 ) | ( ~n3676 & n3831 ) ;
  assign n3833 = ( x101 & ~n3689 ) | ( x101 & n3832 ) | ( ~n3689 & n3832 ) ;
  assign n3834 = ( x102 & ~n3690 ) | ( x102 & n3833 ) | ( ~n3690 & n3833 ) ;
  assign n3835 = ( x103 & ~n3687 ) | ( x103 & n3834 ) | ( ~n3687 & n3834 ) ;
  assign n3836 = ( x104 & ~n3779 ) | ( x104 & n3835 ) | ( ~n3779 & n3835 ) ;
  assign n3837 = n162 | n3836 ;
  assign n3838 = n3827 ^ n3675 ^ x96 ;
  assign n3839 = n3837 ^ n3675 ^ 1'b0 ;
  assign n3840 = ( n3675 & n3838 ) | ( n3675 & ~n3839 ) | ( n3838 & ~n3839 ) ;
  assign n3841 = n3826 ^ n3667 ^ x95 ;
  assign n3842 = n3837 ^ n3667 ^ 1'b0 ;
  assign n3843 = ( n3667 & n3841 ) | ( n3667 & ~n3842 ) | ( n3841 & ~n3842 ) ;
  assign n3844 = n3837 ^ n3753 ^ 1'b0 ;
  assign n3845 = ( n3753 & n3821 ) | ( n3753 & ~n3844 ) | ( n3821 & ~n3844 ) ;
  assign n3846 = n3837 ^ n3696 ^ 1'b0 ;
  assign n3847 = ( n3696 & n3817 ) | ( n3696 & ~n3846 ) | ( n3817 & ~n3846 ) ;
  assign n3848 = n3837 ^ n3702 ^ 1'b0 ;
  assign n3849 = ( n3702 & n3816 ) | ( n3702 & ~n3848 ) | ( n3816 & ~n3848 ) ;
  assign n3850 = n3837 ^ n3705 ^ 1'b0 ;
  assign n3851 = ( n3705 & n3815 ) | ( n3705 & ~n3850 ) | ( n3815 & ~n3850 ) ;
  assign n3852 = n3837 ^ n3716 ^ 1'b0 ;
  assign n3853 = ( n3716 & n3813 ) | ( n3716 & ~n3852 ) | ( n3813 & ~n3852 ) ;
  assign n3854 = n3837 ^ n3717 ^ 1'b0 ;
  assign n3855 = ( n3717 & n3810 ) | ( n3717 & ~n3854 ) | ( n3810 & ~n3854 ) ;
  assign n3856 = n3837 ^ n3720 ^ 1'b0 ;
  assign n3857 = ( n3720 & n3807 ) | ( n3720 & ~n3856 ) | ( n3807 & ~n3856 ) ;
  assign n3858 = n3837 ^ n3726 ^ 1'b0 ;
  assign n3859 = ( n3726 & n3804 ) | ( n3726 & ~n3858 ) | ( n3804 & ~n3858 ) ;
  assign n3860 = n3837 ^ n3729 ^ 1'b0 ;
  assign n3861 = ( n3729 & n3811 ) | ( n3729 & ~n3860 ) | ( n3811 & ~n3860 ) ;
  assign n3862 = n3837 ^ n3771 ^ 1'b0 ;
  assign n3863 = ( n3771 & n3812 ) | ( n3771 & ~n3862 ) | ( n3812 & ~n3862 ) ;
  assign n3864 = n3837 ^ n3735 ^ 1'b0 ;
  assign n3865 = ( n3735 & n3814 ) | ( n3735 & ~n3864 ) | ( n3814 & ~n3864 ) ;
  assign n3866 = n3837 ^ n3679 ^ 1'b0 ;
  assign n3867 = ( n3679 & n3820 ) | ( n3679 & ~n3866 ) | ( n3820 & ~n3866 ) ;
  assign n3868 = n3837 ^ n3784 ^ 1'b0 ;
  assign n3869 = ( n3681 & n3784 ) | ( n3681 & n3868 ) | ( n3784 & n3868 ) ;
  assign n3870 = n3837 ^ n3782 ^ 1'b0 ;
  assign n3871 = ( n3778 & n3782 ) | ( n3778 & n3870 ) | ( n3782 & n3870 ) ;
  assign n3872 = n3834 ^ n3687 ^ x103 ;
  assign n3873 = n3872 ^ n3837 ^ 1'b0 ;
  assign n3874 = ( n3687 & n3872 ) | ( n3687 & n3873 ) | ( n3872 & n3873 ) ;
  assign n3875 = n3837 ^ n3690 ^ 1'b0 ;
  assign n3876 = n3832 ^ n3689 ^ x101 ;
  assign n3877 = n3837 ^ n3689 ^ 1'b0 ;
  assign n3878 = ( n3689 & n3876 ) | ( n3689 & ~n3877 ) | ( n3876 & ~n3877 ) ;
  assign n3879 = n3831 ^ n3676 ^ x100 ;
  assign n3880 = n3837 ^ n3676 ^ 1'b0 ;
  assign n3881 = ( n3676 & n3879 ) | ( n3676 & ~n3880 ) | ( n3879 & ~n3880 ) ;
  assign n3882 = n3830 ^ n3741 ^ x99 ;
  assign n3883 = n3837 ^ n3741 ^ 1'b0 ;
  assign n3884 = ( n3741 & n3882 ) | ( n3741 & ~n3883 ) | ( n3882 & ~n3883 ) ;
  assign n3885 = n3829 ^ n3685 ^ x98 ;
  assign n3886 = n3837 ^ n3685 ^ 1'b0 ;
  assign n3887 = ( n3685 & n3885 ) | ( n3685 & ~n3886 ) | ( n3885 & ~n3886 ) ;
  assign n3888 = n3828 ^ n3688 ^ x97 ;
  assign n3889 = n3837 ^ n3688 ^ 1'b0 ;
  assign n3890 = ( n3688 & n3888 ) | ( n3688 & ~n3889 ) | ( n3888 & ~n3889 ) ;
  assign n3891 = n3833 ^ n3690 ^ x102 ;
  assign n3892 = ( n3690 & ~n3875 ) | ( n3690 & n3891 ) | ( ~n3875 & n3891 ) ;
  assign n3893 = n3825 ^ n3670 ^ x94 ;
  assign n3894 = n3837 ^ n3670 ^ 1'b0 ;
  assign n3895 = ( n3670 & n3893 ) | ( n3670 & ~n3894 ) | ( n3893 & ~n3894 ) ;
  assign n3896 = n3824 ^ n3744 ^ x93 ;
  assign n3897 = n3837 ^ n3744 ^ 1'b0 ;
  assign n3898 = ( n3744 & n3896 ) | ( n3744 & ~n3897 ) | ( n3896 & ~n3897 ) ;
  assign n3899 = n3823 ^ n3693 ^ x92 ;
  assign n3900 = n3837 ^ n3693 ^ 1'b0 ;
  assign n3901 = ( n3693 & n3899 ) | ( n3693 & ~n3900 ) | ( n3899 & ~n3900 ) ;
  assign n3902 = n3822 ^ n3747 ^ x91 ;
  assign n3903 = n3837 ^ n3747 ^ 1'b0 ;
  assign n3904 = ( n3747 & n3902 ) | ( n3747 & ~n3903 ) | ( n3902 & ~n3903 ) ;
  assign n3905 = n3819 ^ n3750 ^ x90 ;
  assign n3906 = n3837 ^ n3750 ^ 1'b0 ;
  assign n3907 = ( n3750 & n3905 ) | ( n3750 & ~n3906 ) | ( n3905 & ~n3906 ) ;
  assign n3908 = n3806 ^ n3769 ^ x87 ;
  assign n3909 = n3837 ^ n3769 ^ 1'b0 ;
  assign n3910 = ( n3769 & n3908 ) | ( n3769 & ~n3909 ) | ( n3908 & ~n3909 ) ;
  assign n3911 = n3805 ^ n3699 ^ x86 ;
  assign n3912 = n3837 ^ n3699 ^ 1'b0 ;
  assign n3913 = ( n3699 & n3911 ) | ( n3699 & ~n3912 ) | ( n3911 & ~n3912 ) ;
  assign n3914 = n3801 ^ n3708 ^ x83 ;
  assign n3915 = n3837 ^ n3708 ^ 1'b0 ;
  assign n3916 = ( n3708 & n3914 ) | ( n3708 & ~n3915 ) | ( n3914 & ~n3915 ) ;
  assign n3917 = n3799 ^ n3757 ^ x81 ;
  assign n3918 = n3837 ^ n3757 ^ 1'b0 ;
  assign n3919 = ( n3757 & n3917 ) | ( n3757 & ~n3918 ) | ( n3917 & ~n3918 ) ;
  assign n3920 = n3798 ^ n3712 ^ x80 ;
  assign n3921 = n3837 ^ n3712 ^ 1'b0 ;
  assign n3922 = ( n3712 & n3920 ) | ( n3712 & ~n3921 ) | ( n3920 & ~n3921 ) ;
  assign n3923 = n3796 ^ n3760 ^ x78 ;
  assign n3924 = n3837 ^ n3760 ^ 1'b0 ;
  assign n3925 = ( n3760 & n3923 ) | ( n3760 & ~n3924 ) | ( n3923 & ~n3924 ) ;
  assign n3926 = n3795 ^ n3763 ^ x77 ;
  assign n3927 = n3837 ^ n3763 ^ 1'b0 ;
  assign n3928 = ( n3763 & n3926 ) | ( n3763 & ~n3927 ) | ( n3926 & ~n3927 ) ;
  assign n3929 = n3793 ^ n3766 ^ x75 ;
  assign n3930 = n3837 ^ n3766 ^ 1'b0 ;
  assign n3931 = ( n3766 & n3929 ) | ( n3766 & ~n3930 ) | ( n3929 & ~n3930 ) ;
  assign n3932 = n3792 ^ n3723 ^ x74 ;
  assign n3933 = n3837 ^ n3723 ^ 1'b0 ;
  assign n3934 = ( n3723 & n3932 ) | ( n3723 & ~n3933 ) | ( n3932 & ~n3933 ) ;
  assign n3935 = n3788 ^ n3732 ^ x70 ;
  assign n3936 = n3837 ^ n3732 ^ 1'b0 ;
  assign n3937 = ( n3732 & n3935 ) | ( n3732 & ~n3936 ) | ( n3935 & ~n3936 ) ;
  assign n3938 = n3786 ^ n3738 ^ x68 ;
  assign n3939 = n3837 ^ n3738 ^ 1'b0 ;
  assign n3940 = ( n3738 & n3938 ) | ( n3738 & ~n3939 ) | ( n3938 & ~n3939 ) ;
  assign n3941 = x23 & ~x64 ;
  assign n3942 = ( x23 & x105 ) | ( x23 & n3836 ) | ( x105 & n3836 ) ;
  assign n3943 = x106 | n3780 ;
  assign n3944 = ( x23 & n183 ) | ( x23 & n3943 ) | ( n183 & n3943 ) ;
  assign n3945 = ( x23 & n3942 ) | ( x23 & n3944 ) | ( n3942 & n3944 ) ;
  assign n3946 = ( x23 & n3941 ) | ( x23 & n3945 ) | ( n3941 & n3945 ) ;
  assign n3947 = ( ~n176 & n3818 ) | ( ~n176 & n3836 ) | ( n3818 & n3836 ) ;
  assign n3948 = ~n3836 & n3947 ;
  assign n3949 = n3946 | n3948 ;
  assign n3950 = ~x22 & x64 ;
  assign n3951 = n3950 ^ n3949 ^ x65 ;
  assign n3952 = ( x65 & n3950 ) | ( x65 & n3951 ) | ( n3950 & n3951 ) ;
  assign n3953 = n3952 ^ n3871 ^ x66 ;
  assign n3954 = ( x66 & n3952 ) | ( x66 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3955 = ( x67 & ~n3869 ) | ( x67 & n3954 ) | ( ~n3869 & n3954 ) ;
  assign n3956 = ( x68 & ~n3867 ) | ( x68 & n3955 ) | ( ~n3867 & n3955 ) ;
  assign n3957 = ( x69 & ~n3940 ) | ( x69 & n3956 ) | ( ~n3940 & n3956 ) ;
  assign n3958 = ( x70 & ~n3865 ) | ( x70 & n3957 ) | ( ~n3865 & n3957 ) ;
  assign n3959 = ( x71 & ~n3937 ) | ( x71 & n3958 ) | ( ~n3937 & n3958 ) ;
  assign n3960 = ( x72 & ~n3863 ) | ( x72 & n3959 ) | ( ~n3863 & n3959 ) ;
  assign n3961 = ( x73 & ~n3861 ) | ( x73 & n3960 ) | ( ~n3861 & n3960 ) ;
  assign n3962 = ( x74 & ~n3859 ) | ( x74 & n3961 ) | ( ~n3859 & n3961 ) ;
  assign n3963 = ( x75 & ~n3934 ) | ( x75 & n3962 ) | ( ~n3934 & n3962 ) ;
  assign n3964 = ( x76 & ~n3931 ) | ( x76 & n3963 ) | ( ~n3931 & n3963 ) ;
  assign n3965 = ( x77 & ~n3857 ) | ( x77 & n3964 ) | ( ~n3857 & n3964 ) ;
  assign n3966 = ( x78 & ~n3928 ) | ( x78 & n3965 ) | ( ~n3928 & n3965 ) ;
  assign n3967 = ( x79 & ~n3925 ) | ( x79 & n3966 ) | ( ~n3925 & n3966 ) ;
  assign n3968 = ( x80 & ~n3855 ) | ( x80 & n3967 ) | ( ~n3855 & n3967 ) ;
  assign n3969 = ( x81 & ~n3922 ) | ( x81 & n3968 ) | ( ~n3922 & n3968 ) ;
  assign n3970 = ( x82 & ~n3919 ) | ( x82 & n3969 ) | ( ~n3919 & n3969 ) ;
  assign n3971 = ( x83 & ~n3853 ) | ( x83 & n3970 ) | ( ~n3853 & n3970 ) ;
  assign n3972 = ( x84 & ~n3916 ) | ( x84 & n3971 ) | ( ~n3916 & n3971 ) ;
  assign n3973 = n3779 & n3837 ;
  assign n3974 = n322 | n3973 ;
  assign n3975 = ( x105 & ~n3943 ) | ( x105 & n3974 ) | ( ~n3943 & n3974 ) ;
  assign n3976 = ( x85 & ~n3851 ) | ( x85 & n3972 ) | ( ~n3851 & n3972 ) ;
  assign n3977 = ( x86 & ~n3849 ) | ( x86 & n3976 ) | ( ~n3849 & n3976 ) ;
  assign n3978 = ( x87 & ~n3913 ) | ( x87 & n3977 ) | ( ~n3913 & n3977 ) ;
  assign n3979 = n3957 ^ n3865 ^ x70 ;
  assign n3980 = n3960 ^ n3861 ^ x73 ;
  assign n3981 = n3961 ^ n3859 ^ x74 ;
  assign n3982 = n3964 ^ n3857 ^ x77 ;
  assign n3983 = n3966 ^ n3925 ^ x79 ;
  assign n3984 = n3967 ^ n3855 ^ x80 ;
  assign n3985 = ( n162 & n322 ) | ( n162 & n3779 ) | ( n322 & n3779 ) ;
  assign n3986 = n3977 ^ n3913 ^ x87 ;
  assign n3987 = n3965 ^ n3928 ^ x78 ;
  assign n3988 = ( x105 & n3943 ) | ( x105 & n3973 ) | ( n3943 & n3973 ) ;
  assign n3989 = ( n183 & n3975 ) | ( n183 & ~n3988 ) | ( n3975 & ~n3988 ) ;
  assign n3990 = ( x88 & ~n3910 ) | ( x88 & n3978 ) | ( ~n3910 & n3978 ) ;
  assign n3991 = n162 & n3974 ;
  assign n3992 = n3978 ^ n3910 ^ x88 ;
  assign n3993 = ( x89 & ~n3847 ) | ( x89 & n3990 ) | ( ~n3847 & n3990 ) ;
  assign n3994 = ( x90 & ~n3845 ) | ( x90 & n3993 ) | ( ~n3845 & n3993 ) ;
  assign n3995 = ( x91 & ~n3907 ) | ( x91 & n3994 ) | ( ~n3907 & n3994 ) ;
  assign n3996 = ( x92 & ~n3904 ) | ( x92 & n3995 ) | ( ~n3904 & n3995 ) ;
  assign n3997 = ( x93 & ~n3901 ) | ( x93 & n3996 ) | ( ~n3901 & n3996 ) ;
  assign n3998 = ( x94 & ~n3898 ) | ( x94 & n3997 ) | ( ~n3898 & n3997 ) ;
  assign n3999 = ( x95 & ~n3895 ) | ( x95 & n3998 ) | ( ~n3895 & n3998 ) ;
  assign n4000 = ( x96 & ~n3843 ) | ( x96 & n3999 ) | ( ~n3843 & n3999 ) ;
  assign n4001 = ( x97 & ~n3840 ) | ( x97 & n4000 ) | ( ~n3840 & n4000 ) ;
  assign n4002 = ( x98 & ~n3890 ) | ( x98 & n4001 ) | ( ~n3890 & n4001 ) ;
  assign n4003 = ( x99 & ~n3887 ) | ( x99 & n4002 ) | ( ~n3887 & n4002 ) ;
  assign n4004 = ( x100 & ~n3884 ) | ( x100 & n4003 ) | ( ~n3884 & n4003 ) ;
  assign n4005 = ( x101 & ~n3881 ) | ( x101 & n4004 ) | ( ~n3881 & n4004 ) ;
  assign n4006 = ( x102 & ~n3878 ) | ( x102 & n4005 ) | ( ~n3878 & n4005 ) ;
  assign n4007 = ( x103 & ~n3892 ) | ( x103 & n4006 ) | ( ~n3892 & n4006 ) ;
  assign n4008 = n4007 ^ n3874 ^ x104 ;
  assign n4009 = ( x104 & ~n3874 ) | ( x104 & n4007 ) | ( ~n3874 & n4007 ) ;
  assign n4010 = ( ~n3943 & n3989 ) | ( ~n3943 & n4009 ) | ( n3989 & n4009 ) ;
  assign n4011 = n3943 | n4010 ;
  assign n4012 = ( ~n3974 & n3991 ) | ( ~n3974 & n4011 ) | ( n3991 & n4011 ) ;
  assign n4013 = n4012 ^ n3874 ^ 1'b0 ;
  assign n4014 = ( n3874 & n4008 ) | ( n3874 & ~n4013 ) | ( n4008 & ~n4013 ) ;
  assign n4015 = n4001 ^ n3890 ^ x98 ;
  assign n4016 = n4012 ^ n3890 ^ 1'b0 ;
  assign n4017 = ( n3890 & n4015 ) | ( n3890 & ~n4016 ) | ( n4015 & ~n4016 ) ;
  assign n4018 = n3995 ^ n3904 ^ x92 ;
  assign n4019 = n4012 ^ n3904 ^ 1'b0 ;
  assign n4020 = ( n3904 & n4018 ) | ( n3904 & ~n4019 ) | ( n4018 & ~n4019 ) ;
  assign n4021 = n4012 ^ n3910 ^ 1'b0 ;
  assign n4022 = ( n3910 & n3992 ) | ( n3910 & ~n4021 ) | ( n3992 & ~n4021 ) ;
  assign n4023 = n4012 ^ n3913 ^ 1'b0 ;
  assign n4024 = ( n3913 & n3986 ) | ( n3913 & ~n4023 ) | ( n3986 & ~n4023 ) ;
  assign n4025 = n4012 ^ n3855 ^ 1'b0 ;
  assign n4026 = ( n3855 & n3984 ) | ( n3855 & ~n4025 ) | ( n3984 & ~n4025 ) ;
  assign n4027 = n4012 ^ n3925 ^ 1'b0 ;
  assign n4028 = ( n3925 & n3983 ) | ( n3925 & ~n4027 ) | ( n3983 & ~n4027 ) ;
  assign n4029 = n4012 ^ n3928 ^ 1'b0 ;
  assign n4030 = ( n3928 & n3987 ) | ( n3928 & ~n4029 ) | ( n3987 & ~n4029 ) ;
  assign n4031 = n4012 ^ n3857 ^ 1'b0 ;
  assign n4032 = ( n3857 & n3982 ) | ( n3857 & ~n4031 ) | ( n3982 & ~n4031 ) ;
  assign n4033 = n4012 ^ n3859 ^ 1'b0 ;
  assign n4034 = ( n3859 & n3981 ) | ( n3859 & ~n4033 ) | ( n3981 & ~n4033 ) ;
  assign n4035 = n4012 ^ n3861 ^ 1'b0 ;
  assign n4036 = ( n3861 & n3980 ) | ( n3861 & ~n4035 ) | ( n3980 & ~n4035 ) ;
  assign n4037 = n4012 ^ n3865 ^ 1'b0 ;
  assign n4038 = ( n3865 & n3979 ) | ( n3865 & ~n4037 ) | ( n3979 & ~n4037 ) ;
  assign n4039 = n4012 ^ n3953 ^ 1'b0 ;
  assign n4040 = ( n3871 & n3953 ) | ( n3871 & n4039 ) | ( n3953 & n4039 ) ;
  assign n4041 = n4012 ^ n3951 ^ 1'b0 ;
  assign n4042 = ( n3949 & n3951 ) | ( n3949 & n4041 ) | ( n3951 & n4041 ) ;
  assign n4043 = n322 | n4011 ;
  assign n4044 = ( n322 & n3985 ) | ( n322 & n4043 ) | ( n3985 & n4043 ) ;
  assign n4045 = n4006 ^ n3892 ^ x103 ;
  assign n4046 = n4005 ^ n3878 ^ x102 ;
  assign n4047 = n4012 ^ n3878 ^ 1'b0 ;
  assign n4048 = ( n3878 & n4046 ) | ( n3878 & ~n4047 ) | ( n4046 & ~n4047 ) ;
  assign n4049 = n4004 ^ n3881 ^ x101 ;
  assign n4050 = n4012 ^ n3881 ^ 1'b0 ;
  assign n4051 = ( n3881 & n4049 ) | ( n3881 & ~n4050 ) | ( n4049 & ~n4050 ) ;
  assign n4052 = n4003 ^ n3884 ^ x100 ;
  assign n4053 = n4012 ^ n3884 ^ 1'b0 ;
  assign n4054 = ( n3884 & n4052 ) | ( n3884 & ~n4053 ) | ( n4052 & ~n4053 ) ;
  assign n4055 = n4002 ^ n3887 ^ x99 ;
  assign n4056 = n4012 ^ n3887 ^ 1'b0 ;
  assign n4057 = ( n3887 & n4055 ) | ( n3887 & ~n4056 ) | ( n4055 & ~n4056 ) ;
  assign n4058 = n4000 ^ n3840 ^ x97 ;
  assign n4059 = n4012 ^ n3840 ^ 1'b0 ;
  assign n4060 = ( n3840 & n4058 ) | ( n3840 & ~n4059 ) | ( n4058 & ~n4059 ) ;
  assign n4061 = n3999 ^ n3843 ^ x96 ;
  assign n4062 = n4012 ^ n3843 ^ 1'b0 ;
  assign n4063 = ( n3843 & n4061 ) | ( n3843 & ~n4062 ) | ( n4061 & ~n4062 ) ;
  assign n4064 = n3998 ^ n3895 ^ x95 ;
  assign n4065 = n4012 ^ n3895 ^ 1'b0 ;
  assign n4066 = ( n3895 & n4064 ) | ( n3895 & ~n4065 ) | ( n4064 & ~n4065 ) ;
  assign n4067 = n3997 ^ n3898 ^ x94 ;
  assign n4068 = n4012 ^ n3898 ^ 1'b0 ;
  assign n4069 = ( n3898 & n4067 ) | ( n3898 & ~n4068 ) | ( n4067 & ~n4068 ) ;
  assign n4070 = n3996 ^ n3901 ^ x93 ;
  assign n4071 = n4012 ^ n3901 ^ 1'b0 ;
  assign n4072 = ( n3901 & n4070 ) | ( n3901 & ~n4071 ) | ( n4070 & ~n4071 ) ;
  assign n4073 = n3994 ^ n3907 ^ x91 ;
  assign n4074 = n4012 ^ n3907 ^ 1'b0 ;
  assign n4075 = ( n3907 & n4073 ) | ( n3907 & ~n4074 ) | ( n4073 & ~n4074 ) ;
  assign n4076 = n3993 ^ n3845 ^ x90 ;
  assign n4077 = n4012 ^ n3845 ^ 1'b0 ;
  assign n4078 = ( n3845 & n4076 ) | ( n3845 & ~n4077 ) | ( n4076 & ~n4077 ) ;
  assign n4079 = n3990 ^ n3847 ^ x89 ;
  assign n4080 = n4012 ^ n3847 ^ 1'b0 ;
  assign n4081 = ( n3847 & n4079 ) | ( n3847 & ~n4080 ) | ( n4079 & ~n4080 ) ;
  assign n4082 = n3976 ^ n3849 ^ x86 ;
  assign n4083 = n4012 ^ n3849 ^ 1'b0 ;
  assign n4084 = ( n3849 & n4082 ) | ( n3849 & ~n4083 ) | ( n4082 & ~n4083 ) ;
  assign n4085 = n3972 ^ n3851 ^ x85 ;
  assign n4086 = n4012 ^ n3851 ^ 1'b0 ;
  assign n4087 = ( n3851 & n4085 ) | ( n3851 & ~n4086 ) | ( n4085 & ~n4086 ) ;
  assign n4088 = n3971 ^ n3916 ^ x84 ;
  assign n4089 = n4012 ^ n3916 ^ 1'b0 ;
  assign n4090 = ( n3916 & n4088 ) | ( n3916 & ~n4089 ) | ( n4088 & ~n4089 ) ;
  assign n4091 = n3970 ^ n3853 ^ x83 ;
  assign n4092 = n4012 ^ n3853 ^ 1'b0 ;
  assign n4093 = ( n3853 & n4091 ) | ( n3853 & ~n4092 ) | ( n4091 & ~n4092 ) ;
  assign n4094 = n3969 ^ n3919 ^ x82 ;
  assign n4095 = n4012 ^ n3919 ^ 1'b0 ;
  assign n4096 = ( n3919 & n4094 ) | ( n3919 & ~n4095 ) | ( n4094 & ~n4095 ) ;
  assign n4097 = n3968 ^ n3922 ^ x81 ;
  assign n4098 = n4012 ^ n3892 ^ 1'b0 ;
  assign n4099 = ( n3892 & n4045 ) | ( n3892 & ~n4098 ) | ( n4045 & ~n4098 ) ;
  assign n4100 = n4012 ^ n3922 ^ 1'b0 ;
  assign n4101 = ( n3922 & n4097 ) | ( n3922 & ~n4100 ) | ( n4097 & ~n4100 ) ;
  assign n4102 = n3963 ^ n3931 ^ x76 ;
  assign n4103 = n4012 ^ n3931 ^ 1'b0 ;
  assign n4104 = ( n3931 & n4102 ) | ( n3931 & ~n4103 ) | ( n4102 & ~n4103 ) ;
  assign n4105 = n3962 ^ n3934 ^ x75 ;
  assign n4106 = n4012 ^ n3934 ^ 1'b0 ;
  assign n4107 = ( n3934 & n4105 ) | ( n3934 & ~n4106 ) | ( n4105 & ~n4106 ) ;
  assign n4108 = n3959 ^ n3863 ^ x72 ;
  assign n4109 = n4012 ^ n3863 ^ 1'b0 ;
  assign n4110 = ( n3863 & n4108 ) | ( n3863 & ~n4109 ) | ( n4108 & ~n4109 ) ;
  assign n4111 = n3958 ^ n3937 ^ x71 ;
  assign n4112 = n4012 ^ n3937 ^ 1'b0 ;
  assign n4113 = ( n3937 & n4111 ) | ( n3937 & ~n4112 ) | ( n4111 & ~n4112 ) ;
  assign n4114 = n3956 ^ n3940 ^ x69 ;
  assign n4115 = n4012 ^ n3940 ^ 1'b0 ;
  assign n4116 = ( n3940 & n4114 ) | ( n3940 & ~n4115 ) | ( n4114 & ~n4115 ) ;
  assign n4117 = n3955 ^ n3867 ^ x68 ;
  assign n4118 = n4012 ^ n3867 ^ 1'b0 ;
  assign n4119 = ( n3867 & n4117 ) | ( n3867 & ~n4118 ) | ( n4117 & ~n4118 ) ;
  assign n4120 = n3954 ^ n3869 ^ x67 ;
  assign n4121 = n4012 ^ n3869 ^ 1'b0 ;
  assign n4122 = ( n3869 & n4120 ) | ( n3869 & ~n4121 ) | ( n4120 & ~n4121 ) ;
  assign n4123 = x64 & n4012 ;
  assign n4124 = ~x21 & x64 ;
  assign n4125 = n4123 ^ x64 ^ x22 ;
  assign n4126 = n4125 ^ n4124 ^ x65 ;
  assign n4127 = ( x65 & n4124 ) | ( x65 & n4126 ) | ( n4124 & n4126 ) ;
  assign n4128 = n4127 ^ n4042 ^ x66 ;
  assign n4129 = ( x66 & n4127 ) | ( x66 & n4128 ) | ( n4127 & n4128 ) ;
  assign n4130 = ( x67 & ~n4040 ) | ( x67 & n4129 ) | ( ~n4040 & n4129 ) ;
  assign n4131 = ( x68 & ~n4122 ) | ( x68 & n4130 ) | ( ~n4122 & n4130 ) ;
  assign n4132 = ( x69 & ~n4119 ) | ( x69 & n4131 ) | ( ~n4119 & n4131 ) ;
  assign n4133 = ( x70 & ~n4116 ) | ( x70 & n4132 ) | ( ~n4116 & n4132 ) ;
  assign n4134 = ( x71 & ~n4038 ) | ( x71 & n4133 ) | ( ~n4038 & n4133 ) ;
  assign n4135 = ( x72 & ~n4113 ) | ( x72 & n4134 ) | ( ~n4113 & n4134 ) ;
  assign n4136 = ( x73 & ~n4110 ) | ( x73 & n4135 ) | ( ~n4110 & n4135 ) ;
  assign n4137 = ( x74 & ~n4036 ) | ( x74 & n4136 ) | ( ~n4036 & n4136 ) ;
  assign n4138 = ( x75 & ~n4034 ) | ( x75 & n4137 ) | ( ~n4034 & n4137 ) ;
  assign n4139 = ( x76 & ~n4107 ) | ( x76 & n4138 ) | ( ~n4107 & n4138 ) ;
  assign n4140 = ( x77 & ~n4104 ) | ( x77 & n4139 ) | ( ~n4104 & n4139 ) ;
  assign n4141 = ( x78 & ~n4032 ) | ( x78 & n4140 ) | ( ~n4032 & n4140 ) ;
  assign n4142 = ( x79 & ~n4030 ) | ( x79 & n4141 ) | ( ~n4030 & n4141 ) ;
  assign n4143 = ( x80 & ~n4028 ) | ( x80 & n4142 ) | ( ~n4028 & n4142 ) ;
  assign n4144 = ( x81 & ~n4026 ) | ( x81 & n4143 ) | ( ~n4026 & n4143 ) ;
  assign n4145 = ( x82 & ~n4101 ) | ( x82 & n4144 ) | ( ~n4101 & n4144 ) ;
  assign n4146 = ( x83 & ~n4096 ) | ( x83 & n4145 ) | ( ~n4096 & n4145 ) ;
  assign n4147 = ( x84 & ~n4093 ) | ( x84 & n4146 ) | ( ~n4093 & n4146 ) ;
  assign n4148 = ( x85 & ~n4090 ) | ( x85 & n4147 ) | ( ~n4090 & n4147 ) ;
  assign n4149 = ( x86 & ~n4087 ) | ( x86 & n4148 ) | ( ~n4087 & n4148 ) ;
  assign n4150 = ( x87 & ~n4084 ) | ( x87 & n4149 ) | ( ~n4084 & n4149 ) ;
  assign n4151 = ( x88 & ~n4024 ) | ( x88 & n4150 ) | ( ~n4024 & n4150 ) ;
  assign n4152 = ( x89 & ~n4022 ) | ( x89 & n4151 ) | ( ~n4022 & n4151 ) ;
  assign n4153 = ( x90 & ~n4081 ) | ( x90 & n4152 ) | ( ~n4081 & n4152 ) ;
  assign n4154 = ( x91 & ~n4078 ) | ( x91 & n4153 ) | ( ~n4078 & n4153 ) ;
  assign n4155 = ( x92 & ~n4075 ) | ( x92 & n4154 ) | ( ~n4075 & n4154 ) ;
  assign n4156 = n4146 ^ n4093 ^ x84 ;
  assign n4157 = n4154 ^ n4075 ^ x92 ;
  assign n4158 = n4148 ^ n4087 ^ x86 ;
  assign n4159 = n4138 ^ n4107 ^ x76 ;
  assign n4160 = n4151 ^ n4022 ^ x89 ;
  assign n4161 = n4153 ^ n4078 ^ x91 ;
  assign n4162 = n4137 ^ n4034 ^ x75 ;
  assign n4163 = n4130 ^ n4122 ^ x68 ;
  assign n4164 = n4135 ^ n4110 ^ x73 ;
  assign n4165 = n4139 ^ n4104 ^ x77 ;
  assign n4166 = ( x93 & ~n4020 ) | ( x93 & n4155 ) | ( ~n4020 & n4155 ) ;
  assign n4167 = ( x94 & ~n4072 ) | ( x94 & n4166 ) | ( ~n4072 & n4166 ) ;
  assign n4168 = ( x95 & ~n4069 ) | ( x95 & n4167 ) | ( ~n4069 & n4167 ) ;
  assign n4169 = ( x96 & ~n4066 ) | ( x96 & n4168 ) | ( ~n4066 & n4168 ) ;
  assign n4170 = ( x97 & ~n4063 ) | ( x97 & n4169 ) | ( ~n4063 & n4169 ) ;
  assign n4171 = ( x98 & ~n4060 ) | ( x98 & n4170 ) | ( ~n4060 & n4170 ) ;
  assign n4172 = ( x99 & ~n4017 ) | ( x99 & n4171 ) | ( ~n4017 & n4171 ) ;
  assign n4173 = ( x100 & ~n4057 ) | ( x100 & n4172 ) | ( ~n4057 & n4172 ) ;
  assign n4174 = ( x101 & ~n4054 ) | ( x101 & n4173 ) | ( ~n4054 & n4173 ) ;
  assign n4175 = ( x102 & ~n4051 ) | ( x102 & n4174 ) | ( ~n4051 & n4174 ) ;
  assign n4176 = ( x103 & ~n4048 ) | ( x103 & n4175 ) | ( ~n4048 & n4175 ) ;
  assign n4177 = ( x104 & ~n4099 ) | ( x104 & n4176 ) | ( ~n4099 & n4176 ) ;
  assign n4178 = ( x105 & ~n4014 ) | ( x105 & n4177 ) | ( ~n4014 & n4177 ) ;
  assign n4179 = ( x106 & ~n4044 ) | ( x106 & n4178 ) | ( ~n4044 & n4178 ) ;
  assign n4180 = n177 | n4179 ;
  assign n4181 = n4175 ^ n4048 ^ x103 ;
  assign n4182 = n4180 ^ n4048 ^ 1'b0 ;
  assign n4183 = ( n4048 & n4181 ) | ( n4048 & ~n4182 ) | ( n4181 & ~n4182 ) ;
  assign n4184 = n4170 ^ n4060 ^ x98 ;
  assign n4185 = n4180 ^ n4060 ^ 1'b0 ;
  assign n4186 = ( n4060 & n4184 ) | ( n4060 & ~n4185 ) | ( n4184 & ~n4185 ) ;
  assign n4187 = n4169 ^ n4063 ^ x97 ;
  assign n4188 = n4180 ^ n4063 ^ 1'b0 ;
  assign n4189 = ( n4063 & n4187 ) | ( n4063 & ~n4188 ) | ( n4187 & ~n4188 ) ;
  assign n4190 = n4155 ^ n4020 ^ x93 ;
  assign n4191 = n4180 ^ n4020 ^ 1'b0 ;
  assign n4192 = ( n4020 & n4190 ) | ( n4020 & ~n4191 ) | ( n4190 & ~n4191 ) ;
  assign n4193 = n4180 ^ n4075 ^ 1'b0 ;
  assign n4194 = ( n4075 & n4157 ) | ( n4075 & ~n4193 ) | ( n4157 & ~n4193 ) ;
  assign n4195 = n4180 ^ n4078 ^ 1'b0 ;
  assign n4196 = ( n4078 & n4161 ) | ( n4078 & ~n4195 ) | ( n4161 & ~n4195 ) ;
  assign n4197 = n4180 ^ n4022 ^ 1'b0 ;
  assign n4198 = ( n4022 & n4160 ) | ( n4022 & ~n4197 ) | ( n4160 & ~n4197 ) ;
  assign n4199 = n4180 ^ n4087 ^ 1'b0 ;
  assign n4200 = ( n4087 & n4158 ) | ( n4087 & ~n4199 ) | ( n4158 & ~n4199 ) ;
  assign n4201 = n4180 ^ n4093 ^ 1'b0 ;
  assign n4202 = ( n4093 & n4156 ) | ( n4093 & ~n4201 ) | ( n4156 & ~n4201 ) ;
  assign n4203 = n4180 ^ n4104 ^ 1'b0 ;
  assign n4204 = ( n4104 & n4165 ) | ( n4104 & ~n4203 ) | ( n4165 & ~n4203 ) ;
  assign n4205 = n4180 ^ n4107 ^ 1'b0 ;
  assign n4206 = ( n4107 & n4159 ) | ( n4107 & ~n4205 ) | ( n4159 & ~n4205 ) ;
  assign n4207 = n4180 ^ n4034 ^ 1'b0 ;
  assign n4208 = ( n4034 & n4162 ) | ( n4034 & ~n4207 ) | ( n4162 & ~n4207 ) ;
  assign n4209 = n4180 ^ n4110 ^ 1'b0 ;
  assign n4210 = ( n4110 & n4164 ) | ( n4110 & ~n4209 ) | ( n4164 & ~n4209 ) ;
  assign n4211 = n4133 ^ n4038 ^ x71 ;
  assign n4212 = n4180 ^ n4038 ^ 1'b0 ;
  assign n4213 = ( n4038 & n4211 ) | ( n4038 & ~n4212 ) | ( n4211 & ~n4212 ) ;
  assign n4214 = n4180 ^ n4122 ^ 1'b0 ;
  assign n4215 = ( n4122 & n4163 ) | ( n4122 & ~n4214 ) | ( n4163 & ~n4214 ) ;
  assign n4216 = n4180 ^ n4128 ^ 1'b0 ;
  assign n4217 = ( n4042 & n4128 ) | ( n4042 & n4216 ) | ( n4128 & n4216 ) ;
  assign n4218 = ( ~x21 & x64 ) | ( ~x21 & n4179 ) | ( x64 & n4179 ) ;
  assign n4219 = n4143 ^ n4026 ^ x81 ;
  assign n4220 = n4171 ^ n4017 ^ x99 ;
  assign n4221 = x64 & ~n4218 ;
  assign n4222 = ( ~x107 & n3273 ) | ( ~x107 & n4221 ) | ( n3273 & n4221 ) ;
  assign n4223 = ~n3273 & n4222 ;
  assign n4224 = n4177 ^ n4014 ^ x105 ;
  assign n4225 = n4134 ^ n4113 ^ x72 ;
  assign n4226 = n4124 & ~n4180 ;
  assign n4227 = ( x21 & ~n4223 ) | ( x21 & n4226 ) | ( ~n4223 & n4226 ) ;
  assign n4228 = n4180 ^ n4026 ^ 1'b0 ;
  assign n4229 = ( n4026 & n4219 ) | ( n4026 & ~n4228 ) | ( n4219 & ~n4228 ) ;
  assign n4230 = n4180 ^ n4113 ^ 1'b0 ;
  assign n4231 = n4180 ^ n4084 ^ 1'b0 ;
  assign n4232 = ( n4113 & n4225 ) | ( n4113 & ~n4230 ) | ( n4225 & ~n4230 ) ;
  assign n4233 = n4180 ^ n4066 ^ 1'b0 ;
  assign n4234 = n4180 ^ n4017 ^ 1'b0 ;
  assign n4235 = n4145 ^ n4096 ^ x83 ;
  assign n4236 = n4168 ^ n4066 ^ x96 ;
  assign n4237 = ( n4017 & n4220 ) | ( n4017 & ~n4234 ) | ( n4220 & ~n4234 ) ;
  assign n4238 = n4149 ^ n4084 ^ x87 ;
  assign n4239 = ( n4084 & ~n4231 ) | ( n4084 & n4238 ) | ( ~n4231 & n4238 ) ;
  assign n4240 = n4166 ^ n4072 ^ x94 ;
  assign n4241 = ( n4066 & ~n4233 ) | ( n4066 & n4236 ) | ( ~n4233 & n4236 ) ;
  assign n4242 = n4224 ^ n4180 ^ 1'b0 ;
  assign n4243 = n4141 ^ n4030 ^ x79 ;
  assign n4244 = ( n4014 & n4224 ) | ( n4014 & n4242 ) | ( n4224 & n4242 ) ;
  assign n4245 = n4180 ^ n4030 ^ 1'b0 ;
  assign n4246 = n4180 ^ n4072 ^ 1'b0 ;
  assign n4247 = ( n4072 & n4240 ) | ( n4072 & ~n4246 ) | ( n4240 & ~n4246 ) ;
  assign n4248 = n4136 ^ n4036 ^ x74 ;
  assign n4249 = n4167 ^ n4069 ^ x95 ;
  assign n4250 = n4180 ^ n4040 ^ 1'b0 ;
  assign n4251 = n4180 ^ n4069 ^ 1'b0 ;
  assign n4252 = n4152 ^ n4081 ^ x90 ;
  assign n4253 = n4129 ^ n4040 ^ x67 ;
  assign n4254 = n4131 ^ n4119 ^ x69 ;
  assign n4255 = n4180 ^ n4081 ^ 1'b0 ;
  assign n4256 = ( n4081 & n4252 ) | ( n4081 & ~n4255 ) | ( n4252 & ~n4255 ) ;
  assign n4257 = ( n4040 & ~n4250 ) | ( n4040 & n4253 ) | ( ~n4250 & n4253 ) ;
  assign n4258 = n4172 ^ n4057 ^ x100 ;
  assign n4259 = n4150 ^ n4024 ^ x88 ;
  assign n4260 = n4180 ^ n4051 ^ 1'b0 ;
  assign n4261 = n4174 ^ n4051 ^ x102 ;
  assign n4262 = ( n4051 & ~n4260 ) | ( n4051 & n4261 ) | ( ~n4260 & n4261 ) ;
  assign n4263 = n4144 ^ n4101 ^ x82 ;
  assign n4264 = n4180 ^ n4028 ^ 1'b0 ;
  assign n4265 = n4176 ^ n4099 ^ x104 ;
  assign n4266 = n4173 ^ n4054 ^ x101 ;
  assign n4267 = n4180 ^ n4032 ^ 1'b0 ;
  assign n4268 = n4180 ^ n4054 ^ 1'b0 ;
  assign n4269 = ( n4054 & n4266 ) | ( n4054 & ~n4268 ) | ( n4266 & ~n4268 ) ;
  assign n4270 = ( n4030 & n4243 ) | ( n4030 & ~n4245 ) | ( n4243 & ~n4245 ) ;
  assign n4271 = n4132 ^ n4116 ^ x70 ;
  assign n4272 = n4180 ^ n4116 ^ 1'b0 ;
  assign n4273 = ( n4116 & n4271 ) | ( n4116 & ~n4272 ) | ( n4271 & ~n4272 ) ;
  assign n4274 = n4180 ^ n4024 ^ 1'b0 ;
  assign n4275 = n4180 ^ n4096 ^ 1'b0 ;
  assign n4276 = ( n4096 & n4235 ) | ( n4096 & ~n4275 ) | ( n4235 & ~n4275 ) ;
  assign n4277 = n4140 ^ n4032 ^ x78 ;
  assign n4278 = n4180 ^ n4119 ^ 1'b0 ;
  assign n4279 = ( n4069 & n4249 ) | ( n4069 & ~n4251 ) | ( n4249 & ~n4251 ) ;
  assign n4280 = n4142 ^ n4028 ^ x80 ;
  assign n4281 = ( n4032 & ~n4267 ) | ( n4032 & n4277 ) | ( ~n4267 & n4277 ) ;
  assign n4282 = n4180 ^ n4101 ^ 1'b0 ;
  assign n4283 = n4180 ^ n4090 ^ 1'b0 ;
  assign n4284 = ( n4119 & n4254 ) | ( n4119 & ~n4278 ) | ( n4254 & ~n4278 ) ;
  assign n4285 = ( n4024 & n4259 ) | ( n4024 & ~n4274 ) | ( n4259 & ~n4274 ) ;
  assign n4286 = n4147 ^ n4090 ^ x85 ;
  assign n4287 = ( n4090 & ~n4283 ) | ( n4090 & n4286 ) | ( ~n4283 & n4286 ) ;
  assign n4288 = n4180 ^ n4057 ^ 1'b0 ;
  assign n4289 = ( n4057 & n4258 ) | ( n4057 & ~n4288 ) | ( n4258 & ~n4288 ) ;
  assign n4290 = n4180 ^ n4036 ^ 1'b0 ;
  assign n4291 = n4180 ^ n4099 ^ 1'b0 ;
  assign n4292 = ( n4028 & ~n4264 ) | ( n4028 & n4280 ) | ( ~n4264 & n4280 ) ;
  assign n4293 = ( n4101 & n4263 ) | ( n4101 & ~n4282 ) | ( n4263 & ~n4282 ) ;
  assign n4294 = ( n4099 & n4265 ) | ( n4099 & ~n4291 ) | ( n4265 & ~n4291 ) ;
  assign n4295 = n4180 ^ n4126 ^ 1'b0 ;
  assign n4296 = ( n4125 & n4126 ) | ( n4125 & n4295 ) | ( n4126 & n4295 ) ;
  assign n4297 = ( n4036 & n4248 ) | ( n4036 & ~n4290 ) | ( n4248 & ~n4290 ) ;
  assign n4298 = ~x20 & x64 ;
  assign n4299 = n4298 ^ n4227 ^ x65 ;
  assign n4300 = ( x65 & n4298 ) | ( x65 & n4299 ) | ( n4298 & n4299 ) ;
  assign n4301 = n4300 ^ n4296 ^ x66 ;
  assign n4302 = ( x66 & n4300 ) | ( x66 & n4301 ) | ( n4300 & n4301 ) ;
  assign n4303 = ( x67 & ~n4217 ) | ( x67 & n4302 ) | ( ~n4217 & n4302 ) ;
  assign n4304 = ( x68 & ~n4257 ) | ( x68 & n4303 ) | ( ~n4257 & n4303 ) ;
  assign n4305 = ( x69 & ~n4215 ) | ( x69 & n4304 ) | ( ~n4215 & n4304 ) ;
  assign n4306 = ( x70 & ~n4284 ) | ( x70 & n4305 ) | ( ~n4284 & n4305 ) ;
  assign n4307 = ( x71 & ~n4273 ) | ( x71 & n4306 ) | ( ~n4273 & n4306 ) ;
  assign n4308 = ( x72 & ~n4213 ) | ( x72 & n4307 ) | ( ~n4213 & n4307 ) ;
  assign n4309 = ( x73 & ~n4232 ) | ( x73 & n4308 ) | ( ~n4232 & n4308 ) ;
  assign n4310 = ( x74 & ~n4210 ) | ( x74 & n4309 ) | ( ~n4210 & n4309 ) ;
  assign n4311 = n4044 & n4180 ;
  assign n4312 = ( x75 & ~n4297 ) | ( x75 & n4310 ) | ( ~n4297 & n4310 ) ;
  assign n4313 = ( x76 & ~n4208 ) | ( x76 & n4312 ) | ( ~n4208 & n4312 ) ;
  assign n4314 = n322 | n4311 ;
  assign n4315 = ( x77 & ~n4206 ) | ( x77 & n4313 ) | ( ~n4206 & n4313 ) ;
  assign n4316 = ( x78 & ~n4204 ) | ( x78 & n4315 ) | ( ~n4204 & n4315 ) ;
  assign n4317 = ( x79 & ~n4281 ) | ( x79 & n4316 ) | ( ~n4281 & n4316 ) ;
  assign n4318 = ( x80 & ~n4270 ) | ( x80 & n4317 ) | ( ~n4270 & n4317 ) ;
  assign n4319 = ( x81 & ~n4292 ) | ( x81 & n4318 ) | ( ~n4292 & n4318 ) ;
  assign n4320 = ( x82 & ~n4229 ) | ( x82 & n4319 ) | ( ~n4229 & n4319 ) ;
  assign n4321 = ( x83 & ~n4293 ) | ( x83 & n4320 ) | ( ~n4293 & n4320 ) ;
  assign n4322 = ( x84 & ~n4276 ) | ( x84 & n4321 ) | ( ~n4276 & n4321 ) ;
  assign n4323 = ( x85 & ~n4202 ) | ( x85 & n4322 ) | ( ~n4202 & n4322 ) ;
  assign n4324 = ( x86 & ~n4287 ) | ( x86 & n4323 ) | ( ~n4287 & n4323 ) ;
  assign n4325 = ( x87 & ~n4200 ) | ( x87 & n4324 ) | ( ~n4200 & n4324 ) ;
  assign n4326 = ( x88 & ~n4239 ) | ( x88 & n4325 ) | ( ~n4239 & n4325 ) ;
  assign n4327 = ( x89 & ~n4285 ) | ( x89 & n4326 ) | ( ~n4285 & n4326 ) ;
  assign n4328 = ( x90 & ~n4198 ) | ( x90 & n4327 ) | ( ~n4198 & n4327 ) ;
  assign n4329 = n177 & n4044 ;
  assign n4330 = ( x91 & ~n4256 ) | ( x91 & n4328 ) | ( ~n4256 & n4328 ) ;
  assign n4331 = ( x92 & ~n4196 ) | ( x92 & n4330 ) | ( ~n4196 & n4330 ) ;
  assign n4332 = ( x93 & ~n4194 ) | ( x93 & n4331 ) | ( ~n4194 & n4331 ) ;
  assign n4333 = n177 & n4314 ;
  assign n4334 = n4309 ^ n4210 ^ x74 ;
  assign n4335 = ( x107 & n3273 ) | ( x107 & ~n4311 ) | ( n3273 & ~n4311 ) ;
  assign n4336 = n4312 ^ n4208 ^ x76 ;
  assign n4337 = n4310 ^ n4297 ^ x75 ;
  assign n4338 = n4306 ^ n4273 ^ x71 ;
  assign n4339 = n4308 ^ n4232 ^ x73 ;
  assign n4340 = n4307 ^ n4213 ^ x72 ;
  assign n4341 = n4303 ^ n4257 ^ x68 ;
  assign n4342 = n4305 ^ n4284 ^ x70 ;
  assign n4343 = ( x94 & ~n4192 ) | ( x94 & n4332 ) | ( ~n4192 & n4332 ) ;
  assign n4344 = ( x95 & ~n4247 ) | ( x95 & n4343 ) | ( ~n4247 & n4343 ) ;
  assign n4345 = ( x96 & ~n4279 ) | ( x96 & n4344 ) | ( ~n4279 & n4344 ) ;
  assign n4346 = ( x97 & ~n4241 ) | ( x97 & n4345 ) | ( ~n4241 & n4345 ) ;
  assign n4347 = ( ~x107 & n3273 ) | ( ~x107 & n4314 ) | ( n3273 & n4314 ) ;
  assign n4348 = ( x98 & ~n4189 ) | ( x98 & n4346 ) | ( ~n4189 & n4346 ) ;
  assign n4349 = ( x99 & ~n4186 ) | ( x99 & n4348 ) | ( ~n4186 & n4348 ) ;
  assign n4350 = ( x100 & ~n4237 ) | ( x100 & n4349 ) | ( ~n4237 & n4349 ) ;
  assign n4351 = ( x101 & ~n4289 ) | ( x101 & n4350 ) | ( ~n4289 & n4350 ) ;
  assign n4352 = ( x102 & ~n4269 ) | ( x102 & n4351 ) | ( ~n4269 & n4351 ) ;
  assign n4353 = ( x103 & ~n4262 ) | ( x103 & n4352 ) | ( ~n4262 & n4352 ) ;
  assign n4354 = ( x104 & ~n4183 ) | ( x104 & n4353 ) | ( ~n4183 & n4353 ) ;
  assign n4355 = ( x105 & ~n4294 ) | ( x105 & n4354 ) | ( ~n4294 & n4354 ) ;
  assign n4356 = ( x106 & ~n4244 ) | ( x106 & n4355 ) | ( ~n4244 & n4355 ) ;
  assign n4357 = n4355 ^ n4244 ^ x106 ;
  assign n4358 = ( n4335 & n4347 ) | ( n4335 & ~n4356 ) | ( n4347 & ~n4356 ) ;
  assign n4359 = n4356 | n4358 ;
  assign n4360 = ( ~n4314 & n4333 ) | ( ~n4314 & n4359 ) | ( n4333 & n4359 ) ;
  assign n4361 = n4360 ^ n4244 ^ 1'b0 ;
  assign n4362 = ( n4244 & n4357 ) | ( n4244 & ~n4361 ) | ( n4357 & ~n4361 ) ;
  assign n4363 = n4354 ^ n4294 ^ x105 ;
  assign n4364 = n4360 ^ n4294 ^ 1'b0 ;
  assign n4365 = ( n4294 & n4363 ) | ( n4294 & ~n4364 ) | ( n4363 & ~n4364 ) ;
  assign n4366 = n4353 ^ n4183 ^ x104 ;
  assign n4367 = n4360 ^ n4183 ^ 1'b0 ;
  assign n4368 = ( n4183 & n4366 ) | ( n4183 & ~n4367 ) | ( n4366 & ~n4367 ) ;
  assign n4369 = n4352 ^ n4262 ^ x103 ;
  assign n4370 = n4360 ^ n4262 ^ 1'b0 ;
  assign n4371 = ( n4262 & n4369 ) | ( n4262 & ~n4370 ) | ( n4369 & ~n4370 ) ;
  assign n4372 = n4351 ^ n4269 ^ x102 ;
  assign n4373 = n4360 ^ n4269 ^ 1'b0 ;
  assign n4374 = ( n4269 & n4372 ) | ( n4269 & ~n4373 ) | ( n4372 & ~n4373 ) ;
  assign n4375 = n4360 ^ n4208 ^ 1'b0 ;
  assign n4376 = ( n4208 & n4336 ) | ( n4208 & ~n4375 ) | ( n4336 & ~n4375 ) ;
  assign n4377 = n4360 ^ n4297 ^ 1'b0 ;
  assign n4378 = ( n4297 & n4337 ) | ( n4297 & ~n4377 ) | ( n4337 & ~n4377 ) ;
  assign n4379 = n4360 ^ n4210 ^ 1'b0 ;
  assign n4380 = ( n4210 & n4334 ) | ( n4210 & ~n4379 ) | ( n4334 & ~n4379 ) ;
  assign n4381 = n4360 ^ n4232 ^ 1'b0 ;
  assign n4382 = ( n4232 & n4339 ) | ( n4232 & ~n4381 ) | ( n4339 & ~n4381 ) ;
  assign n4383 = n4360 ^ n4213 ^ 1'b0 ;
  assign n4384 = ( n4213 & n4340 ) | ( n4213 & ~n4383 ) | ( n4340 & ~n4383 ) ;
  assign n4385 = n4360 ^ n4273 ^ 1'b0 ;
  assign n4386 = ( n4273 & n4338 ) | ( n4273 & ~n4385 ) | ( n4338 & ~n4385 ) ;
  assign n4387 = n4360 ^ n4284 ^ 1'b0 ;
  assign n4388 = ( n4284 & n4342 ) | ( n4284 & ~n4387 ) | ( n4342 & ~n4387 ) ;
  assign n4389 = n4360 ^ n4257 ^ 1'b0 ;
  assign n4390 = ( n4257 & n4341 ) | ( n4257 & ~n4389 ) | ( n4341 & ~n4389 ) ;
  assign n4391 = n4360 ^ n4301 ^ 1'b0 ;
  assign n4392 = ( n4296 & n4301 ) | ( n4296 & n4391 ) | ( n4301 & n4391 ) ;
  assign n4393 = n4360 ^ n4299 ^ 1'b0 ;
  assign n4394 = ( n4227 & n4299 ) | ( n4227 & n4393 ) | ( n4299 & n4393 ) ;
  assign n4395 = n4329 & n4359 ;
  assign n4396 = n4350 ^ n4289 ^ x101 ;
  assign n4397 = n4360 ^ n4289 ^ 1'b0 ;
  assign n4398 = ( n4289 & n4396 ) | ( n4289 & ~n4397 ) | ( n4396 & ~n4397 ) ;
  assign n4399 = n4324 ^ n4200 ^ x87 ;
  assign n4400 = n4360 ^ n4200 ^ 1'b0 ;
  assign n4401 = ( n4200 & n4399 ) | ( n4200 & ~n4400 ) | ( n4399 & ~n4400 ) ;
  assign n4402 = n4323 ^ n4287 ^ x86 ;
  assign n4403 = n4360 ^ n4287 ^ 1'b0 ;
  assign n4404 = ( n4287 & n4402 ) | ( n4287 & ~n4403 ) | ( n4402 & ~n4403 ) ;
  assign n4405 = n4322 ^ n4202 ^ x85 ;
  assign n4406 = n4360 ^ n4202 ^ 1'b0 ;
  assign n4407 = ( n4202 & n4405 ) | ( n4202 & ~n4406 ) | ( n4405 & ~n4406 ) ;
  assign n4408 = n4321 ^ n4276 ^ x84 ;
  assign n4409 = n4360 ^ n4276 ^ 1'b0 ;
  assign n4410 = ( n4276 & n4408 ) | ( n4276 & ~n4409 ) | ( n4408 & ~n4409 ) ;
  assign n4411 = n4320 ^ n4293 ^ x83 ;
  assign n4412 = n4360 ^ n4293 ^ 1'b0 ;
  assign n4413 = ( n4293 & n4411 ) | ( n4293 & ~n4412 ) | ( n4411 & ~n4412 ) ;
  assign n4414 = n4319 ^ n4229 ^ x82 ;
  assign n4415 = n4360 ^ n4229 ^ 1'b0 ;
  assign n4416 = ( n4229 & n4414 ) | ( n4229 & ~n4415 ) | ( n4414 & ~n4415 ) ;
  assign n4417 = n4318 ^ n4292 ^ x81 ;
  assign n4418 = n4360 ^ n4292 ^ 1'b0 ;
  assign n4419 = ( n4292 & n4417 ) | ( n4292 & ~n4418 ) | ( n4417 & ~n4418 ) ;
  assign n4420 = n4317 ^ n4270 ^ x80 ;
  assign n4421 = n4360 ^ n4270 ^ 1'b0 ;
  assign n4422 = ( n4270 & n4420 ) | ( n4270 & ~n4421 ) | ( n4420 & ~n4421 ) ;
  assign n4423 = n4316 ^ n4281 ^ x79 ;
  assign n4424 = n4360 ^ n4281 ^ 1'b0 ;
  assign n4425 = ( n4281 & n4423 ) | ( n4281 & ~n4424 ) | ( n4423 & ~n4424 ) ;
  assign n4426 = n4315 ^ n4204 ^ x78 ;
  assign n4427 = n4360 ^ n4204 ^ 1'b0 ;
  assign n4428 = ( n4204 & n4426 ) | ( n4204 & ~n4427 ) | ( n4426 & ~n4427 ) ;
  assign n4429 = n4313 ^ n4206 ^ x77 ;
  assign n4430 = n4360 ^ n4206 ^ 1'b0 ;
  assign n4431 = ( n4206 & n4429 ) | ( n4206 & ~n4430 ) | ( n4429 & ~n4430 ) ;
  assign n4432 = n4304 ^ n4215 ^ x69 ;
  assign n4433 = n4360 ^ n4215 ^ 1'b0 ;
  assign n4434 = ( n4215 & n4432 ) | ( n4215 & ~n4433 ) | ( n4432 & ~n4433 ) ;
  assign n4435 = n4302 ^ n4217 ^ x67 ;
  assign n4436 = n4360 ^ n4217 ^ 1'b0 ;
  assign n4437 = ( n4217 & n4435 ) | ( n4217 & ~n4436 ) | ( n4435 & ~n4436 ) ;
  assign n4438 = n4349 ^ n4237 ^ x100 ;
  assign n4439 = n4360 ^ n4237 ^ 1'b0 ;
  assign n4440 = ( n4237 & n4438 ) | ( n4237 & ~n4439 ) | ( n4438 & ~n4439 ) ;
  assign n4441 = n4348 ^ n4186 ^ x99 ;
  assign n4442 = n4360 ^ n4186 ^ 1'b0 ;
  assign n4443 = ( n4186 & n4441 ) | ( n4186 & ~n4442 ) | ( n4441 & ~n4442 ) ;
  assign n4444 = n4346 ^ n4189 ^ x98 ;
  assign n4445 = n4360 ^ n4189 ^ 1'b0 ;
  assign n4446 = ( n4189 & n4444 ) | ( n4189 & ~n4445 ) | ( n4444 & ~n4445 ) ;
  assign n4447 = n4345 ^ n4241 ^ x97 ;
  assign n4448 = n4360 ^ n4241 ^ 1'b0 ;
  assign n4449 = ( n4241 & n4447 ) | ( n4241 & ~n4448 ) | ( n4447 & ~n4448 ) ;
  assign n4450 = n4344 ^ n4279 ^ x96 ;
  assign n4451 = n4360 ^ n4279 ^ 1'b0 ;
  assign n4452 = ( n4279 & n4450 ) | ( n4279 & ~n4451 ) | ( n4450 & ~n4451 ) ;
  assign n4453 = n4343 ^ n4247 ^ x95 ;
  assign n4454 = n4360 ^ n4247 ^ 1'b0 ;
  assign n4455 = ( n4247 & n4453 ) | ( n4247 & ~n4454 ) | ( n4453 & ~n4454 ) ;
  assign n4456 = n4332 ^ n4192 ^ x94 ;
  assign n4457 = n4360 ^ n4192 ^ 1'b0 ;
  assign n4458 = ( n4192 & n4456 ) | ( n4192 & ~n4457 ) | ( n4456 & ~n4457 ) ;
  assign n4459 = n4331 ^ n4194 ^ x93 ;
  assign n4460 = n4360 ^ n4194 ^ 1'b0 ;
  assign n4461 = ( n4194 & n4459 ) | ( n4194 & ~n4460 ) | ( n4459 & ~n4460 ) ;
  assign n4462 = n4330 ^ n4196 ^ x92 ;
  assign n4463 = n4360 ^ n4196 ^ 1'b0 ;
  assign n4464 = ( n4196 & n4462 ) | ( n4196 & ~n4463 ) | ( n4462 & ~n4463 ) ;
  assign n4465 = n4328 ^ n4256 ^ x91 ;
  assign n4466 = n4360 ^ n4256 ^ 1'b0 ;
  assign n4467 = ( n4256 & n4465 ) | ( n4256 & ~n4466 ) | ( n4465 & ~n4466 ) ;
  assign n4468 = n4327 ^ n4198 ^ x90 ;
  assign n4469 = n4360 ^ n4198 ^ 1'b0 ;
  assign n4470 = ( n4198 & n4468 ) | ( n4198 & ~n4469 ) | ( n4468 & ~n4469 ) ;
  assign n4471 = n4326 ^ n4285 ^ x89 ;
  assign n4472 = n4360 ^ n4285 ^ 1'b0 ;
  assign n4473 = ( n4285 & n4471 ) | ( n4285 & ~n4472 ) | ( n4471 & ~n4472 ) ;
  assign n4474 = n4325 ^ n4239 ^ x88 ;
  assign n4475 = n4360 ^ n4239 ^ 1'b0 ;
  assign n4476 = ( n4239 & n4474 ) | ( n4239 & ~n4475 ) | ( n4474 & ~n4475 ) ;
  assign n4477 = x64 & n4360 ;
  assign n4478 = n4477 ^ x64 ^ x20 ;
  assign n4479 = ~x19 & x64 ;
  assign n4480 = n4479 ^ n4478 ^ x65 ;
  assign n4481 = ( x65 & n4479 ) | ( x65 & n4480 ) | ( n4479 & n4480 ) ;
  assign n4482 = n4481 ^ n4394 ^ x66 ;
  assign n4483 = ( x66 & n4481 ) | ( x66 & n4482 ) | ( n4481 & n4482 ) ;
  assign n4484 = ( x67 & ~n4392 ) | ( x67 & n4483 ) | ( ~n4392 & n4483 ) ;
  assign n4485 = ( x68 & ~n4437 ) | ( x68 & n4484 ) | ( ~n4437 & n4484 ) ;
  assign n4486 = ( x69 & ~n4390 ) | ( x69 & n4485 ) | ( ~n4390 & n4485 ) ;
  assign n4487 = ( x70 & ~n4434 ) | ( x70 & n4486 ) | ( ~n4434 & n4486 ) ;
  assign n4488 = ( x71 & ~n4388 ) | ( x71 & n4487 ) | ( ~n4388 & n4487 ) ;
  assign n4489 = ( x72 & ~n4386 ) | ( x72 & n4488 ) | ( ~n4386 & n4488 ) ;
  assign n4490 = ( x73 & ~n4384 ) | ( x73 & n4489 ) | ( ~n4384 & n4489 ) ;
  assign n4491 = ( x74 & ~n4382 ) | ( x74 & n4490 ) | ( ~n4382 & n4490 ) ;
  assign n4492 = ( x75 & ~n4380 ) | ( x75 & n4491 ) | ( ~n4380 & n4491 ) ;
  assign n4493 = n4484 ^ n4437 ^ x68 ;
  assign n4494 = ( x76 & ~n4378 ) | ( x76 & n4492 ) | ( ~n4378 & n4492 ) ;
  assign n4495 = ( x77 & ~n4376 ) | ( x77 & n4494 ) | ( ~n4376 & n4494 ) ;
  assign n4496 = n322 | n4395 ;
  assign n4497 = ( x78 & ~n4431 ) | ( x78 & n4495 ) | ( ~n4431 & n4495 ) ;
  assign n4498 = n4494 ^ n4376 ^ x77 ;
  assign n4499 = ( x79 & ~n4428 ) | ( x79 & n4497 ) | ( ~n4428 & n4497 ) ;
  assign n4500 = ( x80 & ~n4425 ) | ( x80 & n4499 ) | ( ~n4425 & n4499 ) ;
  assign n4501 = ( x81 & ~n4422 ) | ( x81 & n4500 ) | ( ~n4422 & n4500 ) ;
  assign n4502 = n4488 ^ n4386 ^ x72 ;
  assign n4503 = ( x82 & ~n4419 ) | ( x82 & n4501 ) | ( ~n4419 & n4501 ) ;
  assign n4504 = ( x83 & ~n4416 ) | ( x83 & n4503 ) | ( ~n4416 & n4503 ) ;
  assign n4505 = ( x84 & ~n4413 ) | ( x84 & n4504 ) | ( ~n4413 & n4504 ) ;
  assign n4506 = ( x108 & n176 ) | ( x108 & ~n4395 ) | ( n176 & ~n4395 ) ;
  assign n4507 = n3273 & n4496 ;
  assign n4508 = n4500 ^ n4422 ^ x81 ;
  assign n4509 = ( x85 & ~n4410 ) | ( x85 & n4505 ) | ( ~n4410 & n4505 ) ;
  assign n4510 = n4499 ^ n4425 ^ x80 ;
  assign n4511 = ( x86 & ~n4407 ) | ( x86 & n4509 ) | ( ~n4407 & n4509 ) ;
  assign n4512 = ( x87 & ~n4404 ) | ( x87 & n4511 ) | ( ~n4404 & n4511 ) ;
  assign n4513 = ( x88 & ~n4401 ) | ( x88 & n4512 ) | ( ~n4401 & n4512 ) ;
  assign n4514 = n4503 ^ n4416 ^ x83 ;
  assign n4515 = ( ~x108 & n176 ) | ( ~x108 & n4496 ) | ( n176 & n4496 ) ;
  assign n4516 = ( x89 & ~n4476 ) | ( x89 & n4513 ) | ( ~n4476 & n4513 ) ;
  assign n4517 = n4511 ^ n4404 ^ x87 ;
  assign n4518 = n4516 ^ n4473 ^ x90 ;
  assign n4519 = n4509 ^ n4407 ^ x86 ;
  assign n4520 = ( x90 & ~n4473 ) | ( x90 & n4516 ) | ( ~n4473 & n4516 ) ;
  assign n4521 = ( x91 & ~n4470 ) | ( x91 & n4520 ) | ( ~n4470 & n4520 ) ;
  assign n4522 = ( x92 & ~n4467 ) | ( x92 & n4521 ) | ( ~n4467 & n4521 ) ;
  assign n4523 = ( x93 & ~n4464 ) | ( x93 & n4522 ) | ( ~n4464 & n4522 ) ;
  assign n4524 = ( x94 & ~n4461 ) | ( x94 & n4523 ) | ( ~n4461 & n4523 ) ;
  assign n4525 = ( x95 & ~n4458 ) | ( x95 & n4524 ) | ( ~n4458 & n4524 ) ;
  assign n4526 = ( x96 & ~n4455 ) | ( x96 & n4525 ) | ( ~n4455 & n4525 ) ;
  assign n4527 = ( x97 & ~n4452 ) | ( x97 & n4526 ) | ( ~n4452 & n4526 ) ;
  assign n4528 = ( x98 & ~n4449 ) | ( x98 & n4527 ) | ( ~n4449 & n4527 ) ;
  assign n4529 = ( x99 & ~n4446 ) | ( x99 & n4528 ) | ( ~n4446 & n4528 ) ;
  assign n4530 = ( x100 & ~n4443 ) | ( x100 & n4529 ) | ( ~n4443 & n4529 ) ;
  assign n4531 = ( x101 & ~n4440 ) | ( x101 & n4530 ) | ( ~n4440 & n4530 ) ;
  assign n4532 = ( x102 & ~n4398 ) | ( x102 & n4531 ) | ( ~n4398 & n4531 ) ;
  assign n4533 = ( x103 & ~n4374 ) | ( x103 & n4532 ) | ( ~n4374 & n4532 ) ;
  assign n4534 = ( x104 & ~n4371 ) | ( x104 & n4533 ) | ( ~n4371 & n4533 ) ;
  assign n4535 = ( x105 & ~n4368 ) | ( x105 & n4534 ) | ( ~n4368 & n4534 ) ;
  assign n4536 = ( x106 & ~n4365 ) | ( x106 & n4535 ) | ( ~n4365 & n4535 ) ;
  assign n4537 = ( x107 & ~n4362 ) | ( x107 & n4536 ) | ( ~n4362 & n4536 ) ;
  assign n4538 = ( n4506 & n4515 ) | ( n4506 & ~n4537 ) | ( n4515 & ~n4537 ) ;
  assign n4539 = n4537 | n4538 ;
  assign n4540 = ( ~n4496 & n4507 ) | ( ~n4496 & n4539 ) | ( n4507 & n4539 ) ;
  assign n4541 = n4532 ^ n4374 ^ x103 ;
  assign n4542 = n4540 ^ n4374 ^ 1'b0 ;
  assign n4543 = ( n4374 & n4541 ) | ( n4374 & ~n4542 ) | ( n4541 & ~n4542 ) ;
  assign n4544 = n4530 ^ n4440 ^ x101 ;
  assign n4545 = n4540 ^ n4440 ^ 1'b0 ;
  assign n4546 = ( n4440 & n4544 ) | ( n4440 & ~n4545 ) | ( n4544 & ~n4545 ) ;
  assign n4547 = n4523 ^ n4461 ^ x94 ;
  assign n4548 = n4540 ^ n4461 ^ 1'b0 ;
  assign n4549 = ( n4461 & n4547 ) | ( n4461 & ~n4548 ) | ( n4547 & ~n4548 ) ;
  assign n4550 = n4522 ^ n4464 ^ x93 ;
  assign n4551 = n4540 ^ n4464 ^ 1'b0 ;
  assign n4552 = ( n4464 & n4550 ) | ( n4464 & ~n4551 ) | ( n4550 & ~n4551 ) ;
  assign n4553 = n4540 ^ n4473 ^ 1'b0 ;
  assign n4554 = ( n4473 & n4518 ) | ( n4473 & ~n4553 ) | ( n4518 & ~n4553 ) ;
  assign n4555 = n4540 ^ n4404 ^ 1'b0 ;
  assign n4556 = ( n4404 & n4517 ) | ( n4404 & ~n4555 ) | ( n4517 & ~n4555 ) ;
  assign n4557 = n4540 ^ n4407 ^ 1'b0 ;
  assign n4558 = ( n4407 & n4519 ) | ( n4407 & ~n4557 ) | ( n4519 & ~n4557 ) ;
  assign n4559 = n4540 ^ n4416 ^ 1'b0 ;
  assign n4560 = ( n4416 & n4514 ) | ( n4416 & ~n4559 ) | ( n4514 & ~n4559 ) ;
  assign n4561 = n4540 ^ n4422 ^ 1'b0 ;
  assign n4562 = ( n4422 & n4508 ) | ( n4422 & ~n4561 ) | ( n4508 & ~n4561 ) ;
  assign n4563 = n4540 ^ n4425 ^ 1'b0 ;
  assign n4564 = ( n4425 & n4510 ) | ( n4425 & ~n4563 ) | ( n4510 & ~n4563 ) ;
  assign n4565 = n4540 ^ n4376 ^ 1'b0 ;
  assign n4566 = ( n4376 & n4498 ) | ( n4376 & ~n4565 ) | ( n4498 & ~n4565 ) ;
  assign n4567 = n4540 ^ n4386 ^ 1'b0 ;
  assign n4568 = ( n4386 & n4502 ) | ( n4386 & ~n4567 ) | ( n4502 & ~n4567 ) ;
  assign n4569 = n4540 ^ n4437 ^ 1'b0 ;
  assign n4570 = ( n4437 & n4493 ) | ( n4437 & ~n4569 ) | ( n4493 & ~n4569 ) ;
  assign n4571 = n4540 ^ n4482 ^ 1'b0 ;
  assign n4572 = ( n4394 & n4482 ) | ( n4394 & n4571 ) | ( n4482 & n4571 ) ;
  assign n4573 = n4540 ^ n4480 ^ 1'b0 ;
  assign n4574 = ( n4478 & n4480 ) | ( n4478 & n4573 ) | ( n4480 & n4573 ) ;
  assign n4575 = n4507 & ~n4539 ;
  assign n4576 = ( n322 & n4507 ) | ( n322 & ~n4575 ) | ( n4507 & ~n4575 ) ;
  assign n4577 = n4536 ^ n4362 ^ x107 ;
  assign n4578 = n4540 ^ n4362 ^ 1'b0 ;
  assign n4579 = ( n4362 & n4577 ) | ( n4362 & ~n4578 ) | ( n4577 & ~n4578 ) ;
  assign n4580 = n4535 ^ n4365 ^ x106 ;
  assign n4581 = n4540 ^ n4365 ^ 1'b0 ;
  assign n4582 = ( n4365 & n4580 ) | ( n4365 & ~n4581 ) | ( n4580 & ~n4581 ) ;
  assign n4583 = n4505 ^ n4410 ^ x85 ;
  assign n4584 = n4540 ^ n4410 ^ 1'b0 ;
  assign n4585 = ( n4410 & n4583 ) | ( n4410 & ~n4584 ) | ( n4583 & ~n4584 ) ;
  assign n4586 = n4504 ^ n4413 ^ x84 ;
  assign n4587 = n4540 ^ n4413 ^ 1'b0 ;
  assign n4588 = ( n4413 & n4586 ) | ( n4413 & ~n4587 ) | ( n4586 & ~n4587 ) ;
  assign n4589 = n4501 ^ n4419 ^ x82 ;
  assign n4590 = n4540 ^ n4419 ^ 1'b0 ;
  assign n4591 = ( n4419 & n4589 ) | ( n4419 & ~n4590 ) | ( n4589 & ~n4590 ) ;
  assign n4592 = n4497 ^ n4428 ^ x79 ;
  assign n4593 = n4540 ^ n4428 ^ 1'b0 ;
  assign n4594 = ( n4428 & n4592 ) | ( n4428 & ~n4593 ) | ( n4592 & ~n4593 ) ;
  assign n4595 = n4495 ^ n4431 ^ x78 ;
  assign n4596 = n4540 ^ n4431 ^ 1'b0 ;
  assign n4597 = ( n4431 & n4595 ) | ( n4431 & ~n4596 ) | ( n4595 & ~n4596 ) ;
  assign n4598 = n4492 ^ n4378 ^ x76 ;
  assign n4599 = n4540 ^ n4378 ^ 1'b0 ;
  assign n4600 = ( n4378 & n4598 ) | ( n4378 & ~n4599 ) | ( n4598 & ~n4599 ) ;
  assign n4601 = n4491 ^ n4380 ^ x75 ;
  assign n4602 = n4540 ^ n4380 ^ 1'b0 ;
  assign n4603 = ( n4380 & n4601 ) | ( n4380 & ~n4602 ) | ( n4601 & ~n4602 ) ;
  assign n4604 = n4490 ^ n4382 ^ x74 ;
  assign n4605 = n4540 ^ n4382 ^ 1'b0 ;
  assign n4606 = ( n4382 & n4604 ) | ( n4382 & ~n4605 ) | ( n4604 & ~n4605 ) ;
  assign n4607 = n4489 ^ n4384 ^ x73 ;
  assign n4608 = n4540 ^ n4384 ^ 1'b0 ;
  assign n4609 = ( n4384 & n4607 ) | ( n4384 & ~n4608 ) | ( n4607 & ~n4608 ) ;
  assign n4610 = n4487 ^ n4388 ^ x71 ;
  assign n4611 = n4540 ^ n4388 ^ 1'b0 ;
  assign n4612 = ( n4388 & n4610 ) | ( n4388 & ~n4611 ) | ( n4610 & ~n4611 ) ;
  assign n4613 = n4486 ^ n4434 ^ x70 ;
  assign n4614 = n4540 ^ n4434 ^ 1'b0 ;
  assign n4615 = ( n4434 & n4613 ) | ( n4434 & ~n4614 ) | ( n4613 & ~n4614 ) ;
  assign n4616 = n4485 ^ n4390 ^ x69 ;
  assign n4617 = n4540 ^ n4390 ^ 1'b0 ;
  assign n4618 = ( n4390 & n4616 ) | ( n4390 & ~n4617 ) | ( n4616 & ~n4617 ) ;
  assign n4619 = n4483 ^ n4392 ^ x67 ;
  assign n4620 = n4540 ^ n4392 ^ 1'b0 ;
  assign n4621 = ( n4392 & n4619 ) | ( n4392 & ~n4620 ) | ( n4619 & ~n4620 ) ;
  assign n4622 = n4534 ^ n4368 ^ x105 ;
  assign n4623 = n4540 ^ n4368 ^ 1'b0 ;
  assign n4624 = ( n4368 & n4622 ) | ( n4368 & ~n4623 ) | ( n4622 & ~n4623 ) ;
  assign n4625 = n4533 ^ n4371 ^ x104 ;
  assign n4626 = n4540 ^ n4371 ^ 1'b0 ;
  assign n4627 = ( n4371 & n4625 ) | ( n4371 & ~n4626 ) | ( n4625 & ~n4626 ) ;
  assign n4628 = n4531 ^ n4398 ^ x102 ;
  assign n4629 = n4540 ^ n4398 ^ 1'b0 ;
  assign n4630 = ( n4398 & n4628 ) | ( n4398 & ~n4629 ) | ( n4628 & ~n4629 ) ;
  assign n4631 = n4529 ^ n4443 ^ x100 ;
  assign n4632 = n4540 ^ n4443 ^ 1'b0 ;
  assign n4633 = ( n4443 & n4631 ) | ( n4443 & ~n4632 ) | ( n4631 & ~n4632 ) ;
  assign n4634 = n4528 ^ n4446 ^ x99 ;
  assign n4635 = n4540 ^ n4446 ^ 1'b0 ;
  assign n4636 = ( n4446 & n4634 ) | ( n4446 & ~n4635 ) | ( n4634 & ~n4635 ) ;
  assign n4637 = n4527 ^ n4449 ^ x98 ;
  assign n4638 = n4540 ^ n4449 ^ 1'b0 ;
  assign n4639 = ( n4449 & n4637 ) | ( n4449 & ~n4638 ) | ( n4637 & ~n4638 ) ;
  assign n4640 = n4526 ^ n4452 ^ x97 ;
  assign n4641 = n4540 ^ n4452 ^ 1'b0 ;
  assign n4642 = ( n4452 & n4640 ) | ( n4452 & ~n4641 ) | ( n4640 & ~n4641 ) ;
  assign n4643 = n4525 ^ n4455 ^ x96 ;
  assign n4644 = n4540 ^ n4455 ^ 1'b0 ;
  assign n4645 = ( n4455 & n4643 ) | ( n4455 & ~n4644 ) | ( n4643 & ~n4644 ) ;
  assign n4646 = n4524 ^ n4458 ^ x95 ;
  assign n4647 = n4540 ^ n4458 ^ 1'b0 ;
  assign n4648 = ( n4458 & n4646 ) | ( n4458 & ~n4647 ) | ( n4646 & ~n4647 ) ;
  assign n4649 = n4521 ^ n4467 ^ x92 ;
  assign n4650 = n4540 ^ n4467 ^ 1'b0 ;
  assign n4651 = ( n4467 & n4649 ) | ( n4467 & ~n4650 ) | ( n4649 & ~n4650 ) ;
  assign n4652 = n4520 ^ n4470 ^ x91 ;
  assign n4653 = n4540 ^ n4470 ^ 1'b0 ;
  assign n4654 = ( n4470 & n4652 ) | ( n4470 & ~n4653 ) | ( n4652 & ~n4653 ) ;
  assign n4655 = n4513 ^ n4476 ^ x89 ;
  assign n4656 = n4540 ^ n4476 ^ 1'b0 ;
  assign n4657 = ( n4476 & n4655 ) | ( n4476 & ~n4656 ) | ( n4655 & ~n4656 ) ;
  assign n4658 = n4512 ^ n4401 ^ x88 ;
  assign n4659 = n4540 ^ n4401 ^ 1'b0 ;
  assign n4660 = ( n4401 & n4658 ) | ( n4401 & ~n4659 ) | ( n4658 & ~n4659 ) ;
  assign n4661 = x64 & n4540 ;
  assign n4662 = n4661 ^ x64 ^ x19 ;
  assign n4663 = ~x18 & x64 ;
  assign n4664 = n4663 ^ n4662 ^ x65 ;
  assign n4665 = ( x65 & n4663 ) | ( x65 & n4664 ) | ( n4663 & n4664 ) ;
  assign n4666 = n4665 ^ n4574 ^ x66 ;
  assign n4667 = ( x66 & n4665 ) | ( x66 & n4666 ) | ( n4665 & n4666 ) ;
  assign n4668 = ( x67 & ~n4572 ) | ( x67 & n4667 ) | ( ~n4572 & n4667 ) ;
  assign n4669 = ( x68 & ~n4621 ) | ( x68 & n4668 ) | ( ~n4621 & n4668 ) ;
  assign n4670 = ( x69 & ~n4570 ) | ( x69 & n4669 ) | ( ~n4570 & n4669 ) ;
  assign n4671 = ( ~x110 & x111 ) | ( ~x110 & n183 ) | ( x111 & n183 ) ;
  assign n4672 = ( x70 & ~n4618 ) | ( x70 & n4670 ) | ( ~n4618 & n4670 ) ;
  assign n4673 = ( x71 & ~n4615 ) | ( x71 & n4672 ) | ( ~n4615 & n4672 ) ;
  assign n4674 = ( x72 & ~n4612 ) | ( x72 & n4673 ) | ( ~n4612 & n4673 ) ;
  assign n4675 = ( x73 & ~n4568 ) | ( x73 & n4674 ) | ( ~n4568 & n4674 ) ;
  assign n4676 = n4669 ^ n4570 ^ x69 ;
  assign n4677 = n4667 ^ n4572 ^ x67 ;
  assign n4678 = n4668 ^ n4621 ^ x68 ;
  assign n4679 = n4670 ^ n4618 ^ x70 ;
  assign n4680 = n4673 ^ n4612 ^ x72 ;
  assign n4681 = n4674 ^ n4568 ^ x73 ;
  assign n4682 = n4675 ^ n4609 ^ x74 ;
  assign n4683 = n4672 ^ n4615 ^ x71 ;
  assign n4684 = ( x74 & ~n4609 ) | ( x74 & n4675 ) | ( ~n4609 & n4675 ) ;
  assign n4685 = ( x75 & ~n4606 ) | ( x75 & n4684 ) | ( ~n4606 & n4684 ) ;
  assign n4686 = ( x76 & ~n4603 ) | ( x76 & n4685 ) | ( ~n4603 & n4685 ) ;
  assign n4687 = n4685 ^ n4603 ^ x76 ;
  assign n4688 = ( x77 & ~n4600 ) | ( x77 & n4686 ) | ( ~n4600 & n4686 ) ;
  assign n4689 = ( x78 & ~n4566 ) | ( x78 & n4688 ) | ( ~n4566 & n4688 ) ;
  assign n4690 = ( x79 & ~n4597 ) | ( x79 & n4689 ) | ( ~n4597 & n4689 ) ;
  assign n4691 = ( x80 & ~n4594 ) | ( x80 & n4690 ) | ( ~n4594 & n4690 ) ;
  assign n4692 = ( x81 & ~n4564 ) | ( x81 & n4691 ) | ( ~n4564 & n4691 ) ;
  assign n4693 = n4684 ^ n4606 ^ x75 ;
  assign n4694 = ( x82 & ~n4562 ) | ( x82 & n4692 ) | ( ~n4562 & n4692 ) ;
  assign n4695 = ( x83 & ~n4591 ) | ( x83 & n4694 ) | ( ~n4591 & n4694 ) ;
  assign n4696 = ( x84 & ~n4560 ) | ( x84 & n4695 ) | ( ~n4560 & n4695 ) ;
  assign n4697 = ( x85 & ~n4588 ) | ( x85 & n4696 ) | ( ~n4588 & n4696 ) ;
  assign n4698 = ( x86 & ~n4585 ) | ( x86 & n4697 ) | ( ~n4585 & n4697 ) ;
  assign n4699 = n4686 ^ n4600 ^ x77 ;
  assign n4700 = n4688 ^ n4566 ^ x78 ;
  assign n4701 = n4689 ^ n4597 ^ x79 ;
  assign n4702 = n4690 ^ n4594 ^ x80 ;
  assign n4703 = n4691 ^ n4564 ^ x81 ;
  assign n4704 = n4692 ^ n4562 ^ x82 ;
  assign n4705 = n4694 ^ n4591 ^ x83 ;
  assign n4706 = n4695 ^ n4560 ^ x84 ;
  assign n4707 = n4696 ^ n4588 ^ x85 ;
  assign n4708 = n4697 ^ n4585 ^ x86 ;
  assign n4709 = ( x87 & ~n4558 ) | ( x87 & n4698 ) | ( ~n4558 & n4698 ) ;
  assign n4710 = ( x88 & ~n4556 ) | ( x88 & n4709 ) | ( ~n4556 & n4709 ) ;
  assign n4711 = ( x89 & ~n4660 ) | ( x89 & n4710 ) | ( ~n4660 & n4710 ) ;
  assign n4712 = x110 | n4671 ;
  assign n4713 = ( x90 & ~n4657 ) | ( x90 & n4711 ) | ( ~n4657 & n4711 ) ;
  assign n4714 = ( x91 & ~n4554 ) | ( x91 & n4713 ) | ( ~n4554 & n4713 ) ;
  assign n4715 = ( x92 & ~n4654 ) | ( x92 & n4714 ) | ( ~n4654 & n4714 ) ;
  assign n4716 = ( x93 & ~n4651 ) | ( x93 & n4715 ) | ( ~n4651 & n4715 ) ;
  assign n4717 = ( x94 & ~n4552 ) | ( x94 & n4716 ) | ( ~n4552 & n4716 ) ;
  assign n4718 = ( x95 & ~n4549 ) | ( x95 & n4717 ) | ( ~n4549 & n4717 ) ;
  assign n4719 = ( x96 & ~n4648 ) | ( x96 & n4718 ) | ( ~n4648 & n4718 ) ;
  assign n4720 = ( x97 & ~n4645 ) | ( x97 & n4719 ) | ( ~n4645 & n4719 ) ;
  assign n4721 = ( x98 & ~n4642 ) | ( x98 & n4720 ) | ( ~n4642 & n4720 ) ;
  assign n4722 = ( x99 & ~n4639 ) | ( x99 & n4721 ) | ( ~n4639 & n4721 ) ;
  assign n4723 = ( x100 & ~n4636 ) | ( x100 & n4722 ) | ( ~n4636 & n4722 ) ;
  assign n4724 = ( x101 & ~n4633 ) | ( x101 & n4723 ) | ( ~n4633 & n4723 ) ;
  assign n4725 = ( x102 & ~n4546 ) | ( x102 & n4724 ) | ( ~n4546 & n4724 ) ;
  assign n4726 = ( x103 & ~n4630 ) | ( x103 & n4725 ) | ( ~n4630 & n4725 ) ;
  assign n4727 = ( x104 & ~n4543 ) | ( x104 & n4726 ) | ( ~n4543 & n4726 ) ;
  assign n4728 = ( x105 & ~n4627 ) | ( x105 & n4727 ) | ( ~n4627 & n4727 ) ;
  assign n4729 = ( x106 & ~n4624 ) | ( x106 & n4728 ) | ( ~n4624 & n4728 ) ;
  assign n4730 = ( x107 & ~n4582 ) | ( x107 & n4729 ) | ( ~n4582 & n4729 ) ;
  assign n4731 = ( x108 & ~n4579 ) | ( x108 & n4730 ) | ( ~n4579 & n4730 ) ;
  assign n4732 = ( x109 & ~n4576 ) | ( x109 & n4731 ) | ( ~n4576 & n4731 ) ;
  assign n4733 = n4712 | n4732 ;
  assign n4734 = n4733 ^ n4708 ^ 1'b0 ;
  assign n4735 = ( n4585 & n4708 ) | ( n4585 & n4734 ) | ( n4708 & n4734 ) ;
  assign n4736 = n4733 ^ n4707 ^ 1'b0 ;
  assign n4737 = ( n4588 & n4707 ) | ( n4588 & n4736 ) | ( n4707 & n4736 ) ;
  assign n4738 = n4733 ^ n4706 ^ 1'b0 ;
  assign n4739 = ( n4560 & n4706 ) | ( n4560 & n4738 ) | ( n4706 & n4738 ) ;
  assign n4740 = n4733 ^ n4705 ^ 1'b0 ;
  assign n4741 = ( n4591 & n4705 ) | ( n4591 & n4740 ) | ( n4705 & n4740 ) ;
  assign n4742 = n4733 ^ n4704 ^ 1'b0 ;
  assign n4743 = ( n4562 & n4704 ) | ( n4562 & n4742 ) | ( n4704 & n4742 ) ;
  assign n4744 = n4733 ^ n4703 ^ 1'b0 ;
  assign n4745 = ( n4564 & n4703 ) | ( n4564 & n4744 ) | ( n4703 & n4744 ) ;
  assign n4746 = n4733 ^ n4702 ^ 1'b0 ;
  assign n4747 = ( n4594 & n4702 ) | ( n4594 & n4746 ) | ( n4702 & n4746 ) ;
  assign n4748 = n4733 ^ n4701 ^ 1'b0 ;
  assign n4749 = ( n4597 & n4701 ) | ( n4597 & n4748 ) | ( n4701 & n4748 ) ;
  assign n4750 = n4733 ^ n4700 ^ 1'b0 ;
  assign n4751 = ( n4566 & n4700 ) | ( n4566 & n4750 ) | ( n4700 & n4750 ) ;
  assign n4752 = n4733 ^ n4699 ^ 1'b0 ;
  assign n4753 = ( n4600 & n4699 ) | ( n4600 & n4752 ) | ( n4699 & n4752 ) ;
  assign n4754 = n4733 ^ n4687 ^ 1'b0 ;
  assign n4755 = ( n4603 & n4687 ) | ( n4603 & n4754 ) | ( n4687 & n4754 ) ;
  assign n4756 = n4733 ^ n4693 ^ 1'b0 ;
  assign n4757 = ( n4606 & n4693 ) | ( n4606 & n4756 ) | ( n4693 & n4756 ) ;
  assign n4758 = n4733 ^ n4682 ^ 1'b0 ;
  assign n4759 = ( n4609 & n4682 ) | ( n4609 & n4758 ) | ( n4682 & n4758 ) ;
  assign n4760 = n4733 ^ n4681 ^ 1'b0 ;
  assign n4761 = ( n4568 & n4681 ) | ( n4568 & n4760 ) | ( n4681 & n4760 ) ;
  assign n4762 = n4733 ^ n4680 ^ 1'b0 ;
  assign n4763 = ( n4612 & n4680 ) | ( n4612 & n4762 ) | ( n4680 & n4762 ) ;
  assign n4764 = n4733 ^ n4683 ^ 1'b0 ;
  assign n4765 = ( n4615 & n4683 ) | ( n4615 & n4764 ) | ( n4683 & n4764 ) ;
  assign n4766 = n4733 ^ n4679 ^ 1'b0 ;
  assign n4767 = ( n4618 & n4679 ) | ( n4618 & n4766 ) | ( n4679 & n4766 ) ;
  assign n4768 = n4733 ^ n4676 ^ 1'b0 ;
  assign n4769 = ( n4570 & n4676 ) | ( n4570 & n4768 ) | ( n4676 & n4768 ) ;
  assign n4770 = n4733 ^ n4678 ^ 1'b0 ;
  assign n4771 = ( n4621 & n4678 ) | ( n4621 & n4770 ) | ( n4678 & n4770 ) ;
  assign n4772 = n4733 ^ n4677 ^ 1'b0 ;
  assign n4773 = ( n4572 & n4677 ) | ( n4572 & n4772 ) | ( n4677 & n4772 ) ;
  assign n4774 = n4733 ^ n4662 ^ 1'b0 ;
  assign n4775 = ( n4662 & n4664 ) | ( n4662 & ~n4774 ) | ( n4664 & ~n4774 ) ;
  assign n4776 = n4731 ^ n4576 ^ x109 ;
  assign n4777 = n4724 ^ n4546 ^ x102 ;
  assign n4778 = n4777 ^ n4733 ^ 1'b0 ;
  assign n4779 = n4714 ^ n4654 ^ x92 ;
  assign n4780 = n4722 ^ n4636 ^ x100 ;
  assign n4781 = ( n4546 & n4777 ) | ( n4546 & n4778 ) | ( n4777 & n4778 ) ;
  assign n4782 = n4723 ^ n4633 ^ x101 ;
  assign n4783 = n4782 ^ n4733 ^ 1'b0 ;
  assign n4784 = ( n4633 & n4782 ) | ( n4633 & n4783 ) | ( n4782 & n4783 ) ;
  assign n4785 = n4698 ^ n4558 ^ x87 ;
  assign n4786 = n4720 ^ n4642 ^ x98 ;
  assign n4787 = n4711 ^ n4657 ^ x90 ;
  assign n4788 = n4787 ^ n4733 ^ 1'b0 ;
  assign n4789 = n4718 ^ n4648 ^ x96 ;
  assign n4790 = n4789 ^ n4733 ^ 1'b0 ;
  assign n4791 = n4710 ^ n4660 ^ x89 ;
  assign n4792 = n4717 ^ n4549 ^ x95 ;
  assign n4793 = n4719 ^ n4645 ^ x97 ;
  assign n4794 = n4793 ^ n4733 ^ 1'b0 ;
  assign n4795 = ( n4648 & n4789 ) | ( n4648 & n4790 ) | ( n4789 & n4790 ) ;
  assign n4796 = n4715 ^ n4651 ^ x93 ;
  assign n4797 = n4796 ^ n4733 ^ 1'b0 ;
  assign n4798 = n4721 ^ n4639 ^ x99 ;
  assign n4799 = n4716 ^ n4552 ^ x94 ;
  assign n4800 = n4779 ^ n4733 ^ 1'b0 ;
  assign n4801 = ( n4654 & n4779 ) | ( n4654 & n4800 ) | ( n4779 & n4800 ) ;
  assign n4802 = n4725 ^ n4630 ^ x103 ;
  assign n4803 = n4802 ^ n4733 ^ 1'b0 ;
  assign n4804 = n4713 ^ n4554 ^ x91 ;
  assign n4805 = n4792 ^ n4733 ^ 1'b0 ;
  assign n4806 = ( n4645 & n4793 ) | ( n4645 & n4794 ) | ( n4793 & n4794 ) ;
  assign n4807 = n4798 ^ n4733 ^ 1'b0 ;
  assign n4808 = n4780 ^ n4733 ^ 1'b0 ;
  assign n4809 = ( n4630 & n4802 ) | ( n4630 & n4803 ) | ( n4802 & n4803 ) ;
  assign n4810 = n4799 ^ n4733 ^ 1'b0 ;
  assign n4811 = ~n4733 & n4776 ;
  assign n4812 = n4804 ^ n4733 ^ 1'b0 ;
  assign n4813 = ( n4651 & n4796 ) | ( n4651 & n4797 ) | ( n4796 & n4797 ) ;
  assign n4814 = n4791 ^ n4733 ^ 1'b0 ;
  assign n4815 = n4785 ^ n4733 ^ 1'b0 ;
  assign n4816 = ( n4636 & n4780 ) | ( n4636 & n4808 ) | ( n4780 & n4808 ) ;
  assign n4817 = n4786 ^ n4733 ^ 1'b0 ;
  assign n4818 = ( n4639 & n4798 ) | ( n4639 & n4807 ) | ( n4798 & n4807 ) ;
  assign n4819 = n4709 ^ n4556 ^ x88 ;
  assign n4820 = ( n4660 & n4791 ) | ( n4660 & n4814 ) | ( n4791 & n4814 ) ;
  assign n4821 = ( n4549 & n4792 ) | ( n4549 & n4805 ) | ( n4792 & n4805 ) ;
  assign n4822 = ( n4554 & n4804 ) | ( n4554 & n4812 ) | ( n4804 & n4812 ) ;
  assign n4823 = ( n4552 & n4799 ) | ( n4552 & n4810 ) | ( n4799 & n4810 ) ;
  assign n4824 = ( n4642 & n4786 ) | ( n4642 & n4817 ) | ( n4786 & n4817 ) ;
  assign n4825 = n4819 ^ n4733 ^ 1'b0 ;
  assign n4826 = ( n4558 & n4785 ) | ( n4558 & n4815 ) | ( n4785 & n4815 ) ;
  assign n4827 = ( n4657 & n4787 ) | ( n4657 & n4788 ) | ( n4787 & n4788 ) ;
  assign n4828 = ( n4556 & n4819 ) | ( n4556 & n4825 ) | ( n4819 & n4825 ) ;
  assign n4829 = n4726 ^ n4543 ^ x104 ;
  assign n4830 = n4733 ^ n4574 ^ 1'b0 ;
  assign n4831 = x18 & x64 ;
  assign n4832 = x110 | n4732 ;
  assign n4833 = ~x17 & x64 ;
  assign n4834 = ( n1298 & n4831 ) | ( n1298 & ~n4832 ) | ( n4831 & ~n4832 ) ;
  assign n4835 = ~n1298 & n4834 ;
  assign n4836 = n4663 & ~n4733 ;
  assign n4837 = n4730 ^ n4579 ^ x108 ;
  assign n4838 = n4576 & n4733 ;
  assign n4839 = ( x18 & ~n4835 ) | ( x18 & n4836 ) | ( ~n4835 & n4836 ) ;
  assign n4840 = ( n4574 & n4666 ) | ( n4574 & ~n4830 ) | ( n4666 & ~n4830 ) ;
  assign n4841 = n4839 ^ n4833 ^ x65 ;
  assign n4842 = n4727 ^ n4627 ^ x105 ;
  assign n4843 = n4728 ^ n4624 ^ x106 ;
  assign n4844 = n322 | n4838 ;
  assign n4845 = n4842 ^ n4733 ^ 1'b0 ;
  assign n4846 = n4843 ^ n4733 ^ 1'b0 ;
  assign n4847 = ( x65 & n4833 ) | ( x65 & n4841 ) | ( n4833 & n4841 ) ;
  assign n4848 = ( n4624 & n4843 ) | ( n4624 & n4846 ) | ( n4843 & n4846 ) ;
  assign n4849 = n4712 & n4844 ;
  assign n4850 = ( n4627 & n4842 ) | ( n4627 & n4845 ) | ( n4842 & n4845 ) ;
  assign n4851 = n4829 ^ n4733 ^ 1'b0 ;
  assign n4852 = n4837 ^ n4733 ^ 1'b0 ;
  assign n4853 = ( n4543 & n4829 ) | ( n4543 & n4851 ) | ( n4829 & n4851 ) ;
  assign n4854 = n4847 ^ n4775 ^ x66 ;
  assign n4855 = ( x66 & n4847 ) | ( x66 & n4854 ) | ( n4847 & n4854 ) ;
  assign n4856 = ( x67 & ~n4840 ) | ( x67 & n4855 ) | ( ~n4840 & n4855 ) ;
  assign n4857 = n4856 ^ n4773 ^ x68 ;
  assign n4858 = ( n4579 & n4837 ) | ( n4579 & n4852 ) | ( n4837 & n4852 ) ;
  assign n4859 = ( n1298 & ~n4811 ) | ( n1298 & n4838 ) | ( ~n4811 & n4838 ) ;
  assign n4860 = n4729 ^ n4582 ^ x107 ;
  assign n4861 = n4860 ^ n4733 ^ 1'b0 ;
  assign n4862 = ( n4582 & n4860 ) | ( n4582 & n4861 ) | ( n4860 & n4861 ) ;
  assign n4863 = ( ~x110 & n1298 ) | ( ~x110 & n4844 ) | ( n1298 & n4844 ) ;
  assign n4864 = n4811 | n4838 ;
  assign n4865 = n4859 ^ n4811 ^ x110 ;
  assign n4866 = ( x68 & ~n4773 ) | ( x68 & n4856 ) | ( ~n4773 & n4856 ) ;
  assign n4867 = ( x69 & ~n4771 ) | ( x69 & n4866 ) | ( ~n4771 & n4866 ) ;
  assign n4868 = n4576 & n4712 ;
  assign n4869 = n4855 ^ n4840 ^ x67 ;
  assign n4870 = ( x110 & n1298 ) | ( x110 & ~n4838 ) | ( n1298 & ~n4838 ) ;
  assign n4871 = n4866 ^ n4771 ^ x69 ;
  assign n4872 = ~n4712 & n4864 ;
  assign n4873 = ( x70 & ~n4769 ) | ( x70 & n4867 ) | ( ~n4769 & n4867 ) ;
  assign n4874 = ( x71 & ~n4767 ) | ( x71 & n4873 ) | ( ~n4767 & n4873 ) ;
  assign n4875 = ( x72 & ~n4765 ) | ( x72 & n4874 ) | ( ~n4765 & n4874 ) ;
  assign n4876 = ( x73 & ~n4763 ) | ( x73 & n4875 ) | ( ~n4763 & n4875 ) ;
  assign n4877 = ( x74 & ~n4761 ) | ( x74 & n4876 ) | ( ~n4761 & n4876 ) ;
  assign n4878 = ( x75 & ~n4759 ) | ( x75 & n4877 ) | ( ~n4759 & n4877 ) ;
  assign n4879 = ( x76 & ~n4757 ) | ( x76 & n4878 ) | ( ~n4757 & n4878 ) ;
  assign n4880 = ( x77 & ~n4755 ) | ( x77 & n4879 ) | ( ~n4755 & n4879 ) ;
  assign n4881 = ( x78 & ~n4753 ) | ( x78 & n4880 ) | ( ~n4753 & n4880 ) ;
  assign n4882 = ( x79 & ~n4751 ) | ( x79 & n4881 ) | ( ~n4751 & n4881 ) ;
  assign n4883 = ( x80 & ~n4749 ) | ( x80 & n4882 ) | ( ~n4749 & n4882 ) ;
  assign n4884 = ( x81 & ~n4747 ) | ( x81 & n4883 ) | ( ~n4747 & n4883 ) ;
  assign n4885 = ( x82 & ~n4745 ) | ( x82 & n4884 ) | ( ~n4745 & n4884 ) ;
  assign n4886 = ( x83 & ~n4743 ) | ( x83 & n4885 ) | ( ~n4743 & n4885 ) ;
  assign n4887 = ( x84 & ~n4741 ) | ( x84 & n4886 ) | ( ~n4741 & n4886 ) ;
  assign n4888 = ( x85 & ~n4739 ) | ( x85 & n4887 ) | ( ~n4739 & n4887 ) ;
  assign n4889 = ( x86 & ~n4737 ) | ( x86 & n4888 ) | ( ~n4737 & n4888 ) ;
  assign n4890 = ( x87 & ~n4735 ) | ( x87 & n4889 ) | ( ~n4735 & n4889 ) ;
  assign n4891 = ( x88 & ~n4826 ) | ( x88 & n4890 ) | ( ~n4826 & n4890 ) ;
  assign n4892 = ( x89 & ~n4828 ) | ( x89 & n4891 ) | ( ~n4828 & n4891 ) ;
  assign n4893 = ( x90 & ~n4820 ) | ( x90 & n4892 ) | ( ~n4820 & n4892 ) ;
  assign n4894 = ( x91 & ~n4827 ) | ( x91 & n4893 ) | ( ~n4827 & n4893 ) ;
  assign n4895 = ( x92 & ~n4822 ) | ( x92 & n4894 ) | ( ~n4822 & n4894 ) ;
  assign n4896 = ( x93 & ~n4801 ) | ( x93 & n4895 ) | ( ~n4801 & n4895 ) ;
  assign n4897 = ( x94 & ~n4813 ) | ( x94 & n4896 ) | ( ~n4813 & n4896 ) ;
  assign n4898 = ( x95 & ~n4823 ) | ( x95 & n4897 ) | ( ~n4823 & n4897 ) ;
  assign n4899 = ( x96 & ~n4821 ) | ( x96 & n4898 ) | ( ~n4821 & n4898 ) ;
  assign n4900 = ( x97 & ~n4795 ) | ( x97 & n4899 ) | ( ~n4795 & n4899 ) ;
  assign n4901 = ( x98 & ~n4806 ) | ( x98 & n4900 ) | ( ~n4806 & n4900 ) ;
  assign n4902 = ( x99 & ~n4824 ) | ( x99 & n4901 ) | ( ~n4824 & n4901 ) ;
  assign n4903 = n4874 ^ n4765 ^ x72 ;
  assign n4904 = n4875 ^ n4763 ^ x73 ;
  assign n4905 = n4895 ^ n4801 ^ x93 ;
  assign n4906 = n4876 ^ n4761 ^ x74 ;
  assign n4907 = n4891 ^ n4828 ^ x89 ;
  assign n4908 = n4878 ^ n4757 ^ x76 ;
  assign n4909 = n4879 ^ n4755 ^ x77 ;
  assign n4910 = n4880 ^ n4753 ^ x78 ;
  assign n4911 = n4881 ^ n4751 ^ x79 ;
  assign n4912 = n4882 ^ n4749 ^ x80 ;
  assign n4913 = n4883 ^ n4747 ^ x81 ;
  assign n4914 = n4884 ^ n4745 ^ x82 ;
  assign n4915 = n4885 ^ n4743 ^ x83 ;
  assign n4916 = n4890 ^ n4826 ^ x88 ;
  assign n4917 = n4887 ^ n4739 ^ x85 ;
  assign n4918 = n4888 ^ n4737 ^ x86 ;
  assign n4919 = n4889 ^ n4735 ^ x87 ;
  assign n4920 = ( x100 & ~n4818 ) | ( x100 & n4902 ) | ( ~n4818 & n4902 ) ;
  assign n4921 = ( x101 & ~n4816 ) | ( x101 & n4920 ) | ( ~n4816 & n4920 ) ;
  assign n4922 = n4892 ^ n4820 ^ x90 ;
  assign n4923 = n4893 ^ n4827 ^ x91 ;
  assign n4924 = n4894 ^ n4822 ^ x92 ;
  assign n4925 = n4920 ^ n4816 ^ x101 ;
  assign n4926 = n4896 ^ n4813 ^ x94 ;
  assign n4927 = n4897 ^ n4823 ^ x95 ;
  assign n4928 = n4898 ^ n4821 ^ x96 ;
  assign n4929 = n4899 ^ n4795 ^ x97 ;
  assign n4930 = n4900 ^ n4806 ^ x98 ;
  assign n4931 = n4901 ^ n4824 ^ x99 ;
  assign n4932 = n4902 ^ n4818 ^ x100 ;
  assign n4933 = ( x102 & ~n4784 ) | ( x102 & n4921 ) | ( ~n4784 & n4921 ) ;
  assign n4934 = n4933 ^ n4781 ^ x103 ;
  assign n4935 = n4921 ^ n4784 ^ x102 ;
  assign n4936 = n4867 ^ n4769 ^ x70 ;
  assign n4937 = ( x103 & ~n4781 ) | ( x103 & n4933 ) | ( ~n4781 & n4933 ) ;
  assign n4938 = ( x104 & ~n4809 ) | ( x104 & n4937 ) | ( ~n4809 & n4937 ) ;
  assign n4939 = ( x105 & ~n4853 ) | ( x105 & n4938 ) | ( ~n4853 & n4938 ) ;
  assign n4940 = ( x106 & ~n4850 ) | ( x106 & n4939 ) | ( ~n4850 & n4939 ) ;
  assign n4941 = ( x107 & ~n4848 ) | ( x107 & n4940 ) | ( ~n4848 & n4940 ) ;
  assign n4942 = ( x108 & ~n4862 ) | ( x108 & n4941 ) | ( ~n4862 & n4941 ) ;
  assign n4943 = ( x109 & ~n4858 ) | ( x109 & n4942 ) | ( ~n4858 & n4942 ) ;
  assign n4944 = ( n4863 & n4870 ) | ( n4863 & ~n4943 ) | ( n4870 & ~n4943 ) ;
  assign n4945 = ( ~n1298 & n4865 ) | ( ~n1298 & n4943 ) | ( n4865 & n4943 ) ;
  assign n4946 = n1298 | n4945 ;
  assign n4947 = n4943 | n4944 ;
  assign n4948 = ( ~n4844 & n4849 ) | ( ~n4844 & n4947 ) | ( n4849 & n4947 ) ;
  assign n4949 = n4948 ^ n4914 ^ 1'b0 ;
  assign n4950 = ~n4872 & n4946 ;
  assign n4951 = n4950 ^ n4745 ^ 1'b0 ;
  assign n4952 = ( n4745 & n4914 ) | ( n4745 & ~n4951 ) | ( n4914 & ~n4951 ) ;
  assign n4953 = n4942 ^ n4858 ^ x109 ;
  assign n4954 = ( n4745 & n4914 ) | ( n4745 & n4949 ) | ( n4914 & n4949 ) ;
  assign n4955 = n4950 ^ n4769 ^ 1'b0 ;
  assign n4956 = n4868 & n4947 ;
  assign n4957 = n4943 ^ n4864 ^ x110 ;
  assign n4958 = n4868 & ~n4946 ;
  assign n4959 = ( n4769 & n4936 ) | ( n4769 & ~n4955 ) | ( n4936 & ~n4955 ) ;
  assign n4960 = n4948 ^ n4869 ^ 1'b0 ;
  assign n4961 = n4950 ^ n4840 ^ 1'b0 ;
  assign n4962 = ( n4840 & n4869 ) | ( n4840 & n4960 ) | ( n4869 & n4960 ) ;
  assign n4963 = ( n4840 & n4869 ) | ( n4840 & ~n4961 ) | ( n4869 & ~n4961 ) ;
  assign n4964 = ~n4950 & n4957 ;
  assign n4965 = n4948 ^ n4931 ^ 1'b0 ;
  assign n4966 = ( n4868 & ~n4958 ) | ( n4868 & n4964 ) | ( ~n4958 & n4964 ) ;
  assign n4967 = n4939 ^ n4850 ^ x106 ;
  assign n4968 = n4948 ^ n4906 ^ 1'b0 ;
  assign n4969 = n4948 ^ n4936 ^ 1'b0 ;
  assign n4970 = n4948 ^ n4924 ^ 1'b0 ;
  assign n4971 = ( n4769 & n4936 ) | ( n4769 & n4969 ) | ( n4936 & n4969 ) ;
  assign n4972 = ( n4761 & n4906 ) | ( n4761 & n4968 ) | ( n4906 & n4968 ) ;
  assign n4973 = n4950 ^ n4749 ^ 1'b0 ;
  assign n4974 = ( n4749 & n4912 ) | ( n4749 & ~n4973 ) | ( n4912 & ~n4973 ) ;
  assign n4975 = n4950 ^ n4761 ^ 1'b0 ;
  assign n4976 = ( n4822 & n4924 ) | ( n4822 & n4970 ) | ( n4924 & n4970 ) ;
  assign n4977 = ( n4761 & n4906 ) | ( n4761 & ~n4975 ) | ( n4906 & ~n4975 ) ;
  assign n4978 = n4948 ^ n4909 ^ 1'b0 ;
  assign n4979 = n4950 ^ n4755 ^ 1'b0 ;
  assign n4980 = ( n4755 & n4909 ) | ( n4755 & ~n4979 ) | ( n4909 & ~n4979 ) ;
  assign n4981 = ( n4755 & n4909 ) | ( n4755 & n4978 ) | ( n4909 & n4978 ) ;
  assign n4982 = n4950 ^ n4824 ^ 1'b0 ;
  assign n4983 = n4941 ^ n4862 ^ x108 ;
  assign n4984 = ( n4824 & n4931 ) | ( n4824 & ~n4982 ) | ( n4931 & ~n4982 ) ;
  assign n4985 = n4948 ^ n4927 ^ 1'b0 ;
  assign n4986 = ( n4824 & n4931 ) | ( n4824 & n4965 ) | ( n4931 & n4965 ) ;
  assign n4987 = n4950 ^ n4822 ^ 1'b0 ;
  assign n4988 = ( n4822 & n4924 ) | ( n4822 & ~n4987 ) | ( n4924 & ~n4987 ) ;
  assign n4989 = n4950 ^ n4823 ^ 1'b0 ;
  assign n4990 = ( n4823 & n4927 ) | ( n4823 & ~n4989 ) | ( n4927 & ~n4989 ) ;
  assign n4991 = ( n4823 & n4927 ) | ( n4823 & n4985 ) | ( n4927 & n4985 ) ;
  assign n4992 = n4950 ^ n4737 ^ 1'b0 ;
  assign n4993 = ( n4737 & n4918 ) | ( n4737 & ~n4992 ) | ( n4918 & ~n4992 ) ;
  assign n4994 = n4948 ^ n4926 ^ 1'b0 ;
  assign n4995 = n4948 ^ n4922 ^ 1'b0 ;
  assign n4996 = ( n4820 & n4922 ) | ( n4820 & n4995 ) | ( n4922 & n4995 ) ;
  assign n4997 = n4950 ^ n4820 ^ 1'b0 ;
  assign n4998 = ( n4820 & n4922 ) | ( n4820 & ~n4997 ) | ( n4922 & ~n4997 ) ;
  assign n4999 = n4950 ^ n4813 ^ 1'b0 ;
  assign n5000 = ( n4813 & n4926 ) | ( n4813 & n4994 ) | ( n4926 & n4994 ) ;
  assign n5001 = n4948 ^ n4903 ^ 1'b0 ;
  assign n5002 = n4940 ^ n4848 ^ x107 ;
  assign n5003 = ( n4765 & n4903 ) | ( n4765 & n5001 ) | ( n4903 & n5001 ) ;
  assign n5004 = ( n4813 & n4926 ) | ( n4813 & ~n4999 ) | ( n4926 & ~n4999 ) ;
  assign n5005 = n4948 ^ n4918 ^ 1'b0 ;
  assign n5006 = n4950 ^ n4806 ^ 1'b0 ;
  assign n5007 = ( n4806 & n4930 ) | ( n4806 & ~n5006 ) | ( n4930 & ~n5006 ) ;
  assign n5008 = ( n4737 & n4918 ) | ( n4737 & n5005 ) | ( n4918 & n5005 ) ;
  assign n5009 = n4950 ^ n4765 ^ 1'b0 ;
  assign n5010 = n4948 ^ n4930 ^ 1'b0 ;
  assign n5011 = ( n4806 & n4930 ) | ( n4806 & n5010 ) | ( n4930 & n5010 ) ;
  assign n5012 = n4948 ^ n4912 ^ 1'b0 ;
  assign n5013 = ( n4749 & n4912 ) | ( n4749 & n5012 ) | ( n4912 & n5012 ) ;
  assign n5014 = ( n4765 & n4903 ) | ( n4765 & ~n5009 ) | ( n4903 & ~n5009 ) ;
  assign n5015 = n4948 ^ n4923 ^ 1'b0 ;
  assign n5016 = ( n4827 & n4923 ) | ( n4827 & n5015 ) | ( n4923 & n5015 ) ;
  assign n5017 = n4937 ^ n4809 ^ x104 ;
  assign n5018 = n4950 ^ n4827 ^ 1'b0 ;
  assign n5019 = ( n4827 & n4923 ) | ( n4827 & ~n5018 ) | ( n4923 & ~n5018 ) ;
  assign n5020 = n4948 ^ n4841 ^ 1'b0 ;
  assign n5021 = ( n4839 & n4841 ) | ( n4839 & n5020 ) | ( n4841 & n5020 ) ;
  assign n5022 = n4950 ^ n4841 ^ 1'b0 ;
  assign n5023 = ( n4839 & n4841 ) | ( n4839 & n5022 ) | ( n4841 & n5022 ) ;
  assign n5024 = n4950 ^ n4771 ^ 1'b0 ;
  assign n5025 = ( n4771 & n4871 ) | ( n4771 & ~n5024 ) | ( n4871 & ~n5024 ) ;
  assign n5026 = n4948 ^ n4871 ^ 1'b0 ;
  assign n5027 = ( n4771 & n4871 ) | ( n4771 & n5026 ) | ( n4871 & n5026 ) ;
  assign n5028 = n4948 ^ n4854 ^ 1'b0 ;
  assign n5029 = ( n4775 & n4854 ) | ( n4775 & n5028 ) | ( n4854 & n5028 ) ;
  assign n5030 = n4886 ^ n4741 ^ x84 ;
  assign n5031 = n4950 ^ n4854 ^ 1'b0 ;
  assign n5032 = ( n4775 & n4854 ) | ( n4775 & n5031 ) | ( n4854 & n5031 ) ;
  assign n5033 = n4948 ^ n4911 ^ 1'b0 ;
  assign n5034 = ( n4751 & n4911 ) | ( n4751 & n5033 ) | ( n4911 & n5033 ) ;
  assign n5035 = n4950 ^ n4751 ^ 1'b0 ;
  assign n5036 = ( n4751 & n4911 ) | ( n4751 & ~n5035 ) | ( n4911 & ~n5035 ) ;
  assign n5037 = n4950 ^ n4862 ^ 1'b0 ;
  assign n5038 = ( n4862 & n4983 ) | ( n4862 & ~n5037 ) | ( n4983 & ~n5037 ) ;
  assign n5039 = n4983 ^ n4948 ^ 1'b0 ;
  assign n5040 = ( n4862 & n4983 ) | ( n4862 & n5039 ) | ( n4983 & n5039 ) ;
  assign n5041 = n4950 ^ n4809 ^ 1'b0 ;
  assign n5042 = ( n4809 & n5017 ) | ( n4809 & ~n5041 ) | ( n5017 & ~n5041 ) ;
  assign n5043 = n5017 ^ n4948 ^ 1'b0 ;
  assign n5044 = ( n4809 & n5017 ) | ( n4809 & n5043 ) | ( n5017 & n5043 ) ;
  assign n5045 = n4950 ^ n4741 ^ 1'b0 ;
  assign n5046 = n5030 ^ n4948 ^ 1'b0 ;
  assign n5047 = ( n4741 & n5030 ) | ( n4741 & n5046 ) | ( n5030 & n5046 ) ;
  assign n5048 = ( n4741 & n5030 ) | ( n4741 & ~n5045 ) | ( n5030 & ~n5045 ) ;
  assign n5049 = n4950 ^ n4753 ^ 1'b0 ;
  assign n5050 = n4877 ^ n4759 ^ x75 ;
  assign n5051 = ( n4753 & n4910 ) | ( n4753 & ~n5049 ) | ( n4910 & ~n5049 ) ;
  assign n5052 = n4948 ^ n4910 ^ 1'b0 ;
  assign n5053 = ( n4753 & n4910 ) | ( n4753 & n5052 ) | ( n4910 & n5052 ) ;
  assign n5054 = n4950 ^ n4739 ^ 1'b0 ;
  assign n5055 = n4948 ^ n4917 ^ 1'b0 ;
  assign n5056 = ( n4739 & n4917 ) | ( n4739 & ~n5054 ) | ( n4917 & ~n5054 ) ;
  assign n5057 = ( n4739 & n4917 ) | ( n4739 & n5055 ) | ( n4917 & n5055 ) ;
  assign n5058 = n4948 ^ n4913 ^ 1'b0 ;
  assign n5059 = n4950 ^ n4747 ^ 1'b0 ;
  assign n5060 = ( n4747 & n4913 ) | ( n4747 & ~n5059 ) | ( n4913 & ~n5059 ) ;
  assign n5061 = ( n4747 & n4913 ) | ( n4747 & n5058 ) | ( n4913 & n5058 ) ;
  assign n5062 = n4948 ^ n4905 ^ 1'b0 ;
  assign n5063 = ( n4801 & n4905 ) | ( n4801 & n5062 ) | ( n4905 & n5062 ) ;
  assign n5064 = n4950 ^ n4801 ^ 1'b0 ;
  assign n5065 = ( n4801 & n4905 ) | ( n4801 & ~n5064 ) | ( n4905 & ~n5064 ) ;
  assign n5066 = n4953 ^ n4948 ^ 1'b0 ;
  assign n5067 = ( n4858 & n4953 ) | ( n4858 & n5066 ) | ( n4953 & n5066 ) ;
  assign n5068 = n4950 ^ n4858 ^ 1'b0 ;
  assign n5069 = ( n4858 & n4953 ) | ( n4858 & ~n5068 ) | ( n4953 & ~n5068 ) ;
  assign n5070 = n4950 ^ n4821 ^ 1'b0 ;
  assign n5071 = n4948 ^ n4928 ^ 1'b0 ;
  assign n5072 = ( n4821 & n4928 ) | ( n4821 & ~n5070 ) | ( n4928 & ~n5070 ) ;
  assign n5073 = ( n4821 & n4928 ) | ( n4821 & n5071 ) | ( n4928 & n5071 ) ;
  assign n5074 = n4948 ^ n4916 ^ 1'b0 ;
  assign n5075 = n4950 ^ n4826 ^ 1'b0 ;
  assign n5076 = ( n4826 & n4916 ) | ( n4826 & ~n5075 ) | ( n4916 & ~n5075 ) ;
  assign n5077 = ( n4826 & n4916 ) | ( n4826 & n5074 ) | ( n4916 & n5074 ) ;
  assign n5078 = n4873 ^ n4767 ^ x71 ;
  assign n5079 = n4950 ^ n4828 ^ 1'b0 ;
  assign n5080 = ( n4828 & n4907 ) | ( n4828 & ~n5079 ) | ( n4907 & ~n5079 ) ;
  assign n5081 = n4948 ^ n4907 ^ 1'b0 ;
  assign n5082 = ( n4828 & n4907 ) | ( n4828 & n5081 ) | ( n4907 & n5081 ) ;
  assign n5083 = n4950 ^ n4735 ^ 1'b0 ;
  assign n5084 = n4948 ^ n4919 ^ 1'b0 ;
  assign n5085 = ( n4735 & n4919 ) | ( n4735 & n5084 ) | ( n4919 & n5084 ) ;
  assign n5086 = ( n4735 & n4919 ) | ( n4735 & ~n5083 ) | ( n4919 & ~n5083 ) ;
  assign n5087 = n4948 ^ n4932 ^ 1'b0 ;
  assign n5088 = n4950 ^ n4818 ^ 1'b0 ;
  assign n5089 = ( n4818 & n4932 ) | ( n4818 & ~n5088 ) | ( n4932 & ~n5088 ) ;
  assign n5090 = ( n4818 & n4932 ) | ( n4818 & n5087 ) | ( n4932 & n5087 ) ;
  assign n5091 = n4950 ^ n4850 ^ 1'b0 ;
  assign n5092 = ( n4850 & n4967 ) | ( n4850 & ~n5091 ) | ( n4967 & ~n5091 ) ;
  assign n5093 = n4967 ^ n4948 ^ 1'b0 ;
  assign n5094 = ( n4850 & n4967 ) | ( n4850 & n5093 ) | ( n4967 & n5093 ) ;
  assign n5095 = n4948 ^ n4915 ^ 1'b0 ;
  assign n5096 = n4950 ^ n4743 ^ 1'b0 ;
  assign n5097 = ( n4743 & n4915 ) | ( n4743 & ~n5096 ) | ( n4915 & ~n5096 ) ;
  assign n5098 = ( n4743 & n4915 ) | ( n4743 & n5095 ) | ( n4915 & n5095 ) ;
  assign n5099 = n4948 ^ n4925 ^ 1'b0 ;
  assign n5100 = ( n4816 & n4925 ) | ( n4816 & n5099 ) | ( n4925 & n5099 ) ;
  assign n5101 = n4950 ^ n4816 ^ 1'b0 ;
  assign n5102 = ( n4816 & n4925 ) | ( n4816 & ~n5101 ) | ( n4925 & ~n5101 ) ;
  assign n5103 = n4950 ^ n4848 ^ 1'b0 ;
  assign n5104 = n5002 ^ n4948 ^ 1'b0 ;
  assign n5105 = ( n4848 & n5002 ) | ( n4848 & n5104 ) | ( n5002 & n5104 ) ;
  assign n5106 = ( n4848 & n5002 ) | ( n4848 & ~n5103 ) | ( n5002 & ~n5103 ) ;
  assign n5107 = n4948 ^ n4908 ^ 1'b0 ;
  assign n5108 = ( n4757 & n4908 ) | ( n4757 & n5107 ) | ( n4908 & n5107 ) ;
  assign n5109 = n4950 ^ n4757 ^ 1'b0 ;
  assign n5110 = ( n4757 & n4908 ) | ( n4757 & ~n5109 ) | ( n4908 & ~n5109 ) ;
  assign n5111 = n4948 ^ n4934 ^ 1'b0 ;
  assign n5112 = n4938 ^ n4853 ^ x105 ;
  assign n5113 = n4950 ^ n4781 ^ 1'b0 ;
  assign n5114 = ( n4781 & n4934 ) | ( n4781 & ~n5113 ) | ( n4934 & ~n5113 ) ;
  assign n5115 = ( n4781 & n4934 ) | ( n4781 & n5111 ) | ( n4934 & n5111 ) ;
  assign n5116 = n4950 ^ n4763 ^ 1'b0 ;
  assign n5117 = n4948 ^ n4904 ^ 1'b0 ;
  assign n5118 = ( n4763 & n4904 ) | ( n4763 & n5117 ) | ( n4904 & n5117 ) ;
  assign n5119 = ( n4763 & n4904 ) | ( n4763 & ~n5116 ) | ( n4904 & ~n5116 ) ;
  assign n5120 = n4950 ^ n4795 ^ 1'b0 ;
  assign n5121 = ( n4795 & n4929 ) | ( n4795 & ~n5120 ) | ( n4929 & ~n5120 ) ;
  assign n5122 = n4948 ^ n4929 ^ 1'b0 ;
  assign n5123 = ( n4795 & n4929 ) | ( n4795 & n5122 ) | ( n4929 & n5122 ) ;
  assign n5124 = n4948 ^ n4935 ^ 1'b0 ;
  assign n5125 = ( n4784 & n4935 ) | ( n4784 & n5124 ) | ( n4935 & n5124 ) ;
  assign n5126 = n4950 ^ n4784 ^ 1'b0 ;
  assign n5127 = ( n4784 & n4935 ) | ( n4784 & ~n5126 ) | ( n4935 & ~n5126 ) ;
  assign n5128 = n4950 ^ n4853 ^ 1'b0 ;
  assign n5129 = n5112 ^ n4948 ^ 1'b0 ;
  assign n5130 = ( n4853 & n5112 ) | ( n4853 & ~n5128 ) | ( n5112 & ~n5128 ) ;
  assign n5131 = ( n4853 & n5112 ) | ( n4853 & n5129 ) | ( n5112 & n5129 ) ;
  assign n5132 = x64 & n4948 ;
  assign n5133 = n5132 ^ x64 ^ x17 ;
  assign n5134 = ~x16 & x64 ;
  assign n5135 = n5134 ^ n5133 ^ x65 ;
  assign n5136 = ( x65 & n5134 ) | ( x65 & n5135 ) | ( n5134 & n5135 ) ;
  assign n5137 = n5136 ^ n5021 ^ x66 ;
  assign n5138 = ( x66 & n5136 ) | ( x66 & n5137 ) | ( n5136 & n5137 ) ;
  assign n5139 = ( x67 & ~n5029 ) | ( x67 & n5138 ) | ( ~n5029 & n5138 ) ;
  assign n5140 = n4948 ^ n4857 ^ 1'b0 ;
  assign n5141 = n5139 ^ n4962 ^ x68 ;
  assign n5142 = ( x68 & ~n4962 ) | ( x68 & n5139 ) | ( ~n4962 & n5139 ) ;
  assign n5143 = n5050 ^ n4948 ^ 1'b0 ;
  assign n5144 = n5078 ^ n4948 ^ 1'b0 ;
  assign n5145 = ( n4767 & n5078 ) | ( n4767 & n5144 ) | ( n5078 & n5144 ) ;
  assign n5146 = ( n4773 & n4857 ) | ( n4773 & n5140 ) | ( n4857 & n5140 ) ;
  assign n5147 = ( x69 & n5142 ) | ( x69 & ~n5146 ) | ( n5142 & ~n5146 ) ;
  assign n5148 = ( x70 & ~n5027 ) | ( x70 & n5147 ) | ( ~n5027 & n5147 ) ;
  assign n5149 = ( x71 & ~n4971 ) | ( x71 & n5148 ) | ( ~n4971 & n5148 ) ;
  assign n5150 = ( x72 & ~n5145 ) | ( x72 & n5149 ) | ( ~n5145 & n5149 ) ;
  assign n5151 = ( x73 & ~n5003 ) | ( x73 & n5150 ) | ( ~n5003 & n5150 ) ;
  assign n5152 = n4950 ^ n4773 ^ 1'b0 ;
  assign n5153 = ( n4759 & n5050 ) | ( n4759 & n5143 ) | ( n5050 & n5143 ) ;
  assign n5154 = ( x74 & ~n5118 ) | ( x74 & n5151 ) | ( ~n5118 & n5151 ) ;
  assign n5155 = ( x75 & ~n4972 ) | ( x75 & n5154 ) | ( ~n4972 & n5154 ) ;
  assign n5156 = n5155 ^ n5153 ^ x76 ;
  assign n5157 = ( x76 & ~n5153 ) | ( x76 & n5155 ) | ( ~n5153 & n5155 ) ;
  assign n5158 = ( x77 & ~n5108 ) | ( x77 & n5157 ) | ( ~n5108 & n5157 ) ;
  assign n5159 = ( x78 & ~n4981 ) | ( x78 & n5158 ) | ( ~n4981 & n5158 ) ;
  assign n5160 = ( x79 & ~n5053 ) | ( x79 & n5159 ) | ( ~n5053 & n5159 ) ;
  assign n5161 = ( x80 & ~n5034 ) | ( x80 & n5160 ) | ( ~n5034 & n5160 ) ;
  assign n5162 = ( x81 & ~n5013 ) | ( x81 & n5161 ) | ( ~n5013 & n5161 ) ;
  assign n5163 = n4950 ^ n4759 ^ 1'b0 ;
  assign n5164 = n5147 ^ n5027 ^ x70 ;
  assign n5165 = n5154 ^ n4972 ^ x75 ;
  assign n5166 = ( x82 & ~n5061 ) | ( x82 & n5162 ) | ( ~n5061 & n5162 ) ;
  assign n5167 = n5150 ^ n5003 ^ x73 ;
  assign n5168 = ( x83 & ~n4954 ) | ( x83 & n5166 ) | ( ~n4954 & n5166 ) ;
  assign n5169 = n5158 ^ n4981 ^ x78 ;
  assign n5170 = ( n4773 & n4857 ) | ( n4773 & ~n5152 ) | ( n4857 & ~n5152 ) ;
  assign n5171 = ( x84 & ~n5098 ) | ( x84 & n5168 ) | ( ~n5098 & n5168 ) ;
  assign n5172 = ( x85 & ~n5047 ) | ( x85 & n5171 ) | ( ~n5047 & n5171 ) ;
  assign n5173 = ( n4759 & n5050 ) | ( n4759 & ~n5163 ) | ( n5050 & ~n5163 ) ;
  assign n5174 = ( x86 & ~n5057 ) | ( x86 & n5172 ) | ( ~n5057 & n5172 ) ;
  assign n5175 = n4950 ^ n4767 ^ 1'b0 ;
  assign n5176 = n5162 ^ n5061 ^ x82 ;
  assign n5177 = n5166 ^ n4954 ^ x83 ;
  assign n5178 = n5151 ^ n5118 ^ x74 ;
  assign n5179 = ( n4767 & n5078 ) | ( n4767 & ~n5175 ) | ( n5078 & ~n5175 ) ;
  assign n5180 = ( x87 & ~n5008 ) | ( x87 & n5174 ) | ( ~n5008 & n5174 ) ;
  assign n5181 = n5174 ^ n5008 ^ x87 ;
  assign n5182 = ( x88 & ~n5085 ) | ( x88 & n5180 ) | ( ~n5085 & n5180 ) ;
  assign n5183 = n5138 ^ n5029 ^ x67 ;
  assign n5184 = ( x89 & ~n5077 ) | ( x89 & n5182 ) | ( ~n5077 & n5182 ) ;
  assign n5185 = ( x90 & ~n5082 ) | ( x90 & n5184 ) | ( ~n5082 & n5184 ) ;
  assign n5186 = ( x91 & ~n4996 ) | ( x91 & n5185 ) | ( ~n4996 & n5185 ) ;
  assign n5187 = ( x92 & ~n5016 ) | ( x92 & n5186 ) | ( ~n5016 & n5186 ) ;
  assign n5188 = ( x93 & ~n4976 ) | ( x93 & n5187 ) | ( ~n4976 & n5187 ) ;
  assign n5189 = ( x94 & ~n5063 ) | ( x94 & n5188 ) | ( ~n5063 & n5188 ) ;
  assign n5190 = ( x95 & ~n5000 ) | ( x95 & n5189 ) | ( ~n5000 & n5189 ) ;
  assign n5191 = ( x96 & ~n4991 ) | ( x96 & n5190 ) | ( ~n4991 & n5190 ) ;
  assign n5192 = ( x97 & ~n5073 ) | ( x97 & n5191 ) | ( ~n5073 & n5191 ) ;
  assign n5193 = ( x98 & ~n5123 ) | ( x98 & n5192 ) | ( ~n5123 & n5192 ) ;
  assign n5194 = ( x99 & ~n5011 ) | ( x99 & n5193 ) | ( ~n5011 & n5193 ) ;
  assign n5195 = ( x100 & ~n4986 ) | ( x100 & n5194 ) | ( ~n4986 & n5194 ) ;
  assign n5196 = ( x101 & ~n5090 ) | ( x101 & n5195 ) | ( ~n5090 & n5195 ) ;
  assign n5197 = ( x102 & ~n5100 ) | ( x102 & n5196 ) | ( ~n5100 & n5196 ) ;
  assign n5198 = ( x103 & ~n5125 ) | ( x103 & n5197 ) | ( ~n5125 & n5197 ) ;
  assign n5199 = ( x104 & ~n5115 ) | ( x104 & n5198 ) | ( ~n5115 & n5198 ) ;
  assign n5200 = ( x105 & ~n5044 ) | ( x105 & n5199 ) | ( ~n5044 & n5199 ) ;
  assign n5201 = ( x106 & ~n5131 ) | ( x106 & n5200 ) | ( ~n5131 & n5200 ) ;
  assign n5202 = ( x107 & ~n5094 ) | ( x107 & n5201 ) | ( ~n5094 & n5201 ) ;
  assign n5203 = ( x108 & ~n5105 ) | ( x108 & n5202 ) | ( ~n5105 & n5202 ) ;
  assign n5204 = ( x109 & ~n5040 ) | ( x109 & n5203 ) | ( ~n5040 & n5203 ) ;
  assign n5205 = n322 | n4956 ;
  assign n5206 = ( x110 & ~n5067 ) | ( x110 & n5204 ) | ( ~n5067 & n5204 ) ;
  assign n5207 = ( x111 & n5205 ) | ( x111 & ~n5206 ) | ( n5205 & ~n5206 ) ;
  assign n5208 = ( x111 & n4956 ) | ( x111 & n5206 ) | ( n4956 & n5206 ) ;
  assign n5209 = ( n183 & n5207 ) | ( n183 & ~n5208 ) | ( n5207 & ~n5208 ) ;
  assign n5210 = n5206 | n5209 ;
  assign n5211 = n1298 & n5205 ;
  assign n5212 = ( ~n5205 & n5210 ) | ( ~n5205 & n5211 ) | ( n5210 & n5211 ) ;
  assign n5213 = n5184 ^ n5082 ^ x90 ;
  assign n5214 = n5212 ^ n5082 ^ 1'b0 ;
  assign n5215 = ( n5082 & n5213 ) | ( n5082 & ~n5214 ) | ( n5213 & ~n5214 ) ;
  assign n5216 = n5182 ^ n5077 ^ x89 ;
  assign n5217 = n5212 ^ n5077 ^ 1'b0 ;
  assign n5218 = ( n5077 & n5216 ) | ( n5077 & ~n5217 ) | ( n5216 & ~n5217 ) ;
  assign n5219 = n5212 ^ n5008 ^ 1'b0 ;
  assign n5220 = ( n5008 & n5181 ) | ( n5008 & ~n5219 ) | ( n5181 & ~n5219 ) ;
  assign n5221 = n5212 ^ n4954 ^ 1'b0 ;
  assign n5222 = ( n4954 & n5177 ) | ( n4954 & ~n5221 ) | ( n5177 & ~n5221 ) ;
  assign n5223 = n5212 ^ n5061 ^ 1'b0 ;
  assign n5224 = ( n5061 & n5176 ) | ( n5061 & ~n5223 ) | ( n5176 & ~n5223 ) ;
  assign n5225 = n5212 ^ n4981 ^ 1'b0 ;
  assign n5226 = ( n4981 & n5169 ) | ( n4981 & ~n5225 ) | ( n5169 & ~n5225 ) ;
  assign n5227 = n5212 ^ n5153 ^ 1'b0 ;
  assign n5228 = ( n5153 & n5156 ) | ( n5153 & ~n5227 ) | ( n5156 & ~n5227 ) ;
  assign n5229 = n5212 ^ n4972 ^ 1'b0 ;
  assign n5230 = ( n4972 & n5165 ) | ( n4972 & ~n5229 ) | ( n5165 & ~n5229 ) ;
  assign n5231 = n5212 ^ n5118 ^ 1'b0 ;
  assign n5232 = ( n5118 & n5178 ) | ( n5118 & ~n5231 ) | ( n5178 & ~n5231 ) ;
  assign n5233 = n5212 ^ n5003 ^ 1'b0 ;
  assign n5234 = ( n5003 & n5167 ) | ( n5003 & ~n5233 ) | ( n5167 & ~n5233 ) ;
  assign n5235 = n5212 ^ n5027 ^ 1'b0 ;
  assign n5236 = ( n5027 & n5164 ) | ( n5027 & ~n5235 ) | ( n5164 & ~n5235 ) ;
  assign n5237 = n5212 ^ n4962 ^ 1'b0 ;
  assign n5238 = ( n4962 & n5141 ) | ( n4962 & ~n5237 ) | ( n5141 & ~n5237 ) ;
  assign n5239 = n5212 ^ n5029 ^ 1'b0 ;
  assign n5240 = ( n5029 & n5183 ) | ( n5029 & ~n5239 ) | ( n5183 & ~n5239 ) ;
  assign n5241 = n5212 ^ n5137 ^ 1'b0 ;
  assign n5242 = ( n5021 & n5137 ) | ( n5021 & n5241 ) | ( n5137 & n5241 ) ;
  assign n5243 = n5212 ^ n5135 ^ 1'b0 ;
  assign n5244 = ( n5133 & n5135 ) | ( n5133 & n5243 ) | ( n5135 & n5243 ) ;
  assign n5245 = ~n5210 & n5211 ;
  assign n5246 = ( n322 & n5211 ) | ( n322 & ~n5245 ) | ( n5211 & ~n5245 ) ;
  assign n5247 = n5201 ^ n5094 ^ x107 ;
  assign n5248 = n5212 ^ n5094 ^ 1'b0 ;
  assign n5249 = ( n5094 & n5247 ) | ( n5094 & ~n5248 ) | ( n5247 & ~n5248 ) ;
  assign n5250 = n5200 ^ n5131 ^ x106 ;
  assign n5251 = n5212 ^ n5131 ^ 1'b0 ;
  assign n5252 = ( n5131 & n5250 ) | ( n5131 & ~n5251 ) | ( n5250 & ~n5251 ) ;
  assign n5253 = n5198 ^ n5115 ^ x104 ;
  assign n5254 = n5212 ^ n5115 ^ 1'b0 ;
  assign n5255 = ( n5115 & n5253 ) | ( n5115 & ~n5254 ) | ( n5253 & ~n5254 ) ;
  assign n5256 = n5196 ^ n5100 ^ x102 ;
  assign n5257 = n5212 ^ n5100 ^ 1'b0 ;
  assign n5258 = ( n5100 & n5256 ) | ( n5100 & ~n5257 ) | ( n5256 & ~n5257 ) ;
  assign n5259 = n5195 ^ n5090 ^ x101 ;
  assign n5260 = n5212 ^ n5090 ^ 1'b0 ;
  assign n5261 = ( n5090 & n5259 ) | ( n5090 & ~n5260 ) | ( n5259 & ~n5260 ) ;
  assign n5262 = n5194 ^ n4986 ^ x100 ;
  assign n5263 = n5212 ^ n4986 ^ 1'b0 ;
  assign n5264 = ( n4986 & n5262 ) | ( n4986 & ~n5263 ) | ( n5262 & ~n5263 ) ;
  assign n5265 = n5193 ^ n5011 ^ x99 ;
  assign n5266 = n5212 ^ n5011 ^ 1'b0 ;
  assign n5267 = ( n5011 & n5265 ) | ( n5011 & ~n5266 ) | ( n5265 & ~n5266 ) ;
  assign n5268 = n5192 ^ n5123 ^ x98 ;
  assign n5269 = n5212 ^ n5123 ^ 1'b0 ;
  assign n5270 = ( n5123 & n5268 ) | ( n5123 & ~n5269 ) | ( n5268 & ~n5269 ) ;
  assign n5271 = n5190 ^ n4991 ^ x96 ;
  assign n5272 = n5212 ^ n4991 ^ 1'b0 ;
  assign n5273 = ( n4991 & n5271 ) | ( n4991 & ~n5272 ) | ( n5271 & ~n5272 ) ;
  assign n5274 = n5189 ^ n5000 ^ x95 ;
  assign n5275 = n5212 ^ n5000 ^ 1'b0 ;
  assign n5276 = ( n5000 & n5274 ) | ( n5000 & ~n5275 ) | ( n5274 & ~n5275 ) ;
  assign n5277 = n5188 ^ n5063 ^ x94 ;
  assign n5278 = n5212 ^ n5063 ^ 1'b0 ;
  assign n5279 = ( n5063 & n5277 ) | ( n5063 & ~n5278 ) | ( n5277 & ~n5278 ) ;
  assign n5280 = n5180 ^ n5085 ^ x88 ;
  assign n5281 = n5212 ^ n5085 ^ 1'b0 ;
  assign n5282 = ( n5085 & n5280 ) | ( n5085 & ~n5281 ) | ( n5280 & ~n5281 ) ;
  assign n5283 = n5168 ^ n5098 ^ x84 ;
  assign n5284 = n5212 ^ n5098 ^ 1'b0 ;
  assign n5285 = ( n5098 & n5283 ) | ( n5098 & ~n5284 ) | ( n5283 & ~n5284 ) ;
  assign n5286 = n5161 ^ n5013 ^ x81 ;
  assign n5287 = n5212 ^ n5013 ^ 1'b0 ;
  assign n5288 = ( n5013 & n5286 ) | ( n5013 & ~n5287 ) | ( n5286 & ~n5287 ) ;
  assign n5289 = n5159 ^ n5053 ^ x79 ;
  assign n5290 = n5212 ^ n5053 ^ 1'b0 ;
  assign n5291 = ( n5053 & n5289 ) | ( n5053 & ~n5290 ) | ( n5289 & ~n5290 ) ;
  assign n5292 = n5157 ^ n5108 ^ x77 ;
  assign n5293 = n5212 ^ n5108 ^ 1'b0 ;
  assign n5294 = ( n5108 & n5292 ) | ( n5108 & ~n5293 ) | ( n5292 & ~n5293 ) ;
  assign n5295 = n5148 ^ n4971 ^ x71 ;
  assign n5296 = n5212 ^ n4971 ^ 1'b0 ;
  assign n5297 = ( n4971 & n5295 ) | ( n4971 & ~n5296 ) | ( n5295 & ~n5296 ) ;
  assign n5298 = n1298 & n4966 ;
  assign n5299 = ( ~x111 & n183 ) | ( ~x111 & n4966 ) | ( n183 & n4966 ) ;
  assign n5300 = n5204 ^ n5067 ^ x110 ;
  assign n5301 = n5212 ^ n5067 ^ 1'b0 ;
  assign n5302 = ( n5067 & n5300 ) | ( n5067 & ~n5301 ) | ( n5300 & ~n5301 ) ;
  assign n5303 = n5203 ^ n5040 ^ x109 ;
  assign n5304 = n5212 ^ n5040 ^ 1'b0 ;
  assign n5305 = ( n5040 & n5303 ) | ( n5040 & ~n5304 ) | ( n5303 & ~n5304 ) ;
  assign n5306 = n5202 ^ n5105 ^ x108 ;
  assign n5307 = n5212 ^ n5105 ^ 1'b0 ;
  assign n5308 = ( n5105 & n5306 ) | ( n5105 & ~n5307 ) | ( n5306 & ~n5307 ) ;
  assign n5309 = n5199 ^ n5044 ^ x105 ;
  assign n5310 = n5212 ^ n5044 ^ 1'b0 ;
  assign n5311 = ( n5044 & n5309 ) | ( n5044 & ~n5310 ) | ( n5309 & ~n5310 ) ;
  assign n5312 = n5197 ^ n5125 ^ x103 ;
  assign n5313 = n5212 ^ n5125 ^ 1'b0 ;
  assign n5314 = ( n5125 & n5312 ) | ( n5125 & ~n5313 ) | ( n5312 & ~n5313 ) ;
  assign n5315 = n5191 ^ n5073 ^ x97 ;
  assign n5316 = n5212 ^ n5073 ^ 1'b0 ;
  assign n5317 = ( n5073 & n5315 ) | ( n5073 & ~n5316 ) | ( n5315 & ~n5316 ) ;
  assign n5318 = n5187 ^ n4976 ^ x93 ;
  assign n5319 = n5212 ^ n4976 ^ 1'b0 ;
  assign n5320 = ( n4976 & n5318 ) | ( n4976 & ~n5319 ) | ( n5318 & ~n5319 ) ;
  assign n5321 = n5186 ^ n5016 ^ x92 ;
  assign n5322 = n5212 ^ n5016 ^ 1'b0 ;
  assign n5323 = ( n5016 & n5321 ) | ( n5016 & ~n5322 ) | ( n5321 & ~n5322 ) ;
  assign n5324 = n5185 ^ n4996 ^ x91 ;
  assign n5325 = n5212 ^ n4996 ^ 1'b0 ;
  assign n5326 = ( n4996 & n5324 ) | ( n4996 & ~n5325 ) | ( n5324 & ~n5325 ) ;
  assign n5327 = n5172 ^ n5057 ^ x86 ;
  assign n5328 = n5212 ^ n5057 ^ 1'b0 ;
  assign n5329 = ( n5057 & n5327 ) | ( n5057 & ~n5328 ) | ( n5327 & ~n5328 ) ;
  assign n5330 = n5171 ^ n5047 ^ x85 ;
  assign n5331 = n5212 ^ n5047 ^ 1'b0 ;
  assign n5332 = ( n5047 & n5330 ) | ( n5047 & ~n5331 ) | ( n5330 & ~n5331 ) ;
  assign n5333 = n5160 ^ n5034 ^ x80 ;
  assign n5334 = n5212 ^ n5034 ^ 1'b0 ;
  assign n5335 = ( n5034 & n5333 ) | ( n5034 & ~n5334 ) | ( n5333 & ~n5334 ) ;
  assign n5336 = n5149 ^ n5145 ^ x72 ;
  assign n5337 = n5212 ^ n5145 ^ 1'b0 ;
  assign n5338 = ( n5145 & n5336 ) | ( n5145 & ~n5337 ) | ( n5336 & ~n5337 ) ;
  assign n5339 = n5146 ^ n5142 ^ x69 ;
  assign n5340 = n5212 ^ n5146 ^ 1'b0 ;
  assign n5341 = ( n5146 & n5339 ) | ( n5146 & ~n5340 ) | ( n5339 & ~n5340 ) ;
  assign n5342 = x64 & n5212 ;
  assign n5343 = x64 & n4950 ;
  assign n5344 = n5343 ^ x64 ^ x17 ;
  assign n5345 = n5344 ^ n5134 ^ x65 ;
  assign n5346 = ( x65 & n5134 ) | ( x65 & n5345 ) | ( n5134 & n5345 ) ;
  assign n5347 = n5346 ^ n5023 ^ x66 ;
  assign n5348 = ( x66 & n5346 ) | ( x66 & n5347 ) | ( n5346 & n5347 ) ;
  assign n5349 = ( x67 & ~n5032 ) | ( x67 & n5348 ) | ( ~n5032 & n5348 ) ;
  assign n5350 = ( x68 & ~n4963 ) | ( x68 & n5349 ) | ( ~n4963 & n5349 ) ;
  assign n5351 = ( x69 & ~n5170 ) | ( x69 & n5350 ) | ( ~n5170 & n5350 ) ;
  assign n5352 = ( x70 & ~n5025 ) | ( x70 & n5351 ) | ( ~n5025 & n5351 ) ;
  assign n5353 = ( x71 & ~n4959 ) | ( x71 & n5352 ) | ( ~n4959 & n5352 ) ;
  assign n5354 = ( x72 & ~n5179 ) | ( x72 & n5353 ) | ( ~n5179 & n5353 ) ;
  assign n5355 = ( x73 & ~n5014 ) | ( x73 & n5354 ) | ( ~n5014 & n5354 ) ;
  assign n5356 = ( x74 & ~n5119 ) | ( x74 & n5355 ) | ( ~n5119 & n5355 ) ;
  assign n5357 = ( x75 & ~n4977 ) | ( x75 & n5356 ) | ( ~n4977 & n5356 ) ;
  assign n5358 = ( x76 & ~n5173 ) | ( x76 & n5357 ) | ( ~n5173 & n5357 ) ;
  assign n5359 = ( x77 & ~n5110 ) | ( x77 & n5358 ) | ( ~n5110 & n5358 ) ;
  assign n5360 = ( x78 & ~n4980 ) | ( x78 & n5359 ) | ( ~n4980 & n5359 ) ;
  assign n5361 = ( x79 & ~n5051 ) | ( x79 & n5360 ) | ( ~n5051 & n5360 ) ;
  assign n5362 = ( x80 & ~n5036 ) | ( x80 & n5361 ) | ( ~n5036 & n5361 ) ;
  assign n5363 = ( x81 & ~n4974 ) | ( x81 & n5362 ) | ( ~n4974 & n5362 ) ;
  assign n5364 = ( x82 & ~n5060 ) | ( x82 & n5363 ) | ( ~n5060 & n5363 ) ;
  assign n5365 = ( x83 & ~n4952 ) | ( x83 & n5364 ) | ( ~n4952 & n5364 ) ;
  assign n5366 = ( x84 & ~n5097 ) | ( x84 & n5365 ) | ( ~n5097 & n5365 ) ;
  assign n5367 = ( x85 & ~n5048 ) | ( x85 & n5366 ) | ( ~n5048 & n5366 ) ;
  assign n5368 = ( x86 & ~n5056 ) | ( x86 & n5367 ) | ( ~n5056 & n5367 ) ;
  assign n5369 = ( x87 & ~n4993 ) | ( x87 & n5368 ) | ( ~n4993 & n5368 ) ;
  assign n5370 = ( x88 & ~n5086 ) | ( x88 & n5369 ) | ( ~n5086 & n5369 ) ;
  assign n5371 = n5364 ^ n4952 ^ x83 ;
  assign n5372 = n5363 ^ n5060 ^ x82 ;
  assign n5373 = n5360 ^ n5051 ^ x79 ;
  assign n5374 = n5359 ^ n4980 ^ x78 ;
  assign n5375 = n5357 ^ n5173 ^ x76 ;
  assign n5376 = ( x89 & ~n5076 ) | ( x89 & n5370 ) | ( ~n5076 & n5370 ) ;
  assign n5377 = ( x90 & ~n5080 ) | ( x90 & n5376 ) | ( ~n5080 & n5376 ) ;
  assign n5378 = n5352 ^ n4959 ^ x71 ;
  assign n5379 = ( x91 & ~n4998 ) | ( x91 & n5377 ) | ( ~n4998 & n5377 ) ;
  assign n5380 = n5379 ^ n5019 ^ x92 ;
  assign n5381 = n5369 ^ n5086 ^ x88 ;
  assign n5382 = ( x92 & ~n5019 ) | ( x92 & n5379 ) | ( ~n5019 & n5379 ) ;
  assign n5383 = n5376 ^ n5080 ^ x90 ;
  assign n5384 = n5370 ^ n5076 ^ x89 ;
  assign n5385 = ( x93 & ~n4988 ) | ( x93 & n5382 ) | ( ~n4988 & n5382 ) ;
  assign n5386 = ( x94 & ~n5065 ) | ( x94 & n5385 ) | ( ~n5065 & n5385 ) ;
  assign n5387 = n5355 ^ n5119 ^ x74 ;
  assign n5388 = ( x95 & ~n5004 ) | ( x95 & n5386 ) | ( ~n5004 & n5386 ) ;
  assign n5389 = n5388 ^ n4990 ^ x96 ;
  assign n5390 = ( x96 & ~n4990 ) | ( x96 & n5388 ) | ( ~n4990 & n5388 ) ;
  assign n5391 = ( x97 & ~n5072 ) | ( x97 & n5390 ) | ( ~n5072 & n5390 ) ;
  assign n5392 = ( x98 & ~n5121 ) | ( x98 & n5391 ) | ( ~n5121 & n5391 ) ;
  assign n5393 = ( x99 & ~n5007 ) | ( x99 & n5392 ) | ( ~n5007 & n5392 ) ;
  assign n5394 = ( x100 & ~n4984 ) | ( x100 & n5393 ) | ( ~n4984 & n5393 ) ;
  assign n5395 = ( x101 & ~n5089 ) | ( x101 & n5394 ) | ( ~n5089 & n5394 ) ;
  assign n5396 = ( x102 & ~n5102 ) | ( x102 & n5395 ) | ( ~n5102 & n5395 ) ;
  assign n5397 = ( x103 & ~n5127 ) | ( x103 & n5396 ) | ( ~n5127 & n5396 ) ;
  assign n5398 = ( x104 & ~n5114 ) | ( x104 & n5397 ) | ( ~n5114 & n5397 ) ;
  assign n5399 = ( x105 & ~n5042 ) | ( x105 & n5398 ) | ( ~n5042 & n5398 ) ;
  assign n5400 = ( x106 & ~n5130 ) | ( x106 & n5399 ) | ( ~n5130 & n5399 ) ;
  assign n5401 = n5349 ^ n4963 ^ x68 ;
  assign n5402 = ( x107 & ~n5092 ) | ( x107 & n5400 ) | ( ~n5092 & n5400 ) ;
  assign n5403 = ( x108 & ~n5106 ) | ( x108 & n5402 ) | ( ~n5106 & n5402 ) ;
  assign n5404 = ( x109 & ~n5038 ) | ( x109 & n5403 ) | ( ~n5038 & n5403 ) ;
  assign n5405 = ( x110 & ~n5069 ) | ( x110 & n5404 ) | ( ~n5069 & n5404 ) ;
  assign n5406 = n5405 ^ n4966 ^ x111 ;
  assign n5407 = n5398 ^ n5042 ^ x105 ;
  assign n5408 = ( x111 & ~n4966 ) | ( x111 & n5405 ) | ( ~n4966 & n5405 ) ;
  assign n5409 = n5299 | n5408 ;
  assign n5410 = ( ~n4966 & n5298 ) | ( ~n4966 & n5409 ) | ( n5298 & n5409 ) ;
  assign n5411 = n5410 ^ n5347 ^ 1'b0 ;
  assign n5412 = ( n5023 & n5347 ) | ( n5023 & n5411 ) | ( n5347 & n5411 ) ;
  assign n5413 = n5410 ^ n5173 ^ 1'b0 ;
  assign n5414 = n5391 ^ n5121 ^ x98 ;
  assign n5415 = n5410 ^ n5345 ^ 1'b0 ;
  assign n5416 = ( n5344 & n5345 ) | ( n5344 & n5415 ) | ( n5345 & n5415 ) ;
  assign n5417 = n5410 ^ n4990 ^ 1'b0 ;
  assign n5418 = n5410 ^ n4980 ^ 1'b0 ;
  assign n5419 = ( n5173 & n5375 ) | ( n5173 & ~n5413 ) | ( n5375 & ~n5413 ) ;
  assign n5420 = n5410 ^ n4959 ^ 1'b0 ;
  assign n5421 = ( n4959 & n5378 ) | ( n4959 & ~n5420 ) | ( n5378 & ~n5420 ) ;
  assign n5422 = n5410 ^ n5080 ^ 1'b0 ;
  assign n5423 = ( n4980 & n5374 ) | ( n4980 & ~n5418 ) | ( n5374 & ~n5418 ) ;
  assign n5424 = n5410 ^ n5042 ^ 1'b0 ;
  assign n5425 = ( n5080 & n5383 ) | ( n5080 & ~n5422 ) | ( n5383 & ~n5422 ) ;
  assign n5426 = n5410 ^ n4963 ^ 1'b0 ;
  assign n5427 = n5410 ^ n5121 ^ 1'b0 ;
  assign n5428 = ( n5121 & n5414 ) | ( n5121 & ~n5427 ) | ( n5414 & ~n5427 ) ;
  assign n5429 = n5410 ^ n5051 ^ 1'b0 ;
  assign n5430 = ( n5051 & n5373 ) | ( n5051 & ~n5429 ) | ( n5373 & ~n5429 ) ;
  assign n5431 = ( n4990 & n5389 ) | ( n4990 & ~n5417 ) | ( n5389 & ~n5417 ) ;
  assign n5432 = n5410 ^ n5119 ^ 1'b0 ;
  assign n5433 = ( n5119 & n5387 ) | ( n5119 & ~n5432 ) | ( n5387 & ~n5432 ) ;
  assign n5434 = n5410 ^ n5086 ^ 1'b0 ;
  assign n5435 = ( n4963 & n5401 ) | ( n4963 & ~n5426 ) | ( n5401 & ~n5426 ) ;
  assign n5436 = n5410 ^ n5019 ^ 1'b0 ;
  assign n5437 = ( n5086 & n5381 ) | ( n5086 & ~n5434 ) | ( n5381 & ~n5434 ) ;
  assign n5438 = n5410 ^ n5076 ^ 1'b0 ;
  assign n5439 = n5410 ^ n4952 ^ 1'b0 ;
  assign n5440 = ( n5019 & n5380 ) | ( n5019 & ~n5436 ) | ( n5380 & ~n5436 ) ;
  assign n5441 = n5298 & ~n5409 ;
  assign n5442 = ( n5042 & n5407 ) | ( n5042 & ~n5424 ) | ( n5407 & ~n5424 ) ;
  assign n5443 = ( n5076 & n5384 ) | ( n5076 & ~n5438 ) | ( n5384 & ~n5438 ) ;
  assign n5444 = n5406 & ~n5410 ;
  assign n5445 = n5410 ^ n5060 ^ 1'b0 ;
  assign n5446 = ( n5060 & n5372 ) | ( n5060 & ~n5445 ) | ( n5372 & ~n5445 ) ;
  assign n5447 = ( n5298 & ~n5441 ) | ( n5298 & n5444 ) | ( ~n5441 & n5444 ) ;
  assign n5448 = ( n4952 & n5371 ) | ( n4952 & ~n5439 ) | ( n5371 & ~n5439 ) ;
  assign n5449 = n5404 ^ n5069 ^ x110 ;
  assign n5450 = n5410 ^ n5069 ^ 1'b0 ;
  assign n5451 = ( n5069 & n5449 ) | ( n5069 & ~n5450 ) | ( n5449 & ~n5450 ) ;
  assign n5452 = n5377 ^ n4998 ^ x91 ;
  assign n5453 = n5410 ^ n4998 ^ 1'b0 ;
  assign n5454 = ( n4998 & n5452 ) | ( n4998 & ~n5453 ) | ( n5452 & ~n5453 ) ;
  assign n5455 = n5368 ^ n4993 ^ x87 ;
  assign n5456 = n5410 ^ n4993 ^ 1'b0 ;
  assign n5457 = ( n4993 & n5455 ) | ( n4993 & ~n5456 ) | ( n5455 & ~n5456 ) ;
  assign n5458 = n5367 ^ n5056 ^ x86 ;
  assign n5459 = n5410 ^ n5056 ^ 1'b0 ;
  assign n5460 = ( n5056 & n5458 ) | ( n5056 & ~n5459 ) | ( n5458 & ~n5459 ) ;
  assign n5461 = n5366 ^ n5048 ^ x85 ;
  assign n5462 = n5410 ^ n5048 ^ 1'b0 ;
  assign n5463 = ( n5048 & n5461 ) | ( n5048 & ~n5462 ) | ( n5461 & ~n5462 ) ;
  assign n5464 = n5365 ^ n5097 ^ x84 ;
  assign n5465 = n5410 ^ n5097 ^ 1'b0 ;
  assign n5466 = ( n5097 & n5464 ) | ( n5097 & ~n5465 ) | ( n5464 & ~n5465 ) ;
  assign n5467 = n5362 ^ n4974 ^ x81 ;
  assign n5468 = n5410 ^ n4974 ^ 1'b0 ;
  assign n5469 = ( n4974 & n5467 ) | ( n4974 & ~n5468 ) | ( n5467 & ~n5468 ) ;
  assign n5470 = n5361 ^ n5036 ^ x80 ;
  assign n5471 = n5410 ^ n5036 ^ 1'b0 ;
  assign n5472 = ( n5036 & n5470 ) | ( n5036 & ~n5471 ) | ( n5470 & ~n5471 ) ;
  assign n5473 = n5358 ^ n5110 ^ x77 ;
  assign n5474 = n5410 ^ n5110 ^ 1'b0 ;
  assign n5475 = ( n5110 & n5473 ) | ( n5110 & ~n5474 ) | ( n5473 & ~n5474 ) ;
  assign n5476 = n5356 ^ n4977 ^ x75 ;
  assign n5477 = n5410 ^ n4977 ^ 1'b0 ;
  assign n5478 = ( n4977 & n5476 ) | ( n4977 & ~n5477 ) | ( n5476 & ~n5477 ) ;
  assign n5479 = n5354 ^ n5014 ^ x73 ;
  assign n5480 = n5410 ^ n5014 ^ 1'b0 ;
  assign n5481 = ( n5014 & n5479 ) | ( n5014 & ~n5480 ) | ( n5479 & ~n5480 ) ;
  assign n5482 = n5353 ^ n5179 ^ x72 ;
  assign n5483 = n5410 ^ n5179 ^ 1'b0 ;
  assign n5484 = ( n5179 & n5482 ) | ( n5179 & ~n5483 ) | ( n5482 & ~n5483 ) ;
  assign n5485 = n5351 ^ n5025 ^ x70 ;
  assign n5486 = n5410 ^ n5025 ^ 1'b0 ;
  assign n5487 = ( n5025 & n5485 ) | ( n5025 & ~n5486 ) | ( n5485 & ~n5486 ) ;
  assign n5488 = n5350 ^ n5170 ^ x69 ;
  assign n5489 = n5410 ^ n5170 ^ 1'b0 ;
  assign n5490 = ( n5170 & n5488 ) | ( n5170 & ~n5489 ) | ( n5488 & ~n5489 ) ;
  assign n5491 = n5348 ^ n5032 ^ x67 ;
  assign n5492 = n5410 ^ n5032 ^ 1'b0 ;
  assign n5493 = ( n5032 & n5491 ) | ( n5032 & ~n5492 ) | ( n5491 & ~n5492 ) ;
  assign n5494 = n5403 ^ n5038 ^ x109 ;
  assign n5495 = n5410 ^ n5038 ^ 1'b0 ;
  assign n5496 = ( n5038 & n5494 ) | ( n5038 & ~n5495 ) | ( n5494 & ~n5495 ) ;
  assign n5497 = n5402 ^ n5106 ^ x108 ;
  assign n5498 = n5410 ^ n5106 ^ 1'b0 ;
  assign n5499 = ( n5106 & n5497 ) | ( n5106 & ~n5498 ) | ( n5497 & ~n5498 ) ;
  assign n5500 = n5400 ^ n5092 ^ x107 ;
  assign n5501 = n5410 ^ n5092 ^ 1'b0 ;
  assign n5502 = ( n5092 & n5500 ) | ( n5092 & ~n5501 ) | ( n5500 & ~n5501 ) ;
  assign n5503 = n5399 ^ n5130 ^ x106 ;
  assign n5504 = n5410 ^ n5130 ^ 1'b0 ;
  assign n5505 = ( n5130 & n5503 ) | ( n5130 & ~n5504 ) | ( n5503 & ~n5504 ) ;
  assign n5506 = n5397 ^ n5114 ^ x104 ;
  assign n5507 = n5410 ^ n5114 ^ 1'b0 ;
  assign n5508 = ( n5114 & n5506 ) | ( n5114 & ~n5507 ) | ( n5506 & ~n5507 ) ;
  assign n5509 = n5396 ^ n5127 ^ x103 ;
  assign n5510 = n5410 ^ n5127 ^ 1'b0 ;
  assign n5511 = ( n5127 & n5509 ) | ( n5127 & ~n5510 ) | ( n5509 & ~n5510 ) ;
  assign n5512 = n5395 ^ n5102 ^ x102 ;
  assign n5513 = n5410 ^ n5102 ^ 1'b0 ;
  assign n5514 = ( n5102 & n5512 ) | ( n5102 & ~n5513 ) | ( n5512 & ~n5513 ) ;
  assign n5515 = n5394 ^ n5089 ^ x101 ;
  assign n5516 = n5410 ^ n5089 ^ 1'b0 ;
  assign n5517 = ( n5089 & n5515 ) | ( n5089 & ~n5516 ) | ( n5515 & ~n5516 ) ;
  assign n5518 = n5393 ^ n4984 ^ x100 ;
  assign n5519 = n5410 ^ n4984 ^ 1'b0 ;
  assign n5520 = ( n4984 & n5518 ) | ( n4984 & ~n5519 ) | ( n5518 & ~n5519 ) ;
  assign n5521 = n5392 ^ n5007 ^ x99 ;
  assign n5522 = n5410 ^ n5007 ^ 1'b0 ;
  assign n5523 = ( n5007 & n5521 ) | ( n5007 & ~n5522 ) | ( n5521 & ~n5522 ) ;
  assign n5524 = n5390 ^ n5072 ^ x97 ;
  assign n5525 = n5410 ^ n5072 ^ 1'b0 ;
  assign n5526 = ( n5072 & n5524 ) | ( n5072 & ~n5525 ) | ( n5524 & ~n5525 ) ;
  assign n5527 = n5386 ^ n5004 ^ x95 ;
  assign n5528 = n5410 ^ n5004 ^ 1'b0 ;
  assign n5529 = ( n5004 & n5527 ) | ( n5004 & ~n5528 ) | ( n5527 & ~n5528 ) ;
  assign n5530 = n5385 ^ n5065 ^ x94 ;
  assign n5531 = n5410 ^ n5065 ^ 1'b0 ;
  assign n5532 = ( n5065 & n5530 ) | ( n5065 & ~n5531 ) | ( n5530 & ~n5531 ) ;
  assign n5533 = n5382 ^ n4988 ^ x93 ;
  assign n5534 = n5410 ^ n4988 ^ 1'b0 ;
  assign n5535 = ( n4988 & n5533 ) | ( n4988 & ~n5534 ) | ( n5533 & ~n5534 ) ;
  assign n5536 = n5342 ^ x64 ^ x16 ;
  assign n5537 = ~x15 & x64 ;
  assign n5538 = n5537 ^ n5536 ^ x65 ;
  assign n5539 = ( x65 & n5537 ) | ( x65 & n5538 ) | ( n5537 & n5538 ) ;
  assign n5540 = n5539 ^ n5244 ^ x66 ;
  assign n5541 = ( x66 & n5539 ) | ( x66 & n5540 ) | ( n5539 & n5540 ) ;
  assign n5542 = ( x67 & ~n5242 ) | ( x67 & n5541 ) | ( ~n5242 & n5541 ) ;
  assign n5543 = ( x68 & ~n5240 ) | ( x68 & n5542 ) | ( ~n5240 & n5542 ) ;
  assign n5544 = ( x69 & ~n5238 ) | ( x69 & n5543 ) | ( ~n5238 & n5543 ) ;
  assign n5545 = ( x70 & ~n5341 ) | ( x70 & n5544 ) | ( ~n5341 & n5544 ) ;
  assign n5546 = ( x71 & ~n5236 ) | ( x71 & n5545 ) | ( ~n5236 & n5545 ) ;
  assign n5547 = ( x72 & ~n5297 ) | ( x72 & n5546 ) | ( ~n5297 & n5546 ) ;
  assign n5548 = ( x73 & ~n5338 ) | ( x73 & n5547 ) | ( ~n5338 & n5547 ) ;
  assign n5549 = ( x74 & ~n5234 ) | ( x74 & n5548 ) | ( ~n5234 & n5548 ) ;
  assign n5550 = ( x75 & ~n5232 ) | ( x75 & n5549 ) | ( ~n5232 & n5549 ) ;
  assign n5551 = ( x76 & ~n5230 ) | ( x76 & n5550 ) | ( ~n5230 & n5550 ) ;
  assign n5552 = ( x77 & ~n5228 ) | ( x77 & n5551 ) | ( ~n5228 & n5551 ) ;
  assign n5553 = ( x78 & ~n5294 ) | ( x78 & n5552 ) | ( ~n5294 & n5552 ) ;
  assign n5554 = ( x79 & ~n5226 ) | ( x79 & n5553 ) | ( ~n5226 & n5553 ) ;
  assign n5555 = ( x80 & ~n5291 ) | ( x80 & n5554 ) | ( ~n5291 & n5554 ) ;
  assign n5556 = ( x81 & ~n5335 ) | ( x81 & n5555 ) | ( ~n5335 & n5555 ) ;
  assign n5557 = ( x82 & ~n5288 ) | ( x82 & n5556 ) | ( ~n5288 & n5556 ) ;
  assign n5558 = ( x83 & ~n5224 ) | ( x83 & n5557 ) | ( ~n5224 & n5557 ) ;
  assign n5559 = ( x84 & ~n5222 ) | ( x84 & n5558 ) | ( ~n5222 & n5558 ) ;
  assign n5560 = ( x85 & ~n5285 ) | ( x85 & n5559 ) | ( ~n5285 & n5559 ) ;
  assign n5561 = ( x86 & ~n5332 ) | ( x86 & n5560 ) | ( ~n5332 & n5560 ) ;
  assign n5562 = ( x87 & ~n5329 ) | ( x87 & n5561 ) | ( ~n5329 & n5561 ) ;
  assign n5563 = ( x88 & ~n5220 ) | ( x88 & n5562 ) | ( ~n5220 & n5562 ) ;
  assign n5564 = ( x89 & ~n5282 ) | ( x89 & n5563 ) | ( ~n5282 & n5563 ) ;
  assign n5565 = ( x90 & ~n5218 ) | ( x90 & n5564 ) | ( ~n5218 & n5564 ) ;
  assign n5566 = ( x91 & ~n5215 ) | ( x91 & n5565 ) | ( ~n5215 & n5565 ) ;
  assign n5567 = n5553 ^ n5226 ^ x79 ;
  assign n5568 = ( x92 & ~n5326 ) | ( x92 & n5566 ) | ( ~n5326 & n5566 ) ;
  assign n5569 = n5552 ^ n5294 ^ x78 ;
  assign n5570 = n5556 ^ n5288 ^ x82 ;
  assign n5571 = n5557 ^ n5224 ^ x83 ;
  assign n5572 = n5558 ^ n5222 ^ x84 ;
  assign n5573 = ( x93 & ~n5323 ) | ( x93 & n5568 ) | ( ~n5323 & n5568 ) ;
  assign n5574 = n5560 ^ n5332 ^ x86 ;
  assign n5575 = ( x94 & ~n5320 ) | ( x94 & n5573 ) | ( ~n5320 & n5573 ) ;
  assign n5576 = n5563 ^ n5282 ^ x89 ;
  assign n5577 = n5568 ^ n5323 ^ x93 ;
  assign n5578 = n5564 ^ n5218 ^ x90 ;
  assign n5579 = n5550 ^ n5230 ^ x76 ;
  assign n5580 = n5549 ^ n5232 ^ x75 ;
  assign n5581 = n5543 ^ n5238 ^ x69 ;
  assign n5582 = n5542 ^ n5240 ^ x68 ;
  assign n5583 = n5541 ^ n5242 ^ x67 ;
  assign n5584 = ( x95 & ~n5279 ) | ( x95 & n5575 ) | ( ~n5279 & n5575 ) ;
  assign n5585 = ( x96 & ~n5276 ) | ( x96 & n5584 ) | ( ~n5276 & n5584 ) ;
  assign n5586 = ( x97 & ~n5273 ) | ( x97 & n5585 ) | ( ~n5273 & n5585 ) ;
  assign n5587 = ( x98 & ~n5317 ) | ( x98 & n5586 ) | ( ~n5317 & n5586 ) ;
  assign n5588 = ( x99 & ~n5270 ) | ( x99 & n5587 ) | ( ~n5270 & n5587 ) ;
  assign n5589 = ( x100 & ~n5267 ) | ( x100 & n5588 ) | ( ~n5267 & n5588 ) ;
  assign n5590 = ( x101 & ~n5264 ) | ( x101 & n5589 ) | ( ~n5264 & n5589 ) ;
  assign n5591 = ( x102 & ~n5261 ) | ( x102 & n5590 ) | ( ~n5261 & n5590 ) ;
  assign n5592 = ( x103 & ~n5258 ) | ( x103 & n5591 ) | ( ~n5258 & n5591 ) ;
  assign n5593 = ( x104 & ~n5314 ) | ( x104 & n5592 ) | ( ~n5314 & n5592 ) ;
  assign n5594 = ( x105 & ~n5255 ) | ( x105 & n5593 ) | ( ~n5255 & n5593 ) ;
  assign n5595 = ( x106 & ~n5311 ) | ( x106 & n5594 ) | ( ~n5311 & n5594 ) ;
  assign n5596 = ( x107 & ~n5252 ) | ( x107 & n5595 ) | ( ~n5252 & n5595 ) ;
  assign n5597 = ( x108 & ~n5249 ) | ( x108 & n5596 ) | ( ~n5249 & n5596 ) ;
  assign n5598 = ( x109 & ~n5308 ) | ( x109 & n5597 ) | ( ~n5308 & n5597 ) ;
  assign n5599 = ( x110 & ~n5305 ) | ( x110 & n5598 ) | ( ~n5305 & n5598 ) ;
  assign n5600 = ( x111 & ~n5302 ) | ( x111 & n5599 ) | ( ~n5302 & n5599 ) ;
  assign n5601 = ( x112 & ~n5246 ) | ( x112 & n5600 ) | ( ~n5246 & n5600 ) ;
  assign n5602 = n158 | n5601 ;
  assign n5603 = n5585 ^ n5273 ^ x97 ;
  assign n5604 = n5602 ^ n5273 ^ 1'b0 ;
  assign n5605 = ( n5273 & n5603 ) | ( n5273 & ~n5604 ) | ( n5603 & ~n5604 ) ;
  assign n5606 = n5573 ^ n5320 ^ x94 ;
  assign n5607 = n5602 ^ n5320 ^ 1'b0 ;
  assign n5608 = ( n5320 & n5606 ) | ( n5320 & ~n5607 ) | ( n5606 & ~n5607 ) ;
  assign n5609 = n5602 ^ n5323 ^ 1'b0 ;
  assign n5610 = ( n5323 & n5577 ) | ( n5323 & ~n5609 ) | ( n5577 & ~n5609 ) ;
  assign n5611 = n5602 ^ n5218 ^ 1'b0 ;
  assign n5612 = ( n5218 & n5578 ) | ( n5218 & ~n5611 ) | ( n5578 & ~n5611 ) ;
  assign n5613 = n5602 ^ n5282 ^ 1'b0 ;
  assign n5614 = ( n5282 & n5576 ) | ( n5282 & ~n5613 ) | ( n5576 & ~n5613 ) ;
  assign n5615 = n5602 ^ n5332 ^ 1'b0 ;
  assign n5616 = ( n5332 & n5574 ) | ( n5332 & ~n5615 ) | ( n5574 & ~n5615 ) ;
  assign n5617 = n5602 ^ n5222 ^ 1'b0 ;
  assign n5618 = ( n5222 & n5572 ) | ( n5222 & ~n5617 ) | ( n5572 & ~n5617 ) ;
  assign n5619 = n5602 ^ n5224 ^ 1'b0 ;
  assign n5620 = ( n5224 & n5571 ) | ( n5224 & ~n5619 ) | ( n5571 & ~n5619 ) ;
  assign n5621 = n5602 ^ n5288 ^ 1'b0 ;
  assign n5622 = ( n5288 & n5570 ) | ( n5288 & ~n5621 ) | ( n5570 & ~n5621 ) ;
  assign n5623 = n5602 ^ n5226 ^ 1'b0 ;
  assign n5624 = ( n5226 & n5567 ) | ( n5226 & ~n5623 ) | ( n5567 & ~n5623 ) ;
  assign n5625 = n5602 ^ n5294 ^ 1'b0 ;
  assign n5626 = ( n5294 & n5569 ) | ( n5294 & ~n5625 ) | ( n5569 & ~n5625 ) ;
  assign n5627 = n5602 ^ n5230 ^ 1'b0 ;
  assign n5628 = ( n5230 & n5579 ) | ( n5230 & ~n5627 ) | ( n5579 & ~n5627 ) ;
  assign n5629 = n5602 ^ n5232 ^ 1'b0 ;
  assign n5630 = ( n5232 & n5580 ) | ( n5232 & ~n5629 ) | ( n5580 & ~n5629 ) ;
  assign n5631 = n5602 ^ n5238 ^ 1'b0 ;
  assign n5632 = ( n5238 & n5581 ) | ( n5238 & ~n5631 ) | ( n5581 & ~n5631 ) ;
  assign n5633 = n5602 ^ n5240 ^ 1'b0 ;
  assign n5634 = ( n5240 & n5582 ) | ( n5240 & ~n5633 ) | ( n5582 & ~n5633 ) ;
  assign n5635 = n5602 ^ n5242 ^ 1'b0 ;
  assign n5636 = ( n5242 & n5583 ) | ( n5242 & ~n5635 ) | ( n5583 & ~n5635 ) ;
  assign n5637 = n5602 ^ n5540 ^ 1'b0 ;
  assign n5638 = ( n5244 & n5540 ) | ( n5244 & n5637 ) | ( n5540 & n5637 ) ;
  assign n5639 = n5602 ^ n5538 ^ 1'b0 ;
  assign n5640 = ( n5536 & n5538 ) | ( n5536 & n5639 ) | ( n5538 & n5639 ) ;
  assign n5641 = n5599 ^ n5302 ^ x111 ;
  assign n5642 = n5602 ^ n5302 ^ 1'b0 ;
  assign n5643 = ( n5302 & n5641 ) | ( n5302 & ~n5642 ) | ( n5641 & ~n5642 ) ;
  assign n5644 = n5598 ^ n5305 ^ x110 ;
  assign n5645 = n5602 ^ n5305 ^ 1'b0 ;
  assign n5646 = ( n5305 & n5644 ) | ( n5305 & ~n5645 ) | ( n5644 & ~n5645 ) ;
  assign n5647 = n5575 ^ n5279 ^ x95 ;
  assign n5648 = n5602 ^ n5279 ^ 1'b0 ;
  assign n5649 = ( n5279 & n5647 ) | ( n5279 & ~n5648 ) | ( n5647 & ~n5648 ) ;
  assign n5650 = n5566 ^ n5326 ^ x92 ;
  assign n5651 = n5602 ^ n5326 ^ 1'b0 ;
  assign n5652 = ( n5326 & n5650 ) | ( n5326 & ~n5651 ) | ( n5650 & ~n5651 ) ;
  assign n5653 = n5565 ^ n5215 ^ x91 ;
  assign n5654 = n5602 ^ n5215 ^ 1'b0 ;
  assign n5655 = ( n5215 & n5653 ) | ( n5215 & ~n5654 ) | ( n5653 & ~n5654 ) ;
  assign n5656 = n5562 ^ n5220 ^ x88 ;
  assign n5657 = n5602 ^ n5220 ^ 1'b0 ;
  assign n5658 = ( n5220 & n5656 ) | ( n5220 & ~n5657 ) | ( n5656 & ~n5657 ) ;
  assign n5659 = n5561 ^ n5329 ^ x87 ;
  assign n5660 = n5602 ^ n5329 ^ 1'b0 ;
  assign n5661 = ( n5329 & n5659 ) | ( n5329 & ~n5660 ) | ( n5659 & ~n5660 ) ;
  assign n5662 = n5559 ^ n5285 ^ x85 ;
  assign n5663 = n5602 ^ n5285 ^ 1'b0 ;
  assign n5664 = ( n5285 & n5662 ) | ( n5285 & ~n5663 ) | ( n5662 & ~n5663 ) ;
  assign n5665 = n5555 ^ n5335 ^ x81 ;
  assign n5666 = n5602 ^ n5335 ^ 1'b0 ;
  assign n5667 = ( n5335 & n5665 ) | ( n5335 & ~n5666 ) | ( n5665 & ~n5666 ) ;
  assign n5668 = n5554 ^ n5291 ^ x80 ;
  assign n5669 = n5602 ^ n5291 ^ 1'b0 ;
  assign n5670 = ( n5291 & n5668 ) | ( n5291 & ~n5669 ) | ( n5668 & ~n5669 ) ;
  assign n5671 = n5551 ^ n5228 ^ x77 ;
  assign n5672 = n5602 ^ n5228 ^ 1'b0 ;
  assign n5673 = ( n5228 & n5671 ) | ( n5228 & ~n5672 ) | ( n5671 & ~n5672 ) ;
  assign n5674 = n5548 ^ n5234 ^ x74 ;
  assign n5675 = n5602 ^ n5234 ^ 1'b0 ;
  assign n5676 = ( n5234 & n5674 ) | ( n5234 & ~n5675 ) | ( n5674 & ~n5675 ) ;
  assign n5677 = n5547 ^ n5338 ^ x73 ;
  assign n5678 = n5602 ^ n5338 ^ 1'b0 ;
  assign n5679 = ( n5338 & n5677 ) | ( n5338 & ~n5678 ) | ( n5677 & ~n5678 ) ;
  assign n5680 = n5546 ^ n5297 ^ x72 ;
  assign n5681 = n5602 ^ n5297 ^ 1'b0 ;
  assign n5682 = ( n5297 & n5680 ) | ( n5297 & ~n5681 ) | ( n5680 & ~n5681 ) ;
  assign n5683 = n5545 ^ n5236 ^ x71 ;
  assign n5684 = n5602 ^ n5236 ^ 1'b0 ;
  assign n5685 = ( n5236 & n5683 ) | ( n5236 & ~n5684 ) | ( n5683 & ~n5684 ) ;
  assign n5686 = n5544 ^ n5341 ^ x70 ;
  assign n5687 = n5602 ^ n5341 ^ 1'b0 ;
  assign n5688 = ( n5341 & n5686 ) | ( n5341 & ~n5687 ) | ( n5686 & ~n5687 ) ;
  assign n5689 = n5597 ^ n5308 ^ x109 ;
  assign n5690 = n5602 ^ n5308 ^ 1'b0 ;
  assign n5691 = ( n5308 & n5689 ) | ( n5308 & ~n5690 ) | ( n5689 & ~n5690 ) ;
  assign n5692 = n5596 ^ n5249 ^ x108 ;
  assign n5693 = n5602 ^ n5249 ^ 1'b0 ;
  assign n5694 = ( n5249 & n5692 ) | ( n5249 & ~n5693 ) | ( n5692 & ~n5693 ) ;
  assign n5695 = n5595 ^ n5252 ^ x107 ;
  assign n5696 = n5602 ^ n5252 ^ 1'b0 ;
  assign n5697 = ( n5252 & n5695 ) | ( n5252 & ~n5696 ) | ( n5695 & ~n5696 ) ;
  assign n5698 = n5594 ^ n5311 ^ x106 ;
  assign n5699 = n5602 ^ n5311 ^ 1'b0 ;
  assign n5700 = ( n5311 & n5698 ) | ( n5311 & ~n5699 ) | ( n5698 & ~n5699 ) ;
  assign n5701 = n5593 ^ n5255 ^ x105 ;
  assign n5702 = n5602 ^ n5255 ^ 1'b0 ;
  assign n5703 = ( n5255 & n5701 ) | ( n5255 & ~n5702 ) | ( n5701 & ~n5702 ) ;
  assign n5704 = n5592 ^ n5314 ^ x104 ;
  assign n5705 = n5602 ^ n5314 ^ 1'b0 ;
  assign n5706 = ( n5314 & n5704 ) | ( n5314 & ~n5705 ) | ( n5704 & ~n5705 ) ;
  assign n5707 = n5591 ^ n5258 ^ x103 ;
  assign n5708 = n5602 ^ n5258 ^ 1'b0 ;
  assign n5709 = ( n5258 & n5707 ) | ( n5258 & ~n5708 ) | ( n5707 & ~n5708 ) ;
  assign n5710 = n5590 ^ n5261 ^ x102 ;
  assign n5711 = n5602 ^ n5261 ^ 1'b0 ;
  assign n5712 = ( n5261 & n5710 ) | ( n5261 & ~n5711 ) | ( n5710 & ~n5711 ) ;
  assign n5713 = n5589 ^ n5264 ^ x101 ;
  assign n5714 = n5602 ^ n5264 ^ 1'b0 ;
  assign n5715 = ( n5264 & n5713 ) | ( n5264 & ~n5714 ) | ( n5713 & ~n5714 ) ;
  assign n5716 = n5588 ^ n5267 ^ x100 ;
  assign n5717 = n5602 ^ n5267 ^ 1'b0 ;
  assign n5718 = ( n5267 & n5716 ) | ( n5267 & ~n5717 ) | ( n5716 & ~n5717 ) ;
  assign n5719 = n5587 ^ n5270 ^ x99 ;
  assign n5720 = n5602 ^ n5270 ^ 1'b0 ;
  assign n5721 = ( n5270 & n5719 ) | ( n5270 & ~n5720 ) | ( n5719 & ~n5720 ) ;
  assign n5722 = n5586 ^ n5317 ^ x98 ;
  assign n5723 = n5602 ^ n5317 ^ 1'b0 ;
  assign n5724 = ( n5317 & n5722 ) | ( n5317 & ~n5723 ) | ( n5722 & ~n5723 ) ;
  assign n5725 = n5584 ^ n5276 ^ x96 ;
  assign n5726 = n5602 ^ n5276 ^ 1'b0 ;
  assign n5727 = ( n5276 & n5725 ) | ( n5276 & ~n5726 ) | ( n5725 & ~n5726 ) ;
  assign n5728 = n5246 & n5602 ;
  assign n5729 = n158 & n5246 ;
  assign n5730 = ( ~x114 & x115 ) | ( ~x114 & n174 ) | ( x115 & n174 ) ;
  assign n5731 = x114 | n5730 ;
  assign n5732 = ~x14 & x64 ;
  assign n5733 = x64 & ~x113 ;
  assign n5734 = ~n5731 & n5733 ;
  assign n5735 = x15 & ~n5734 ;
  assign n5736 = ~n158 & n5537 ;
  assign n5737 = n5601 | n5736 ;
  assign n5738 = ( x15 & ~n5601 ) | ( x15 & n5737 ) | ( ~n5601 & n5737 ) ;
  assign n5739 = ( n5735 & n5737 ) | ( n5735 & n5738 ) | ( n5737 & n5738 ) ;
  assign n5740 = n5739 ^ n5732 ^ x65 ;
  assign n5741 = ( x65 & n5732 ) | ( x65 & n5740 ) | ( n5732 & n5740 ) ;
  assign n5742 = n5741 ^ n5640 ^ x66 ;
  assign n5743 = ( x66 & n5741 ) | ( x66 & n5742 ) | ( n5741 & n5742 ) ;
  assign n5744 = ( x67 & ~n5638 ) | ( x67 & n5743 ) | ( ~n5638 & n5743 ) ;
  assign n5745 = ( x68 & ~n5636 ) | ( x68 & n5744 ) | ( ~n5636 & n5744 ) ;
  assign n5746 = ( x69 & ~n5634 ) | ( x69 & n5745 ) | ( ~n5634 & n5745 ) ;
  assign n5747 = ( x70 & ~n5632 ) | ( x70 & n5746 ) | ( ~n5632 & n5746 ) ;
  assign n5748 = ( x71 & ~n5688 ) | ( x71 & n5747 ) | ( ~n5688 & n5747 ) ;
  assign n5749 = ( x72 & ~n5685 ) | ( x72 & n5748 ) | ( ~n5685 & n5748 ) ;
  assign n5750 = ( x73 & ~n5682 ) | ( x73 & n5749 ) | ( ~n5682 & n5749 ) ;
  assign n5751 = ( x74 & ~n5679 ) | ( x74 & n5750 ) | ( ~n5679 & n5750 ) ;
  assign n5752 = ( x75 & ~n5676 ) | ( x75 & n5751 ) | ( ~n5676 & n5751 ) ;
  assign n5753 = ( x76 & ~n5630 ) | ( x76 & n5752 ) | ( ~n5630 & n5752 ) ;
  assign n5754 = ( x77 & ~n5628 ) | ( x77 & n5753 ) | ( ~n5628 & n5753 ) ;
  assign n5755 = ( x78 & ~n5673 ) | ( x78 & n5754 ) | ( ~n5673 & n5754 ) ;
  assign n5756 = ( x79 & ~n5626 ) | ( x79 & n5755 ) | ( ~n5626 & n5755 ) ;
  assign n5757 = ( x80 & ~n5624 ) | ( x80 & n5756 ) | ( ~n5624 & n5756 ) ;
  assign n5758 = ( x81 & ~n5670 ) | ( x81 & n5757 ) | ( ~n5670 & n5757 ) ;
  assign n5759 = ( x82 & ~n5667 ) | ( x82 & n5758 ) | ( ~n5667 & n5758 ) ;
  assign n5760 = ( x83 & ~n5622 ) | ( x83 & n5759 ) | ( ~n5622 & n5759 ) ;
  assign n5761 = ( x84 & ~n5620 ) | ( x84 & n5760 ) | ( ~n5620 & n5760 ) ;
  assign n5762 = ( x85 & ~n5618 ) | ( x85 & n5761 ) | ( ~n5618 & n5761 ) ;
  assign n5763 = ( x86 & ~n5664 ) | ( x86 & n5762 ) | ( ~n5664 & n5762 ) ;
  assign n5764 = ( x87 & ~n5616 ) | ( x87 & n5763 ) | ( ~n5616 & n5763 ) ;
  assign n5765 = ( x88 & ~n5661 ) | ( x88 & n5764 ) | ( ~n5661 & n5764 ) ;
  assign n5766 = ( x89 & ~n5658 ) | ( x89 & n5765 ) | ( ~n5658 & n5765 ) ;
  assign n5767 = ( x90 & ~n5614 ) | ( x90 & n5766 ) | ( ~n5614 & n5766 ) ;
  assign n5768 = ( x91 & ~n5612 ) | ( x91 & n5767 ) | ( ~n5612 & n5767 ) ;
  assign n5769 = ( x92 & ~n5655 ) | ( x92 & n5768 ) | ( ~n5655 & n5768 ) ;
  assign n5770 = ( x93 & ~n5652 ) | ( x93 & n5769 ) | ( ~n5652 & n5769 ) ;
  assign n5771 = n5758 ^ n5667 ^ x82 ;
  assign n5772 = n5757 ^ n5670 ^ x81 ;
  assign n5773 = n5763 ^ n5616 ^ x87 ;
  assign n5774 = ( x94 & ~n5610 ) | ( x94 & n5770 ) | ( ~n5610 & n5770 ) ;
  assign n5775 = n322 | n5728 ;
  assign n5776 = n5770 ^ n5610 ^ x94 ;
  assign n5777 = n5753 ^ n5628 ^ x77 ;
  assign n5778 = n5752 ^ n5630 ^ x76 ;
  assign n5779 = n5749 ^ n5682 ^ x73 ;
  assign n5780 = n5747 ^ n5688 ^ x71 ;
  assign n5781 = n5743 ^ n5638 ^ x67 ;
  assign n5782 = ( x95 & ~n5608 ) | ( x95 & n5774 ) | ( ~n5608 & n5774 ) ;
  assign n5783 = ( x96 & ~n5649 ) | ( x96 & n5782 ) | ( ~n5649 & n5782 ) ;
  assign n5784 = ( x97 & ~n5727 ) | ( x97 & n5783 ) | ( ~n5727 & n5783 ) ;
  assign n5785 = ( x98 & ~n5605 ) | ( x98 & n5784 ) | ( ~n5605 & n5784 ) ;
  assign n5786 = ( x99 & ~n5724 ) | ( x99 & n5785 ) | ( ~n5724 & n5785 ) ;
  assign n5787 = ( x100 & ~n5721 ) | ( x100 & n5786 ) | ( ~n5721 & n5786 ) ;
  assign n5788 = ( x101 & ~n5718 ) | ( x101 & n5787 ) | ( ~n5718 & n5787 ) ;
  assign n5789 = ( x102 & ~n5715 ) | ( x102 & n5788 ) | ( ~n5715 & n5788 ) ;
  assign n5790 = ( x103 & ~n5712 ) | ( x103 & n5789 ) | ( ~n5712 & n5789 ) ;
  assign n5791 = ( x104 & ~n5709 ) | ( x104 & n5790 ) | ( ~n5709 & n5790 ) ;
  assign n5792 = ( x105 & ~n5706 ) | ( x105 & n5791 ) | ( ~n5706 & n5791 ) ;
  assign n5793 = ( x106 & ~n5703 ) | ( x106 & n5792 ) | ( ~n5703 & n5792 ) ;
  assign n5794 = ( x107 & ~n5700 ) | ( x107 & n5793 ) | ( ~n5700 & n5793 ) ;
  assign n5795 = ( x108 & ~n5697 ) | ( x108 & n5794 ) | ( ~n5697 & n5794 ) ;
  assign n5796 = ( x109 & ~n5694 ) | ( x109 & n5795 ) | ( ~n5694 & n5795 ) ;
  assign n5797 = ( x110 & ~n5691 ) | ( x110 & n5796 ) | ( ~n5691 & n5796 ) ;
  assign n5798 = ( x111 & ~n5646 ) | ( x111 & n5797 ) | ( ~n5646 & n5797 ) ;
  assign n5799 = n5798 ^ n5643 ^ x112 ;
  assign n5800 = ( x112 & ~n5643 ) | ( x112 & n5798 ) | ( ~n5643 & n5798 ) ;
  assign n5801 = ( x113 & n5775 ) | ( x113 & ~n5800 ) | ( n5775 & ~n5800 ) ;
  assign n5802 = ( x113 & n5728 ) | ( x113 & n5800 ) | ( n5728 & n5800 ) ;
  assign n5803 = ( n5731 & n5801 ) | ( n5731 & ~n5802 ) | ( n5801 & ~n5802 ) ;
  assign n5804 = n5800 | n5803 ;
  assign n5805 = n158 & n5775 ;
  assign n5806 = ( ~n5775 & n5804 ) | ( ~n5775 & n5805 ) | ( n5804 & n5805 ) ;
  assign n5807 = n5796 ^ n5691 ^ x110 ;
  assign n5808 = n5806 ^ n5691 ^ 1'b0 ;
  assign n5809 = ( n5691 & n5807 ) | ( n5691 & ~n5808 ) | ( n5807 & ~n5808 ) ;
  assign n5810 = n5795 ^ n5694 ^ x109 ;
  assign n5811 = n5806 ^ n5694 ^ 1'b0 ;
  assign n5812 = ( n5694 & n5810 ) | ( n5694 & ~n5811 ) | ( n5810 & ~n5811 ) ;
  assign n5813 = n5786 ^ n5721 ^ x100 ;
  assign n5814 = n5806 ^ n5721 ^ 1'b0 ;
  assign n5815 = ( n5721 & n5813 ) | ( n5721 & ~n5814 ) | ( n5813 & ~n5814 ) ;
  assign n5816 = n5806 ^ n5643 ^ 1'b0 ;
  assign n5817 = ( n5643 & n5799 ) | ( n5643 & ~n5816 ) | ( n5799 & ~n5816 ) ;
  assign n5818 = n5782 ^ n5649 ^ x96 ;
  assign n5819 = n5806 ^ n5649 ^ 1'b0 ;
  assign n5820 = ( n5649 & n5818 ) | ( n5649 & ~n5819 ) | ( n5818 & ~n5819 ) ;
  assign n5821 = n5806 ^ n5610 ^ 1'b0 ;
  assign n5822 = ( n5610 & n5776 ) | ( n5610 & ~n5821 ) | ( n5776 & ~n5821 ) ;
  assign n5823 = n5806 ^ n5616 ^ 1'b0 ;
  assign n5824 = ( n5616 & n5773 ) | ( n5616 & ~n5823 ) | ( n5773 & ~n5823 ) ;
  assign n5825 = n5806 ^ n5667 ^ 1'b0 ;
  assign n5826 = ( n5667 & n5771 ) | ( n5667 & ~n5825 ) | ( n5771 & ~n5825 ) ;
  assign n5827 = n5806 ^ n5670 ^ 1'b0 ;
  assign n5828 = ( n5670 & n5772 ) | ( n5670 & ~n5827 ) | ( n5772 & ~n5827 ) ;
  assign n5829 = n5806 ^ n5628 ^ 1'b0 ;
  assign n5830 = ( n5628 & n5777 ) | ( n5628 & ~n5829 ) | ( n5777 & ~n5829 ) ;
  assign n5831 = n5806 ^ n5630 ^ 1'b0 ;
  assign n5832 = ( n5630 & n5778 ) | ( n5630 & ~n5831 ) | ( n5778 & ~n5831 ) ;
  assign n5833 = n5806 ^ n5682 ^ 1'b0 ;
  assign n5834 = ( n5682 & n5779 ) | ( n5682 & ~n5833 ) | ( n5779 & ~n5833 ) ;
  assign n5835 = n5806 ^ n5688 ^ 1'b0 ;
  assign n5836 = ( n5688 & n5780 ) | ( n5688 & ~n5835 ) | ( n5780 & ~n5835 ) ;
  assign n5837 = n5806 ^ n5638 ^ 1'b0 ;
  assign n5838 = ( n5638 & n5781 ) | ( n5638 & ~n5837 ) | ( n5781 & ~n5837 ) ;
  assign n5839 = n5806 ^ n5742 ^ 1'b0 ;
  assign n5840 = ( n5640 & n5742 ) | ( n5640 & n5839 ) | ( n5742 & n5839 ) ;
  assign n5841 = n5806 ^ n5740 ^ 1'b0 ;
  assign n5842 = ( n5739 & n5740 ) | ( n5739 & n5841 ) | ( n5740 & n5841 ) ;
  assign n5843 = n5729 & n5804 ;
  assign n5844 = n5797 ^ n5646 ^ x111 ;
  assign n5845 = n5806 ^ n5646 ^ 1'b0 ;
  assign n5846 = ( n5646 & n5844 ) | ( n5646 & ~n5845 ) | ( n5844 & ~n5845 ) ;
  assign n5847 = n5794 ^ n5697 ^ x108 ;
  assign n5848 = n5806 ^ n5697 ^ 1'b0 ;
  assign n5849 = ( n5697 & n5847 ) | ( n5697 & ~n5848 ) | ( n5847 & ~n5848 ) ;
  assign n5850 = n5765 ^ n5658 ^ x89 ;
  assign n5851 = n5806 ^ n5658 ^ 1'b0 ;
  assign n5852 = ( n5658 & n5850 ) | ( n5658 & ~n5851 ) | ( n5850 & ~n5851 ) ;
  assign n5853 = n5764 ^ n5661 ^ x88 ;
  assign n5854 = n5806 ^ n5661 ^ 1'b0 ;
  assign n5855 = ( n5661 & n5853 ) | ( n5661 & ~n5854 ) | ( n5853 & ~n5854 ) ;
  assign n5856 = n5762 ^ n5664 ^ x86 ;
  assign n5857 = n5806 ^ n5664 ^ 1'b0 ;
  assign n5858 = ( n5664 & n5856 ) | ( n5664 & ~n5857 ) | ( n5856 & ~n5857 ) ;
  assign n5859 = n5761 ^ n5618 ^ x85 ;
  assign n5860 = n5806 ^ n5618 ^ 1'b0 ;
  assign n5861 = ( n5618 & n5859 ) | ( n5618 & ~n5860 ) | ( n5859 & ~n5860 ) ;
  assign n5862 = n5760 ^ n5620 ^ x84 ;
  assign n5863 = n5806 ^ n5620 ^ 1'b0 ;
  assign n5864 = ( n5620 & n5862 ) | ( n5620 & ~n5863 ) | ( n5862 & ~n5863 ) ;
  assign n5865 = n5759 ^ n5622 ^ x83 ;
  assign n5866 = n5806 ^ n5622 ^ 1'b0 ;
  assign n5867 = ( n5622 & n5865 ) | ( n5622 & ~n5866 ) | ( n5865 & ~n5866 ) ;
  assign n5868 = n5756 ^ n5624 ^ x80 ;
  assign n5869 = n5806 ^ n5624 ^ 1'b0 ;
  assign n5870 = ( n5624 & n5868 ) | ( n5624 & ~n5869 ) | ( n5868 & ~n5869 ) ;
  assign n5871 = n5755 ^ n5626 ^ x79 ;
  assign n5872 = n5806 ^ n5626 ^ 1'b0 ;
  assign n5873 = ( n5626 & n5871 ) | ( n5626 & ~n5872 ) | ( n5871 & ~n5872 ) ;
  assign n5874 = n5754 ^ n5673 ^ x78 ;
  assign n5875 = n5806 ^ n5673 ^ 1'b0 ;
  assign n5876 = ( n5673 & n5874 ) | ( n5673 & ~n5875 ) | ( n5874 & ~n5875 ) ;
  assign n5877 = n5751 ^ n5676 ^ x75 ;
  assign n5878 = n5806 ^ n5676 ^ 1'b0 ;
  assign n5879 = ( n5676 & n5877 ) | ( n5676 & ~n5878 ) | ( n5877 & ~n5878 ) ;
  assign n5880 = n5750 ^ n5679 ^ x74 ;
  assign n5881 = n5806 ^ n5679 ^ 1'b0 ;
  assign n5882 = ( n5679 & n5880 ) | ( n5679 & ~n5881 ) | ( n5880 & ~n5881 ) ;
  assign n5883 = n5748 ^ n5685 ^ x72 ;
  assign n5884 = n5806 ^ n5685 ^ 1'b0 ;
  assign n5885 = ( n5685 & n5883 ) | ( n5685 & ~n5884 ) | ( n5883 & ~n5884 ) ;
  assign n5886 = n5746 ^ n5632 ^ x70 ;
  assign n5887 = n5806 ^ n5632 ^ 1'b0 ;
  assign n5888 = ( n5632 & n5886 ) | ( n5632 & ~n5887 ) | ( n5886 & ~n5887 ) ;
  assign n5889 = n5745 ^ n5634 ^ x69 ;
  assign n5890 = n5806 ^ n5634 ^ 1'b0 ;
  assign n5891 = ( n5634 & n5889 ) | ( n5634 & ~n5890 ) | ( n5889 & ~n5890 ) ;
  assign n5892 = n5744 ^ n5636 ^ x68 ;
  assign n5893 = n5806 ^ n5636 ^ 1'b0 ;
  assign n5894 = ( n5636 & n5892 ) | ( n5636 & ~n5893 ) | ( n5892 & ~n5893 ) ;
  assign n5895 = n5793 ^ n5700 ^ x107 ;
  assign n5896 = n5806 ^ n5700 ^ 1'b0 ;
  assign n5897 = ( n5700 & n5895 ) | ( n5700 & ~n5896 ) | ( n5895 & ~n5896 ) ;
  assign n5898 = n5792 ^ n5703 ^ x106 ;
  assign n5899 = n5806 ^ n5703 ^ 1'b0 ;
  assign n5900 = ( n5703 & n5898 ) | ( n5703 & ~n5899 ) | ( n5898 & ~n5899 ) ;
  assign n5901 = n5791 ^ n5706 ^ x105 ;
  assign n5902 = n5806 ^ n5706 ^ 1'b0 ;
  assign n5903 = ( n5706 & n5901 ) | ( n5706 & ~n5902 ) | ( n5901 & ~n5902 ) ;
  assign n5904 = n5790 ^ n5709 ^ x104 ;
  assign n5905 = n5806 ^ n5709 ^ 1'b0 ;
  assign n5906 = ( n5709 & n5904 ) | ( n5709 & ~n5905 ) | ( n5904 & ~n5905 ) ;
  assign n5907 = n5789 ^ n5712 ^ x103 ;
  assign n5908 = n5806 ^ n5712 ^ 1'b0 ;
  assign n5909 = ( n5712 & n5907 ) | ( n5712 & ~n5908 ) | ( n5907 & ~n5908 ) ;
  assign n5910 = n5788 ^ n5715 ^ x102 ;
  assign n5911 = n5806 ^ n5715 ^ 1'b0 ;
  assign n5912 = ( n5715 & n5910 ) | ( n5715 & ~n5911 ) | ( n5910 & ~n5911 ) ;
  assign n5913 = n5787 ^ n5718 ^ x101 ;
  assign n5914 = n5806 ^ n5718 ^ 1'b0 ;
  assign n5915 = ( n5718 & n5913 ) | ( n5718 & ~n5914 ) | ( n5913 & ~n5914 ) ;
  assign n5916 = n5785 ^ n5724 ^ x99 ;
  assign n5917 = n5806 ^ n5724 ^ 1'b0 ;
  assign n5918 = ( n5724 & n5916 ) | ( n5724 & ~n5917 ) | ( n5916 & ~n5917 ) ;
  assign n5919 = n5784 ^ n5605 ^ x98 ;
  assign n5920 = n5806 ^ n5605 ^ 1'b0 ;
  assign n5921 = ( n5605 & n5919 ) | ( n5605 & ~n5920 ) | ( n5919 & ~n5920 ) ;
  assign n5922 = n5783 ^ n5727 ^ x97 ;
  assign n5923 = n5806 ^ n5727 ^ 1'b0 ;
  assign n5924 = ( n5727 & n5922 ) | ( n5727 & ~n5923 ) | ( n5922 & ~n5923 ) ;
  assign n5925 = n5774 ^ n5608 ^ x95 ;
  assign n5926 = n5806 ^ n5608 ^ 1'b0 ;
  assign n5927 = ( n5608 & n5925 ) | ( n5608 & ~n5926 ) | ( n5925 & ~n5926 ) ;
  assign n5928 = n5769 ^ n5652 ^ x93 ;
  assign n5929 = n5806 ^ n5652 ^ 1'b0 ;
  assign n5930 = ( n5652 & n5928 ) | ( n5652 & ~n5929 ) | ( n5928 & ~n5929 ) ;
  assign n5931 = n5768 ^ n5655 ^ x92 ;
  assign n5932 = n5806 ^ n5655 ^ 1'b0 ;
  assign n5933 = ( n5655 & n5931 ) | ( n5655 & ~n5932 ) | ( n5931 & ~n5932 ) ;
  assign n5934 = n5767 ^ n5612 ^ x91 ;
  assign n5935 = n5806 ^ n5612 ^ 1'b0 ;
  assign n5936 = ( n5612 & n5934 ) | ( n5612 & ~n5935 ) | ( n5934 & ~n5935 ) ;
  assign n5937 = n5766 ^ n5614 ^ x90 ;
  assign n5938 = n5806 ^ n5614 ^ 1'b0 ;
  assign n5939 = ( n5614 & n5937 ) | ( n5614 & ~n5938 ) | ( n5937 & ~n5938 ) ;
  assign n5940 = x64 & n5410 ;
  assign n5941 = n5940 ^ x64 ^ x16 ;
  assign n5942 = n5941 ^ n5537 ^ x65 ;
  assign n5943 = ( x65 & n5537 ) | ( x65 & n5942 ) | ( n5537 & n5942 ) ;
  assign n5944 = n5943 ^ n5416 ^ x66 ;
  assign n5945 = ( x66 & n5943 ) | ( x66 & n5944 ) | ( n5943 & n5944 ) ;
  assign n5946 = ( x67 & ~n5412 ) | ( x67 & n5945 ) | ( ~n5412 & n5945 ) ;
  assign n5947 = ( x68 & ~n5493 ) | ( x68 & n5946 ) | ( ~n5493 & n5946 ) ;
  assign n5948 = ( x69 & ~n5435 ) | ( x69 & n5947 ) | ( ~n5435 & n5947 ) ;
  assign n5949 = ( x70 & ~n5490 ) | ( x70 & n5948 ) | ( ~n5490 & n5948 ) ;
  assign n5950 = ( x71 & ~n5487 ) | ( x71 & n5949 ) | ( ~n5487 & n5949 ) ;
  assign n5951 = ( x72 & ~n5421 ) | ( x72 & n5950 ) | ( ~n5421 & n5950 ) ;
  assign n5952 = ( x73 & ~n5484 ) | ( x73 & n5951 ) | ( ~n5484 & n5951 ) ;
  assign n5953 = ( x74 & ~n5481 ) | ( x74 & n5952 ) | ( ~n5481 & n5952 ) ;
  assign n5954 = ( x75 & ~n5433 ) | ( x75 & n5953 ) | ( ~n5433 & n5953 ) ;
  assign n5955 = ( x76 & ~n5478 ) | ( x76 & n5954 ) | ( ~n5478 & n5954 ) ;
  assign n5956 = ( x77 & ~n5419 ) | ( x77 & n5955 ) | ( ~n5419 & n5955 ) ;
  assign n5957 = ( x78 & ~n5475 ) | ( x78 & n5956 ) | ( ~n5475 & n5956 ) ;
  assign n5958 = ( x79 & ~n5423 ) | ( x79 & n5957 ) | ( ~n5423 & n5957 ) ;
  assign n5959 = ( x80 & ~n5430 ) | ( x80 & n5958 ) | ( ~n5430 & n5958 ) ;
  assign n5960 = ( x81 & ~n5472 ) | ( x81 & n5959 ) | ( ~n5472 & n5959 ) ;
  assign n5961 = ( x82 & ~n5469 ) | ( x82 & n5960 ) | ( ~n5469 & n5960 ) ;
  assign n5962 = ( x83 & ~n5446 ) | ( x83 & n5961 ) | ( ~n5446 & n5961 ) ;
  assign n5963 = ( x84 & ~n5448 ) | ( x84 & n5962 ) | ( ~n5448 & n5962 ) ;
  assign n5964 = ( x85 & ~n5466 ) | ( x85 & n5963 ) | ( ~n5466 & n5963 ) ;
  assign n5965 = ( x86 & ~n5463 ) | ( x86 & n5964 ) | ( ~n5463 & n5964 ) ;
  assign n5966 = ( x87 & ~n5460 ) | ( x87 & n5965 ) | ( ~n5460 & n5965 ) ;
  assign n5967 = ( x88 & ~n5457 ) | ( x88 & n5966 ) | ( ~n5457 & n5966 ) ;
  assign n5968 = ( x89 & ~n5437 ) | ( x89 & n5967 ) | ( ~n5437 & n5967 ) ;
  assign n5969 = ( x90 & ~n5443 ) | ( x90 & n5968 ) | ( ~n5443 & n5968 ) ;
  assign n5970 = ( x91 & ~n5425 ) | ( x91 & n5969 ) | ( ~n5425 & n5969 ) ;
  assign n5971 = ( x92 & ~n5454 ) | ( x92 & n5970 ) | ( ~n5454 & n5970 ) ;
  assign n5972 = ( x93 & ~n5440 ) | ( x93 & n5971 ) | ( ~n5440 & n5971 ) ;
  assign n5973 = ( x94 & ~n5535 ) | ( x94 & n5972 ) | ( ~n5535 & n5972 ) ;
  assign n5974 = ( x95 & ~n5532 ) | ( x95 & n5973 ) | ( ~n5532 & n5973 ) ;
  assign n5975 = n5961 ^ n5446 ^ x83 ;
  assign n5976 = n5962 ^ n5448 ^ x84 ;
  assign n5977 = n5960 ^ n5469 ^ x82 ;
  assign n5978 = n5964 ^ n5463 ^ x86 ;
  assign n5979 = n5963 ^ n5466 ^ x85 ;
  assign n5980 = n5958 ^ n5430 ^ x80 ;
  assign n5981 = n5957 ^ n5423 ^ x79 ;
  assign n5982 = n5956 ^ n5475 ^ x78 ;
  assign n5983 = n5954 ^ n5478 ^ x76 ;
  assign n5984 = n5950 ^ n5421 ^ x72 ;
  assign n5985 = n5949 ^ n5487 ^ x71 ;
  assign n5986 = n5972 ^ n5535 ^ x94 ;
  assign n5987 = n5973 ^ n5532 ^ x95 ;
  assign n5988 = n5974 ^ n5529 ^ x96 ;
  assign n5989 = ( x96 & ~n5529 ) | ( x96 & n5974 ) | ( ~n5529 & n5974 ) ;
  assign n5990 = ( x97 & ~n5431 ) | ( x97 & n5989 ) | ( ~n5431 & n5989 ) ;
  assign n5991 = ( x98 & ~n5526 ) | ( x98 & n5990 ) | ( ~n5526 & n5990 ) ;
  assign n5992 = ( x99 & ~n5428 ) | ( x99 & n5991 ) | ( ~n5428 & n5991 ) ;
  assign n5993 = ( x100 & ~n5523 ) | ( x100 & n5992 ) | ( ~n5523 & n5992 ) ;
  assign n5994 = ( x101 & ~n5520 ) | ( x101 & n5993 ) | ( ~n5520 & n5993 ) ;
  assign n5995 = ( x102 & ~n5517 ) | ( x102 & n5994 ) | ( ~n5517 & n5994 ) ;
  assign n5996 = ( x103 & ~n5514 ) | ( x103 & n5995 ) | ( ~n5514 & n5995 ) ;
  assign n5997 = ( x104 & ~n5511 ) | ( x104 & n5996 ) | ( ~n5511 & n5996 ) ;
  assign n5998 = ( x105 & ~n5508 ) | ( x105 & n5997 ) | ( ~n5508 & n5997 ) ;
  assign n5999 = ( x106 & ~n5442 ) | ( x106 & n5998 ) | ( ~n5442 & n5998 ) ;
  assign n6000 = ( x107 & ~n5505 ) | ( x107 & n5999 ) | ( ~n5505 & n5999 ) ;
  assign n6001 = ( x108 & ~n5502 ) | ( x108 & n6000 ) | ( ~n5502 & n6000 ) ;
  assign n6002 = ( x109 & ~n5499 ) | ( x109 & n6001 ) | ( ~n5499 & n6001 ) ;
  assign n6003 = ( x110 & ~n5496 ) | ( x110 & n6002 ) | ( ~n5496 & n6002 ) ;
  assign n6004 = ( x111 & ~n5451 ) | ( x111 & n6003 ) | ( ~n5451 & n6003 ) ;
  assign n6005 = ( x112 & ~n5447 ) | ( x112 & n6004 ) | ( ~n5447 & n6004 ) ;
  assign n6006 = n158 | n6005 ;
  assign n6007 = n5736 | n6005 ;
  assign n6008 = ( x15 & ~n6005 ) | ( x15 & n6007 ) | ( ~n6005 & n6007 ) ;
  assign n6009 = ~n5734 & n6008 ;
  assign n6010 = n5992 ^ n5523 ^ x100 ;
  assign n6011 = ( n6007 & n6008 ) | ( n6007 & n6009 ) | ( n6008 & n6009 ) ;
  assign n6012 = n6006 ^ n5466 ^ 1'b0 ;
  assign n6013 = ( n5466 & n5979 ) | ( n5466 & ~n6012 ) | ( n5979 & ~n6012 ) ;
  assign n6014 = n6006 ^ n5535 ^ 1'b0 ;
  assign n6015 = n6006 ^ n5430 ^ 1'b0 ;
  assign n6016 = n6006 ^ n5421 ^ 1'b0 ;
  assign n6017 = ( n5421 & n5984 ) | ( n5421 & ~n6016 ) | ( n5984 & ~n6016 ) ;
  assign n6018 = ( n5430 & n5980 ) | ( n5430 & ~n6015 ) | ( n5980 & ~n6015 ) ;
  assign n6019 = n6006 ^ n5523 ^ 1'b0 ;
  assign n6020 = ( n5535 & n5986 ) | ( n5535 & ~n6014 ) | ( n5986 & ~n6014 ) ;
  assign n6021 = n6006 ^ n5944 ^ 1'b0 ;
  assign n6022 = n6006 ^ n5529 ^ 1'b0 ;
  assign n6023 = n6006 ^ n5478 ^ 1'b0 ;
  assign n6024 = n6006 ^ n5448 ^ 1'b0 ;
  assign n6025 = ( n5529 & n5988 ) | ( n5529 & ~n6022 ) | ( n5988 & ~n6022 ) ;
  assign n6026 = ( n5478 & n5983 ) | ( n5478 & ~n6023 ) | ( n5983 & ~n6023 ) ;
  assign n6027 = n5991 ^ n5428 ^ x99 ;
  assign n6028 = n6006 ^ n5428 ^ 1'b0 ;
  assign n6029 = ( n5428 & n6027 ) | ( n5428 & ~n6028 ) | ( n6027 & ~n6028 ) ;
  assign n6030 = ( n5416 & n5944 ) | ( n5416 & n6021 ) | ( n5944 & n6021 ) ;
  assign n6031 = n6006 ^ n5487 ^ 1'b0 ;
  assign n6032 = n6006 ^ n5463 ^ 1'b0 ;
  assign n6033 = n6006 ^ n5423 ^ 1'b0 ;
  assign n6034 = ( n5423 & n5981 ) | ( n5423 & ~n6033 ) | ( n5981 & ~n6033 ) ;
  assign n6035 = n6006 ^ n5532 ^ 1'b0 ;
  assign n6036 = n6006 ^ n5446 ^ 1'b0 ;
  assign n6037 = n6006 ^ n5475 ^ 1'b0 ;
  assign n6038 = ( n5475 & n5982 ) | ( n5475 & ~n6037 ) | ( n5982 & ~n6037 ) ;
  assign n6039 = n6006 ^ n5942 ^ 1'b0 ;
  assign n6040 = ( n5941 & n5942 ) | ( n5941 & n6039 ) | ( n5942 & n6039 ) ;
  assign n6041 = n6006 ^ n5469 ^ 1'b0 ;
  assign n6042 = ( n5469 & n5977 ) | ( n5469 & ~n6041 ) | ( n5977 & ~n6041 ) ;
  assign n6043 = ( n5448 & n5976 ) | ( n5448 & ~n6024 ) | ( n5976 & ~n6024 ) ;
  assign n6044 = ( n5532 & n5987 ) | ( n5532 & ~n6035 ) | ( n5987 & ~n6035 ) ;
  assign n6045 = ( n5523 & n6010 ) | ( n5523 & ~n6019 ) | ( n6010 & ~n6019 ) ;
  assign n6046 = ( n5487 & n5985 ) | ( n5487 & ~n6031 ) | ( n5985 & ~n6031 ) ;
  assign n6047 = ( n5463 & n5978 ) | ( n5463 & ~n6032 ) | ( n5978 & ~n6032 ) ;
  assign n6048 = ( n5446 & n5975 ) | ( n5446 & ~n6036 ) | ( n5975 & ~n6036 ) ;
  assign n6049 = n6002 ^ n5496 ^ x110 ;
  assign n6050 = n6006 ^ n5496 ^ 1'b0 ;
  assign n6051 = ( n5496 & n6049 ) | ( n5496 & ~n6050 ) | ( n6049 & ~n6050 ) ;
  assign n6052 = n6001 ^ n5499 ^ x109 ;
  assign n6053 = n6006 ^ n5499 ^ 1'b0 ;
  assign n6054 = ( n5499 & n6052 ) | ( n5499 & ~n6053 ) | ( n6052 & ~n6053 ) ;
  assign n6055 = n5999 ^ n5505 ^ x107 ;
  assign n6056 = n6006 ^ n5505 ^ 1'b0 ;
  assign n6057 = ( n5505 & n6055 ) | ( n5505 & ~n6056 ) | ( n6055 & ~n6056 ) ;
  assign n6058 = n5996 ^ n5511 ^ x104 ;
  assign n6059 = n6006 ^ n5511 ^ 1'b0 ;
  assign n6060 = ( n5511 & n6058 ) | ( n5511 & ~n6059 ) | ( n6058 & ~n6059 ) ;
  assign n6061 = n5995 ^ n5514 ^ x103 ;
  assign n6062 = n6006 ^ n5514 ^ 1'b0 ;
  assign n6063 = ( n5514 & n6061 ) | ( n5514 & ~n6062 ) | ( n6061 & ~n6062 ) ;
  assign n6064 = n5994 ^ n5517 ^ x102 ;
  assign n6065 = n6006 ^ n5517 ^ 1'b0 ;
  assign n6066 = ( n5517 & n6064 ) | ( n5517 & ~n6065 ) | ( n6064 & ~n6065 ) ;
  assign n6067 = n5993 ^ n5520 ^ x101 ;
  assign n6068 = n6006 ^ n5520 ^ 1'b0 ;
  assign n6069 = ( n5520 & n6067 ) | ( n5520 & ~n6068 ) | ( n6067 & ~n6068 ) ;
  assign n6070 = n5990 ^ n5526 ^ x98 ;
  assign n6071 = n6006 ^ n5526 ^ 1'b0 ;
  assign n6072 = ( n5526 & n6070 ) | ( n5526 & ~n6071 ) | ( n6070 & ~n6071 ) ;
  assign n6073 = n5968 ^ n5443 ^ x90 ;
  assign n6074 = n6006 ^ n5443 ^ 1'b0 ;
  assign n6075 = ( n5443 & n6073 ) | ( n5443 & ~n6074 ) | ( n6073 & ~n6074 ) ;
  assign n6076 = n5966 ^ n5457 ^ x88 ;
  assign n6077 = n6006 ^ n5457 ^ 1'b0 ;
  assign n6078 = ( n5457 & n6076 ) | ( n5457 & ~n6077 ) | ( n6076 & ~n6077 ) ;
  assign n6079 = n5965 ^ n5460 ^ x87 ;
  assign n6080 = n6006 ^ n5460 ^ 1'b0 ;
  assign n6081 = ( n5460 & n6079 ) | ( n5460 & ~n6080 ) | ( n6079 & ~n6080 ) ;
  assign n6082 = n5953 ^ n5433 ^ x75 ;
  assign n6083 = n6006 ^ n5433 ^ 1'b0 ;
  assign n6084 = ( n5433 & n6082 ) | ( n5433 & ~n6083 ) | ( n6082 & ~n6083 ) ;
  assign n6085 = n5952 ^ n5481 ^ x74 ;
  assign n6086 = n6006 ^ n5481 ^ 1'b0 ;
  assign n6087 = ( n5481 & n6085 ) | ( n5481 & ~n6086 ) | ( n6085 & ~n6086 ) ;
  assign n6088 = n5951 ^ n5484 ^ x73 ;
  assign n6089 = n6006 ^ n5484 ^ 1'b0 ;
  assign n6090 = ( n5484 & n6088 ) | ( n5484 & ~n6089 ) | ( n6088 & ~n6089 ) ;
  assign n6091 = n5948 ^ n5490 ^ x70 ;
  assign n6092 = n6006 ^ n5490 ^ 1'b0 ;
  assign n6093 = ( n5490 & n6091 ) | ( n5490 & ~n6092 ) | ( n6091 & ~n6092 ) ;
  assign n6094 = n5947 ^ n5435 ^ x69 ;
  assign n6095 = n6006 ^ n5435 ^ 1'b0 ;
  assign n6096 = ( n5435 & n6094 ) | ( n5435 & ~n6095 ) | ( n6094 & ~n6095 ) ;
  assign n6097 = n5946 ^ n5493 ^ x68 ;
  assign n6098 = n6006 ^ n5493 ^ 1'b0 ;
  assign n6099 = ( n5493 & n6097 ) | ( n5493 & ~n6098 ) | ( n6097 & ~n6098 ) ;
  assign n6100 = n6003 ^ n5451 ^ x111 ;
  assign n6101 = n5967 ^ n5437 ^ x89 ;
  assign n6102 = x64 & n5806 ;
  assign n6103 = n5971 ^ n5440 ^ x93 ;
  assign n6104 = n5970 ^ n5454 ^ x92 ;
  assign n6105 = n5945 ^ n5412 ^ x67 ;
  assign n6106 = n5955 ^ n5419 ^ x77 ;
  assign n6107 = n6000 ^ n5502 ^ x108 ;
  assign n6108 = n5998 ^ n5442 ^ x106 ;
  assign n6109 = n5989 ^ n5431 ^ x97 ;
  assign n6110 = n5959 ^ n5472 ^ x81 ;
  assign n6111 = n6006 ^ n5440 ^ 1'b0 ;
  assign n6112 = ( n5440 & n6103 ) | ( n5440 & ~n6111 ) | ( n6103 & ~n6111 ) ;
  assign n6113 = n6006 ^ n5412 ^ 1'b0 ;
  assign n6114 = n6006 ^ n5454 ^ 1'b0 ;
  assign n6115 = ( n5454 & n6104 ) | ( n5454 & ~n6114 ) | ( n6104 & ~n6114 ) ;
  assign n6116 = n6006 ^ n5442 ^ 1'b0 ;
  assign n6117 = ( n5442 & n6108 ) | ( n5442 & ~n6116 ) | ( n6108 & ~n6116 ) ;
  assign n6118 = n6006 ^ n5451 ^ 1'b0 ;
  assign n6119 = n6006 ^ n5425 ^ 1'b0 ;
  assign n6120 = ( n5412 & n6105 ) | ( n5412 & ~n6113 ) | ( n6105 & ~n6113 ) ;
  assign n6121 = ( n5451 & n6100 ) | ( n5451 & ~n6118 ) | ( n6100 & ~n6118 ) ;
  assign n6122 = n6006 ^ n5508 ^ 1'b0 ;
  assign n6123 = n6006 ^ n5431 ^ 1'b0 ;
  assign n6124 = n6006 ^ n5502 ^ 1'b0 ;
  assign n6125 = n5997 ^ n5508 ^ x105 ;
  assign n6126 = n6102 ^ x64 ^ x14 ;
  assign n6127 = n6006 ^ n5472 ^ 1'b0 ;
  assign n6128 = ( n5431 & n6109 ) | ( n5431 & ~n6123 ) | ( n6109 & ~n6123 ) ;
  assign n6129 = ( n5508 & ~n6122 ) | ( n5508 & n6125 ) | ( ~n6122 & n6125 ) ;
  assign n6130 = ( n5472 & n6110 ) | ( n5472 & ~n6127 ) | ( n6110 & ~n6127 ) ;
  assign n6131 = n158 & n5447 ;
  assign n6132 = n6004 ^ n5447 ^ x112 ;
  assign n6133 = n6132 ^ n6006 ^ 1'b0 ;
  assign n6134 = ( n5447 & n6132 ) | ( n5447 & n6133 ) | ( n6132 & n6133 ) ;
  assign n6135 = n5969 ^ n5425 ^ x91 ;
  assign n6136 = ( n5502 & n6107 ) | ( n5502 & ~n6124 ) | ( n6107 & ~n6124 ) ;
  assign n6137 = n158 & n6134 ;
  assign n6138 = n6006 ^ n5437 ^ 1'b0 ;
  assign n6139 = ( n5437 & n6101 ) | ( n5437 & ~n6138 ) | ( n6101 & ~n6138 ) ;
  assign n6140 = n6006 ^ n5419 ^ 1'b0 ;
  assign n6141 = ( n5425 & ~n6119 ) | ( n5425 & n6135 ) | ( ~n6119 & n6135 ) ;
  assign n6142 = ( n5419 & n6106 ) | ( n5419 & ~n6140 ) | ( n6106 & ~n6140 ) ;
  assign n6143 = n6011 ^ n5732 ^ x65 ;
  assign n6144 = ( x65 & n5732 ) | ( x65 & n6143 ) | ( n5732 & n6143 ) ;
  assign n6145 = n6144 ^ n6040 ^ x66 ;
  assign n6146 = ( x66 & n6144 ) | ( x66 & n6145 ) | ( n6144 & n6145 ) ;
  assign n6147 = ( x67 & ~n6030 ) | ( x67 & n6146 ) | ( ~n6030 & n6146 ) ;
  assign n6148 = ( x68 & ~n6120 ) | ( x68 & n6147 ) | ( ~n6120 & n6147 ) ;
  assign n6149 = ( x69 & ~n6099 ) | ( x69 & n6148 ) | ( ~n6099 & n6148 ) ;
  assign n6150 = ( x70 & ~n6096 ) | ( x70 & n6149 ) | ( ~n6096 & n6149 ) ;
  assign n6151 = ( x71 & ~n6093 ) | ( x71 & n6150 ) | ( ~n6093 & n6150 ) ;
  assign n6152 = ( x72 & ~n6046 ) | ( x72 & n6151 ) | ( ~n6046 & n6151 ) ;
  assign n6153 = ( x73 & ~n6017 ) | ( x73 & n6152 ) | ( ~n6017 & n6152 ) ;
  assign n6154 = ( x74 & ~n6090 ) | ( x74 & n6153 ) | ( ~n6090 & n6153 ) ;
  assign n6155 = ( x75 & ~n6087 ) | ( x75 & n6154 ) | ( ~n6087 & n6154 ) ;
  assign n6156 = ( x76 & ~n6084 ) | ( x76 & n6155 ) | ( ~n6084 & n6155 ) ;
  assign n6157 = ( x77 & ~n6026 ) | ( x77 & n6156 ) | ( ~n6026 & n6156 ) ;
  assign n6158 = ( x78 & ~n6142 ) | ( x78 & n6157 ) | ( ~n6142 & n6157 ) ;
  assign n6159 = ( x79 & ~n6038 ) | ( x79 & n6158 ) | ( ~n6038 & n6158 ) ;
  assign n6160 = ( x80 & ~n6034 ) | ( x80 & n6159 ) | ( ~n6034 & n6159 ) ;
  assign n6161 = ( x81 & ~n6018 ) | ( x81 & n6160 ) | ( ~n6018 & n6160 ) ;
  assign n6162 = ( x82 & ~n6130 ) | ( x82 & n6161 ) | ( ~n6130 & n6161 ) ;
  assign n6163 = ( x83 & ~n6042 ) | ( x83 & n6162 ) | ( ~n6042 & n6162 ) ;
  assign n6164 = ( x84 & ~n6048 ) | ( x84 & n6163 ) | ( ~n6048 & n6163 ) ;
  assign n6165 = ( x85 & ~n6043 ) | ( x85 & n6164 ) | ( ~n6043 & n6164 ) ;
  assign n6166 = ( x86 & ~n6013 ) | ( x86 & n6165 ) | ( ~n6013 & n6165 ) ;
  assign n6167 = ( x87 & ~n6047 ) | ( x87 & n6166 ) | ( ~n6047 & n6166 ) ;
  assign n6168 = ( x88 & ~n6081 ) | ( x88 & n6167 ) | ( ~n6081 & n6167 ) ;
  assign n6169 = ( x89 & ~n6078 ) | ( x89 & n6168 ) | ( ~n6078 & n6168 ) ;
  assign n6170 = ( x90 & ~n6139 ) | ( x90 & n6169 ) | ( ~n6139 & n6169 ) ;
  assign n6171 = ( x91 & ~n6075 ) | ( x91 & n6170 ) | ( ~n6075 & n6170 ) ;
  assign n6172 = ( x92 & ~n6141 ) | ( x92 & n6171 ) | ( ~n6141 & n6171 ) ;
  assign n6173 = ( x93 & ~n6115 ) | ( x93 & n6172 ) | ( ~n6115 & n6172 ) ;
  assign n6174 = ( x94 & ~n6112 ) | ( x94 & n6173 ) | ( ~n6112 & n6173 ) ;
  assign n6175 = ( x95 & ~n6020 ) | ( x95 & n6174 ) | ( ~n6020 & n6174 ) ;
  assign n6176 = n6160 ^ n6018 ^ x81 ;
  assign n6177 = n6161 ^ n6130 ^ x82 ;
  assign n6178 = n6156 ^ n6026 ^ x77 ;
  assign n6179 = n6163 ^ n6048 ^ x84 ;
  assign n6180 = n6164 ^ n6043 ^ x85 ;
  assign n6181 = n6165 ^ n6013 ^ x86 ;
  assign n6182 = n6157 ^ n6142 ^ x78 ;
  assign n6183 = ( x96 & ~n6044 ) | ( x96 & n6175 ) | ( ~n6044 & n6175 ) ;
  assign n6184 = n6159 ^ n6034 ^ x80 ;
  assign n6185 = n6175 ^ n6044 ^ x96 ;
  assign n6186 = n6170 ^ n6075 ^ x91 ;
  assign n6187 = n6171 ^ n6141 ^ x92 ;
  assign n6188 = n6152 ^ n6017 ^ x73 ;
  assign n6189 = n6150 ^ n6093 ^ x71 ;
  assign n6190 = n6149 ^ n6096 ^ x70 ;
  assign n6191 = n6148 ^ n6099 ^ x69 ;
  assign n6192 = n6147 ^ n6120 ^ x68 ;
  assign n6193 = ( x97 & ~n6025 ) | ( x97 & n6183 ) | ( ~n6025 & n6183 ) ;
  assign n6194 = ( x98 & ~n6128 ) | ( x98 & n6193 ) | ( ~n6128 & n6193 ) ;
  assign n6195 = ( x99 & ~n6072 ) | ( x99 & n6194 ) | ( ~n6072 & n6194 ) ;
  assign n6196 = ( x100 & ~n6029 ) | ( x100 & n6195 ) | ( ~n6029 & n6195 ) ;
  assign n6197 = ( x101 & ~n6045 ) | ( x101 & n6196 ) | ( ~n6045 & n6196 ) ;
  assign n6198 = ( x102 & ~n6069 ) | ( x102 & n6197 ) | ( ~n6069 & n6197 ) ;
  assign n6199 = ( x103 & ~n6066 ) | ( x103 & n6198 ) | ( ~n6066 & n6198 ) ;
  assign n6200 = ( x104 & ~n6063 ) | ( x104 & n6199 ) | ( ~n6063 & n6199 ) ;
  assign n6201 = ( x105 & ~n6060 ) | ( x105 & n6200 ) | ( ~n6060 & n6200 ) ;
  assign n6202 = ( x106 & ~n6129 ) | ( x106 & n6201 ) | ( ~n6129 & n6201 ) ;
  assign n6203 = ( x107 & ~n6117 ) | ( x107 & n6202 ) | ( ~n6117 & n6202 ) ;
  assign n6204 = ( x108 & ~n6057 ) | ( x108 & n6203 ) | ( ~n6057 & n6203 ) ;
  assign n6205 = ( x109 & ~n6136 ) | ( x109 & n6204 ) | ( ~n6136 & n6204 ) ;
  assign n6206 = ( x110 & ~n6054 ) | ( x110 & n6205 ) | ( ~n6054 & n6205 ) ;
  assign n6207 = ( x111 & ~n6051 ) | ( x111 & n6206 ) | ( ~n6051 & n6206 ) ;
  assign n6208 = ( x112 & ~n6121 ) | ( x112 & n6207 ) | ( ~n6121 & n6207 ) ;
  assign n6209 = ( x113 & ~n6134 ) | ( x113 & n6208 ) | ( ~n6134 & n6208 ) ;
  assign n6210 = ( ~x113 & n5731 ) | ( ~x113 & n6134 ) | ( n5731 & n6134 ) ;
  assign n6211 = n6209 | n6210 ;
  assign n6212 = ( ~n6134 & n6137 ) | ( ~n6134 & n6211 ) | ( n6137 & n6211 ) ;
  assign n6213 = n6212 ^ n6044 ^ 1'b0 ;
  assign n6214 = ( n6044 & n6185 ) | ( n6044 & ~n6213 ) | ( n6185 & ~n6213 ) ;
  assign n6215 = n6212 ^ n6141 ^ 1'b0 ;
  assign n6216 = ( n6141 & n6187 ) | ( n6141 & ~n6215 ) | ( n6187 & ~n6215 ) ;
  assign n6217 = n6212 ^ n6075 ^ 1'b0 ;
  assign n6218 = ( n6075 & n6186 ) | ( n6075 & ~n6217 ) | ( n6186 & ~n6217 ) ;
  assign n6219 = n6212 ^ n6013 ^ 1'b0 ;
  assign n6220 = ( n6013 & n6181 ) | ( n6013 & ~n6219 ) | ( n6181 & ~n6219 ) ;
  assign n6221 = n6212 ^ n6043 ^ 1'b0 ;
  assign n6222 = ( n6043 & n6180 ) | ( n6043 & ~n6221 ) | ( n6180 & ~n6221 ) ;
  assign n6223 = n6212 ^ n6048 ^ 1'b0 ;
  assign n6224 = ( n6048 & n6179 ) | ( n6048 & ~n6223 ) | ( n6179 & ~n6223 ) ;
  assign n6225 = n6212 ^ n6130 ^ 1'b0 ;
  assign n6226 = ( n6130 & n6177 ) | ( n6130 & ~n6225 ) | ( n6177 & ~n6225 ) ;
  assign n6227 = n6212 ^ n6018 ^ 1'b0 ;
  assign n6228 = ( n6018 & n6176 ) | ( n6018 & ~n6227 ) | ( n6176 & ~n6227 ) ;
  assign n6229 = n6212 ^ n6034 ^ 1'b0 ;
  assign n6230 = ( n6034 & n6184 ) | ( n6034 & ~n6229 ) | ( n6184 & ~n6229 ) ;
  assign n6231 = n6212 ^ n6142 ^ 1'b0 ;
  assign n6232 = ( n6142 & n6182 ) | ( n6142 & ~n6231 ) | ( n6182 & ~n6231 ) ;
  assign n6233 = n6212 ^ n6026 ^ 1'b0 ;
  assign n6234 = ( n6026 & n6178 ) | ( n6026 & ~n6233 ) | ( n6178 & ~n6233 ) ;
  assign n6235 = n6212 ^ n6017 ^ 1'b0 ;
  assign n6236 = ( n6017 & n6188 ) | ( n6017 & ~n6235 ) | ( n6188 & ~n6235 ) ;
  assign n6237 = n6212 ^ n6093 ^ 1'b0 ;
  assign n6238 = ( n6093 & n6189 ) | ( n6093 & ~n6237 ) | ( n6189 & ~n6237 ) ;
  assign n6239 = n6212 ^ n6096 ^ 1'b0 ;
  assign n6240 = ( n6096 & n6190 ) | ( n6096 & ~n6239 ) | ( n6190 & ~n6239 ) ;
  assign n6241 = n6212 ^ n6099 ^ 1'b0 ;
  assign n6242 = ( n6099 & n6191 ) | ( n6099 & ~n6241 ) | ( n6191 & ~n6241 ) ;
  assign n6243 = n6212 ^ n6120 ^ 1'b0 ;
  assign n6244 = ( n6120 & n6192 ) | ( n6120 & ~n6243 ) | ( n6192 & ~n6243 ) ;
  assign n6245 = n6212 ^ n6145 ^ 1'b0 ;
  assign n6246 = ( n6040 & n6145 ) | ( n6040 & n6245 ) | ( n6145 & n6245 ) ;
  assign n6247 = n6212 ^ n6143 ^ 1'b0 ;
  assign n6248 = ( n6011 & n6143 ) | ( n6011 & n6247 ) | ( n6143 & n6247 ) ;
  assign n6249 = n6208 ^ n6134 ^ x113 ;
  assign n6250 = ~n6212 & n6249 ;
  assign n6251 = n6131 & ~n6211 ;
  assign n6252 = ( n6131 & n6250 ) | ( n6131 & ~n6251 ) | ( n6250 & ~n6251 ) ;
  assign n6253 = n6207 ^ n6121 ^ x112 ;
  assign n6254 = n6212 ^ n6121 ^ 1'b0 ;
  assign n6255 = ( n6121 & n6253 ) | ( n6121 & ~n6254 ) | ( n6253 & ~n6254 ) ;
  assign n6256 = n6206 ^ n6051 ^ x111 ;
  assign n6257 = n6212 ^ n6051 ^ 1'b0 ;
  assign n6258 = ( n6051 & n6256 ) | ( n6051 & ~n6257 ) | ( n6256 & ~n6257 ) ;
  assign n6259 = n6174 ^ n6020 ^ x95 ;
  assign n6260 = n6212 ^ n6020 ^ 1'b0 ;
  assign n6261 = ( n6020 & n6259 ) | ( n6020 & ~n6260 ) | ( n6259 & ~n6260 ) ;
  assign n6262 = n6173 ^ n6112 ^ x94 ;
  assign n6263 = n6212 ^ n6112 ^ 1'b0 ;
  assign n6264 = ( n6112 & n6262 ) | ( n6112 & ~n6263 ) | ( n6262 & ~n6263 ) ;
  assign n6265 = n6172 ^ n6115 ^ x93 ;
  assign n6266 = n6212 ^ n6115 ^ 1'b0 ;
  assign n6267 = ( n6115 & n6265 ) | ( n6115 & ~n6266 ) | ( n6265 & ~n6266 ) ;
  assign n6268 = n6169 ^ n6139 ^ x90 ;
  assign n6269 = n6212 ^ n6139 ^ 1'b0 ;
  assign n6270 = ( n6139 & n6268 ) | ( n6139 & ~n6269 ) | ( n6268 & ~n6269 ) ;
  assign n6271 = n6212 ^ n6078 ^ 1'b0 ;
  assign n6272 = n6167 ^ n6081 ^ x88 ;
  assign n6273 = n6212 ^ n6081 ^ 1'b0 ;
  assign n6274 = ( n6081 & n6272 ) | ( n6081 & ~n6273 ) | ( n6272 & ~n6273 ) ;
  assign n6275 = n6166 ^ n6047 ^ x87 ;
  assign n6276 = n6212 ^ n6047 ^ 1'b0 ;
  assign n6277 = n6168 ^ n6078 ^ x89 ;
  assign n6278 = ( n6078 & ~n6271 ) | ( n6078 & n6277 ) | ( ~n6271 & n6277 ) ;
  assign n6279 = ( n6047 & n6275 ) | ( n6047 & ~n6276 ) | ( n6275 & ~n6276 ) ;
  assign n6280 = n6162 ^ n6042 ^ x83 ;
  assign n6281 = n6212 ^ n6042 ^ 1'b0 ;
  assign n6282 = ( n6042 & n6280 ) | ( n6042 & ~n6281 ) | ( n6280 & ~n6281 ) ;
  assign n6283 = n6158 ^ n6038 ^ x79 ;
  assign n6284 = n6212 ^ n6038 ^ 1'b0 ;
  assign n6285 = ( n6038 & n6283 ) | ( n6038 & ~n6284 ) | ( n6283 & ~n6284 ) ;
  assign n6286 = n6155 ^ n6084 ^ x76 ;
  assign n6287 = n6212 ^ n6084 ^ 1'b0 ;
  assign n6288 = ( n6084 & n6286 ) | ( n6084 & ~n6287 ) | ( n6286 & ~n6287 ) ;
  assign n6289 = n6154 ^ n6087 ^ x75 ;
  assign n6290 = n6212 ^ n6087 ^ 1'b0 ;
  assign n6291 = ( n6087 & n6289 ) | ( n6087 & ~n6290 ) | ( n6289 & ~n6290 ) ;
  assign n6292 = n6153 ^ n6090 ^ x74 ;
  assign n6293 = n6212 ^ n6090 ^ 1'b0 ;
  assign n6294 = ( n6090 & n6292 ) | ( n6090 & ~n6293 ) | ( n6292 & ~n6293 ) ;
  assign n6295 = n6151 ^ n6046 ^ x72 ;
  assign n6296 = n6212 ^ n6046 ^ 1'b0 ;
  assign n6297 = ( n6046 & n6295 ) | ( n6046 & ~n6296 ) | ( n6295 & ~n6296 ) ;
  assign n6298 = n6146 ^ n6030 ^ x67 ;
  assign n6299 = n6212 ^ n6030 ^ 1'b0 ;
  assign n6300 = ( n6030 & n6298 ) | ( n6030 & ~n6299 ) | ( n6298 & ~n6299 ) ;
  assign n6301 = n6205 ^ n6054 ^ x110 ;
  assign n6302 = n6212 ^ n6054 ^ 1'b0 ;
  assign n6303 = ( n6054 & n6301 ) | ( n6054 & ~n6302 ) | ( n6301 & ~n6302 ) ;
  assign n6304 = n6204 ^ n6136 ^ x109 ;
  assign n6305 = n6212 ^ n6136 ^ 1'b0 ;
  assign n6306 = ( n6136 & n6304 ) | ( n6136 & ~n6305 ) | ( n6304 & ~n6305 ) ;
  assign n6307 = n6203 ^ n6057 ^ x108 ;
  assign n6308 = n6212 ^ n6057 ^ 1'b0 ;
  assign n6309 = ( n6057 & n6307 ) | ( n6057 & ~n6308 ) | ( n6307 & ~n6308 ) ;
  assign n6310 = n6202 ^ n6117 ^ x107 ;
  assign n6311 = n6212 ^ n6117 ^ 1'b0 ;
  assign n6312 = ( n6117 & n6310 ) | ( n6117 & ~n6311 ) | ( n6310 & ~n6311 ) ;
  assign n6313 = n6201 ^ n6129 ^ x106 ;
  assign n6314 = n6212 ^ n6129 ^ 1'b0 ;
  assign n6315 = ( n6129 & n6313 ) | ( n6129 & ~n6314 ) | ( n6313 & ~n6314 ) ;
  assign n6316 = n6200 ^ n6060 ^ x105 ;
  assign n6317 = n6212 ^ n6060 ^ 1'b0 ;
  assign n6318 = ( n6060 & n6316 ) | ( n6060 & ~n6317 ) | ( n6316 & ~n6317 ) ;
  assign n6319 = n6199 ^ n6063 ^ x104 ;
  assign n6320 = n6212 ^ n6063 ^ 1'b0 ;
  assign n6321 = ( n6063 & n6319 ) | ( n6063 & ~n6320 ) | ( n6319 & ~n6320 ) ;
  assign n6322 = n6198 ^ n6066 ^ x103 ;
  assign n6323 = n6212 ^ n6066 ^ 1'b0 ;
  assign n6324 = ( n6066 & n6322 ) | ( n6066 & ~n6323 ) | ( n6322 & ~n6323 ) ;
  assign n6325 = n6197 ^ n6069 ^ x102 ;
  assign n6326 = n6212 ^ n6069 ^ 1'b0 ;
  assign n6327 = ( n6069 & n6325 ) | ( n6069 & ~n6326 ) | ( n6325 & ~n6326 ) ;
  assign n6328 = n6196 ^ n6045 ^ x101 ;
  assign n6329 = n6212 ^ n6045 ^ 1'b0 ;
  assign n6330 = ( n6045 & n6328 ) | ( n6045 & ~n6329 ) | ( n6328 & ~n6329 ) ;
  assign n6331 = n6195 ^ n6029 ^ x100 ;
  assign n6332 = n6212 ^ n6029 ^ 1'b0 ;
  assign n6333 = ( n6029 & n6331 ) | ( n6029 & ~n6332 ) | ( n6331 & ~n6332 ) ;
  assign n6334 = n6194 ^ n6072 ^ x99 ;
  assign n6335 = n6212 ^ n6072 ^ 1'b0 ;
  assign n6336 = ( n6072 & n6334 ) | ( n6072 & ~n6335 ) | ( n6334 & ~n6335 ) ;
  assign n6337 = n6193 ^ n6128 ^ x98 ;
  assign n6338 = n6212 ^ n6128 ^ 1'b0 ;
  assign n6339 = ( n6128 & n6337 ) | ( n6128 & ~n6338 ) | ( n6337 & ~n6338 ) ;
  assign n6340 = n6183 ^ n6025 ^ x97 ;
  assign n6341 = n6212 ^ n6025 ^ 1'b0 ;
  assign n6342 = ( n6025 & n6340 ) | ( n6025 & ~n6341 ) | ( n6340 & ~n6341 ) ;
  assign n6343 = ~x13 & x64 ;
  assign n6344 = n6343 ^ n6126 ^ x65 ;
  assign n6345 = ( x65 & n6343 ) | ( x65 & n6344 ) | ( n6343 & n6344 ) ;
  assign n6346 = n6345 ^ n5842 ^ x66 ;
  assign n6347 = ( x66 & n6345 ) | ( x66 & n6346 ) | ( n6345 & n6346 ) ;
  assign n6348 = ( x67 & ~n5840 ) | ( x67 & n6347 ) | ( ~n5840 & n6347 ) ;
  assign n6349 = ( x68 & ~n5838 ) | ( x68 & n6348 ) | ( ~n5838 & n6348 ) ;
  assign n6350 = ( x69 & ~n5894 ) | ( x69 & n6349 ) | ( ~n5894 & n6349 ) ;
  assign n6351 = ( x70 & ~n5891 ) | ( x70 & n6350 ) | ( ~n5891 & n6350 ) ;
  assign n6352 = ( x71 & ~n5888 ) | ( x71 & n6351 ) | ( ~n5888 & n6351 ) ;
  assign n6353 = ( x72 & ~n5836 ) | ( x72 & n6352 ) | ( ~n5836 & n6352 ) ;
  assign n6354 = ( x73 & ~n5885 ) | ( x73 & n6353 ) | ( ~n5885 & n6353 ) ;
  assign n6355 = ( x74 & ~n5834 ) | ( x74 & n6354 ) | ( ~n5834 & n6354 ) ;
  assign n6356 = ( x75 & ~n5882 ) | ( x75 & n6355 ) | ( ~n5882 & n6355 ) ;
  assign n6357 = ( x76 & ~n5879 ) | ( x76 & n6356 ) | ( ~n5879 & n6356 ) ;
  assign n6358 = ( x77 & ~n5832 ) | ( x77 & n6357 ) | ( ~n5832 & n6357 ) ;
  assign n6359 = ( x78 & ~n5830 ) | ( x78 & n6358 ) | ( ~n5830 & n6358 ) ;
  assign n6360 = ( x79 & ~n5876 ) | ( x79 & n6359 ) | ( ~n5876 & n6359 ) ;
  assign n6361 = ( x80 & ~n5873 ) | ( x80 & n6360 ) | ( ~n5873 & n6360 ) ;
  assign n6362 = ( x81 & ~n5870 ) | ( x81 & n6361 ) | ( ~n5870 & n6361 ) ;
  assign n6363 = ( x82 & ~n5828 ) | ( x82 & n6362 ) | ( ~n5828 & n6362 ) ;
  assign n6364 = n322 | n5843 ;
  assign n6365 = ( x114 & n182 ) | ( x114 & ~n5843 ) | ( n182 & ~n5843 ) ;
  assign n6366 = ( x83 & ~n5826 ) | ( x83 & n6363 ) | ( ~n5826 & n6363 ) ;
  assign n6367 = ( x84 & ~n5867 ) | ( x84 & n6366 ) | ( ~n5867 & n6366 ) ;
  assign n6368 = ( x85 & ~n5864 ) | ( x85 & n6367 ) | ( ~n5864 & n6367 ) ;
  assign n6369 = ( x86 & ~n5861 ) | ( x86 & n6368 ) | ( ~n5861 & n6368 ) ;
  assign n6370 = ( x87 & ~n5858 ) | ( x87 & n6369 ) | ( ~n5858 & n6369 ) ;
  assign n6371 = ( x88 & ~n5824 ) | ( x88 & n6370 ) | ( ~n5824 & n6370 ) ;
  assign n6372 = ( x89 & ~n5855 ) | ( x89 & n6371 ) | ( ~n5855 & n6371 ) ;
  assign n6373 = ( x90 & ~n5852 ) | ( x90 & n6372 ) | ( ~n5852 & n6372 ) ;
  assign n6374 = ( x91 & ~n5939 ) | ( x91 & n6373 ) | ( ~n5939 & n6373 ) ;
  assign n6375 = n6359 ^ n5876 ^ x79 ;
  assign n6376 = n6360 ^ n5873 ^ x80 ;
  assign n6377 = ( x92 & ~n5936 ) | ( x92 & n6374 ) | ( ~n5936 & n6374 ) ;
  assign n6378 = n6362 ^ n5828 ^ x82 ;
  assign n6379 = n6367 ^ n5864 ^ x85 ;
  assign n6380 = n6366 ^ n5867 ^ x84 ;
  assign n6381 = n6369 ^ n5858 ^ x87 ;
  assign n6382 = ( x93 & ~n5933 ) | ( x93 & n6377 ) | ( ~n5933 & n6377 ) ;
  assign n6383 = ( x94 & ~n5930 ) | ( x94 & n6382 ) | ( ~n5930 & n6382 ) ;
  assign n6384 = n6370 ^ n5824 ^ x88 ;
  assign n6385 = n6371 ^ n5855 ^ x89 ;
  assign n6386 = n6372 ^ n5852 ^ x90 ;
  assign n6387 = n6352 ^ n5836 ^ x72 ;
  assign n6388 = n6383 ^ n5822 ^ x95 ;
  assign n6389 = n6353 ^ n5885 ^ x73 ;
  assign n6390 = n6382 ^ n5930 ^ x94 ;
  assign n6391 = ( x95 & ~n5822 ) | ( x95 & n6383 ) | ( ~n5822 & n6383 ) ;
  assign n6392 = ( x96 & ~n5927 ) | ( x96 & n6391 ) | ( ~n5927 & n6391 ) ;
  assign n6393 = n6349 ^ n5894 ^ x69 ;
  assign n6394 = ( x97 & ~n5820 ) | ( x97 & n6392 ) | ( ~n5820 & n6392 ) ;
  assign n6395 = ( x98 & ~n5924 ) | ( x98 & n6394 ) | ( ~n5924 & n6394 ) ;
  assign n6396 = ( x99 & ~n5921 ) | ( x99 & n6395 ) | ( ~n5921 & n6395 ) ;
  assign n6397 = ( x100 & ~n5918 ) | ( x100 & n6396 ) | ( ~n5918 & n6396 ) ;
  assign n6398 = ( x101 & ~n5815 ) | ( x101 & n6397 ) | ( ~n5815 & n6397 ) ;
  assign n6399 = ( x102 & ~n5915 ) | ( x102 & n6398 ) | ( ~n5915 & n6398 ) ;
  assign n6400 = ( x103 & ~n5912 ) | ( x103 & n6399 ) | ( ~n5912 & n6399 ) ;
  assign n6401 = ( x104 & ~n5909 ) | ( x104 & n6400 ) | ( ~n5909 & n6400 ) ;
  assign n6402 = ( x105 & ~n5906 ) | ( x105 & n6401 ) | ( ~n5906 & n6401 ) ;
  assign n6403 = ( x106 & ~n5903 ) | ( x106 & n6402 ) | ( ~n5903 & n6402 ) ;
  assign n6404 = ( x107 & ~n5900 ) | ( x107 & n6403 ) | ( ~n5900 & n6403 ) ;
  assign n6405 = ( x108 & ~n5897 ) | ( x108 & n6404 ) | ( ~n5897 & n6404 ) ;
  assign n6406 = ( x109 & ~n5849 ) | ( x109 & n6405 ) | ( ~n5849 & n6405 ) ;
  assign n6407 = ( x110 & ~n5812 ) | ( x110 & n6406 ) | ( ~n5812 & n6406 ) ;
  assign n6408 = ( x111 & ~n5809 ) | ( x111 & n6407 ) | ( ~n5809 & n6407 ) ;
  assign n6409 = ( x112 & ~n5846 ) | ( x112 & n6408 ) | ( ~n5846 & n6408 ) ;
  assign n6410 = ( x113 & ~n5817 ) | ( x113 & n6409 ) | ( ~n5817 & n6409 ) ;
  assign n6411 = ( ~x114 & n182 ) | ( ~x114 & n6364 ) | ( n182 & n6364 ) ;
  assign n6412 = ( n6365 & ~n6410 ) | ( n6365 & n6411 ) | ( ~n6410 & n6411 ) ;
  assign n6413 = n6410 | n6412 ;
  assign n6414 = n5731 & n6364 ;
  assign n6415 = ( ~n6364 & n6413 ) | ( ~n6364 & n6414 ) | ( n6413 & n6414 ) ;
  assign n6416 = n6400 ^ n5909 ^ x104 ;
  assign n6417 = n6415 ^ n5909 ^ 1'b0 ;
  assign n6418 = ( n5909 & n6416 ) | ( n5909 & ~n6417 ) | ( n6416 & ~n6417 ) ;
  assign n6419 = n6394 ^ n5924 ^ x98 ;
  assign n6420 = n6415 ^ n5924 ^ 1'b0 ;
  assign n6421 = ( n5924 & n6419 ) | ( n5924 & ~n6420 ) | ( n6419 & ~n6420 ) ;
  assign n6422 = n6415 ^ n5822 ^ 1'b0 ;
  assign n6423 = ( n5822 & n6388 ) | ( n5822 & ~n6422 ) | ( n6388 & ~n6422 ) ;
  assign n6424 = n6415 ^ n5930 ^ 1'b0 ;
  assign n6425 = ( n5930 & n6390 ) | ( n5930 & ~n6424 ) | ( n6390 & ~n6424 ) ;
  assign n6426 = n6415 ^ n5852 ^ 1'b0 ;
  assign n6427 = ( n5852 & n6386 ) | ( n5852 & ~n6426 ) | ( n6386 & ~n6426 ) ;
  assign n6428 = n6415 ^ n5855 ^ 1'b0 ;
  assign n6429 = ( n5855 & n6385 ) | ( n5855 & ~n6428 ) | ( n6385 & ~n6428 ) ;
  assign n6430 = n6415 ^ n5824 ^ 1'b0 ;
  assign n6431 = ( n5824 & n6384 ) | ( n5824 & ~n6430 ) | ( n6384 & ~n6430 ) ;
  assign n6432 = n6415 ^ n5858 ^ 1'b0 ;
  assign n6433 = ( n5858 & n6381 ) | ( n5858 & ~n6432 ) | ( n6381 & ~n6432 ) ;
  assign n6434 = n6415 ^ n5864 ^ 1'b0 ;
  assign n6435 = ( n5864 & n6379 ) | ( n5864 & ~n6434 ) | ( n6379 & ~n6434 ) ;
  assign n6436 = n6415 ^ n5867 ^ 1'b0 ;
  assign n6437 = ( n5867 & n6380 ) | ( n5867 & ~n6436 ) | ( n6380 & ~n6436 ) ;
  assign n6438 = n6415 ^ n5828 ^ 1'b0 ;
  assign n6439 = ( n5828 & n6378 ) | ( n5828 & ~n6438 ) | ( n6378 & ~n6438 ) ;
  assign n6440 = n6415 ^ n5873 ^ 1'b0 ;
  assign n6441 = ( n5873 & n6376 ) | ( n5873 & ~n6440 ) | ( n6376 & ~n6440 ) ;
  assign n6442 = n6415 ^ n5876 ^ 1'b0 ;
  assign n6443 = ( n5876 & n6375 ) | ( n5876 & ~n6442 ) | ( n6375 & ~n6442 ) ;
  assign n6444 = n6415 ^ n5885 ^ 1'b0 ;
  assign n6445 = ( n5885 & n6389 ) | ( n5885 & ~n6444 ) | ( n6389 & ~n6444 ) ;
  assign n6446 = n6415 ^ n5836 ^ 1'b0 ;
  assign n6447 = ( n5836 & n6387 ) | ( n5836 & ~n6446 ) | ( n6387 & ~n6446 ) ;
  assign n6448 = n6415 ^ n5894 ^ 1'b0 ;
  assign n6449 = ( n5894 & n6393 ) | ( n5894 & ~n6448 ) | ( n6393 & ~n6448 ) ;
  assign n6450 = n6415 ^ n6346 ^ 1'b0 ;
  assign n6451 = ( n5842 & n6346 ) | ( n5842 & n6450 ) | ( n6346 & n6450 ) ;
  assign n6452 = n6415 ^ n6344 ^ 1'b0 ;
  assign n6453 = ( n6126 & n6344 ) | ( n6126 & n6452 ) | ( n6344 & n6452 ) ;
  assign n6454 = ~n6413 & n6414 ;
  assign n6455 = ( n322 & n6414 ) | ( n322 & ~n6454 ) | ( n6414 & ~n6454 ) ;
  assign n6456 = n6409 ^ n5817 ^ x113 ;
  assign n6457 = n6415 ^ n5817 ^ 1'b0 ;
  assign n6458 = ( n5817 & n6456 ) | ( n5817 & ~n6457 ) | ( n6456 & ~n6457 ) ;
  assign n6459 = n6408 ^ n5846 ^ x112 ;
  assign n6460 = n6415 ^ n5846 ^ 1'b0 ;
  assign n6461 = ( n5846 & n6459 ) | ( n5846 & ~n6460 ) | ( n6459 & ~n6460 ) ;
  assign n6462 = n6407 ^ n5809 ^ x111 ;
  assign n6463 = n6415 ^ n5809 ^ 1'b0 ;
  assign n6464 = ( n5809 & n6462 ) | ( n5809 & ~n6463 ) | ( n6462 & ~n6463 ) ;
  assign n6465 = n6374 ^ n5936 ^ x92 ;
  assign n6466 = n6415 ^ n5936 ^ 1'b0 ;
  assign n6467 = ( n5936 & n6465 ) | ( n5936 & ~n6466 ) | ( n6465 & ~n6466 ) ;
  assign n6468 = n6373 ^ n5939 ^ x91 ;
  assign n6469 = n6415 ^ n5939 ^ 1'b0 ;
  assign n6470 = ( n5939 & n6468 ) | ( n5939 & ~n6469 ) | ( n6468 & ~n6469 ) ;
  assign n6471 = n6368 ^ n5861 ^ x86 ;
  assign n6472 = n6415 ^ n5861 ^ 1'b0 ;
  assign n6473 = ( n5861 & n6471 ) | ( n5861 & ~n6472 ) | ( n6471 & ~n6472 ) ;
  assign n6474 = n6363 ^ n5826 ^ x83 ;
  assign n6475 = n6415 ^ n5826 ^ 1'b0 ;
  assign n6476 = ( n5826 & n6474 ) | ( n5826 & ~n6475 ) | ( n6474 & ~n6475 ) ;
  assign n6477 = n6361 ^ n5870 ^ x81 ;
  assign n6478 = n6415 ^ n5870 ^ 1'b0 ;
  assign n6479 = ( n5870 & n6477 ) | ( n5870 & ~n6478 ) | ( n6477 & ~n6478 ) ;
  assign n6480 = n6358 ^ n5830 ^ x78 ;
  assign n6481 = n6415 ^ n5830 ^ 1'b0 ;
  assign n6482 = ( n5830 & n6480 ) | ( n5830 & ~n6481 ) | ( n6480 & ~n6481 ) ;
  assign n6483 = n6357 ^ n5832 ^ x77 ;
  assign n6484 = n6415 ^ n5832 ^ 1'b0 ;
  assign n6485 = ( n5832 & n6483 ) | ( n5832 & ~n6484 ) | ( n6483 & ~n6484 ) ;
  assign n6486 = n6356 ^ n5879 ^ x76 ;
  assign n6487 = n6415 ^ n5879 ^ 1'b0 ;
  assign n6488 = ( n5879 & n6486 ) | ( n5879 & ~n6487 ) | ( n6486 & ~n6487 ) ;
  assign n6489 = n6355 ^ n5882 ^ x75 ;
  assign n6490 = n6415 ^ n5882 ^ 1'b0 ;
  assign n6491 = ( n5882 & n6489 ) | ( n5882 & ~n6490 ) | ( n6489 & ~n6490 ) ;
  assign n6492 = n6354 ^ n5834 ^ x74 ;
  assign n6493 = n6415 ^ n5834 ^ 1'b0 ;
  assign n6494 = ( n5834 & n6492 ) | ( n5834 & ~n6493 ) | ( n6492 & ~n6493 ) ;
  assign n6495 = n6351 ^ n5888 ^ x71 ;
  assign n6496 = n6415 ^ n5888 ^ 1'b0 ;
  assign n6497 = ( n5888 & n6495 ) | ( n5888 & ~n6496 ) | ( n6495 & ~n6496 ) ;
  assign n6498 = n6350 ^ n5891 ^ x70 ;
  assign n6499 = n6415 ^ n5891 ^ 1'b0 ;
  assign n6500 = ( n5891 & n6498 ) | ( n5891 & ~n6499 ) | ( n6498 & ~n6499 ) ;
  assign n6501 = n6348 ^ n5838 ^ x68 ;
  assign n6502 = n6415 ^ n5838 ^ 1'b0 ;
  assign n6503 = ( n5838 & n6501 ) | ( n5838 & ~n6502 ) | ( n6501 & ~n6502 ) ;
  assign n6504 = n6347 ^ n5840 ^ x67 ;
  assign n6505 = n6415 ^ n5840 ^ 1'b0 ;
  assign n6506 = ( n5840 & n6504 ) | ( n5840 & ~n6505 ) | ( n6504 & ~n6505 ) ;
  assign n6507 = n6406 ^ n5812 ^ x110 ;
  assign n6508 = n6415 ^ n5812 ^ 1'b0 ;
  assign n6509 = ( n5812 & n6507 ) | ( n5812 & ~n6508 ) | ( n6507 & ~n6508 ) ;
  assign n6510 = n6405 ^ n5849 ^ x109 ;
  assign n6511 = n6415 ^ n5849 ^ 1'b0 ;
  assign n6512 = ( n5849 & n6510 ) | ( n5849 & ~n6511 ) | ( n6510 & ~n6511 ) ;
  assign n6513 = n6404 ^ n5897 ^ x108 ;
  assign n6514 = n6415 ^ n5897 ^ 1'b0 ;
  assign n6515 = ( n5897 & n6513 ) | ( n5897 & ~n6514 ) | ( n6513 & ~n6514 ) ;
  assign n6516 = n6403 ^ n5900 ^ x107 ;
  assign n6517 = n6415 ^ n5900 ^ 1'b0 ;
  assign n6518 = ( n5900 & n6516 ) | ( n5900 & ~n6517 ) | ( n6516 & ~n6517 ) ;
  assign n6519 = n6402 ^ n5903 ^ x106 ;
  assign n6520 = n6415 ^ n5903 ^ 1'b0 ;
  assign n6521 = ( n5903 & n6519 ) | ( n5903 & ~n6520 ) | ( n6519 & ~n6520 ) ;
  assign n6522 = n6401 ^ n5906 ^ x105 ;
  assign n6523 = n6415 ^ n5906 ^ 1'b0 ;
  assign n6524 = ( n5906 & n6522 ) | ( n5906 & ~n6523 ) | ( n6522 & ~n6523 ) ;
  assign n6525 = n6399 ^ n5912 ^ x103 ;
  assign n6526 = n6415 ^ n5912 ^ 1'b0 ;
  assign n6527 = ( n5912 & n6525 ) | ( n5912 & ~n6526 ) | ( n6525 & ~n6526 ) ;
  assign n6528 = n6398 ^ n5915 ^ x102 ;
  assign n6529 = n6415 ^ n5915 ^ 1'b0 ;
  assign n6530 = ( n5915 & n6528 ) | ( n5915 & ~n6529 ) | ( n6528 & ~n6529 ) ;
  assign n6531 = n6397 ^ n5815 ^ x101 ;
  assign n6532 = n6415 ^ n5815 ^ 1'b0 ;
  assign n6533 = ( n5815 & n6531 ) | ( n5815 & ~n6532 ) | ( n6531 & ~n6532 ) ;
  assign n6534 = n6396 ^ n5918 ^ x100 ;
  assign n6535 = n6415 ^ n5918 ^ 1'b0 ;
  assign n6536 = ( n5918 & n6534 ) | ( n5918 & ~n6535 ) | ( n6534 & ~n6535 ) ;
  assign n6537 = n6395 ^ n5921 ^ x99 ;
  assign n6538 = n6415 ^ n5921 ^ 1'b0 ;
  assign n6539 = ( n5921 & n6537 ) | ( n5921 & ~n6538 ) | ( n6537 & ~n6538 ) ;
  assign n6540 = n6392 ^ n5820 ^ x97 ;
  assign n6541 = n6415 ^ n5820 ^ 1'b0 ;
  assign n6542 = ( n5820 & n6540 ) | ( n5820 & ~n6541 ) | ( n6540 & ~n6541 ) ;
  assign n6543 = n6391 ^ n5927 ^ x96 ;
  assign n6544 = n6415 ^ n5927 ^ 1'b0 ;
  assign n6545 = ( n5927 & n6543 ) | ( n5927 & ~n6544 ) | ( n6543 & ~n6544 ) ;
  assign n6546 = n6377 ^ n5933 ^ x93 ;
  assign n6547 = n6415 ^ n5933 ^ 1'b0 ;
  assign n6548 = ( n5933 & n6546 ) | ( n5933 & ~n6547 ) | ( n6546 & ~n6547 ) ;
  assign n6549 = x64 & n6212 ;
  assign n6550 = n6549 ^ x64 ^ x14 ;
  assign n6551 = n6550 ^ n6343 ^ x65 ;
  assign n6552 = ( x65 & n6343 ) | ( x65 & n6551 ) | ( n6343 & n6551 ) ;
  assign n6553 = n6552 ^ n6248 ^ x66 ;
  assign n6554 = ( x66 & n6552 ) | ( x66 & n6553 ) | ( n6552 & n6553 ) ;
  assign n6555 = ( x67 & ~n6246 ) | ( x67 & n6554 ) | ( ~n6246 & n6554 ) ;
  assign n6556 = ( x68 & ~n6300 ) | ( x68 & n6555 ) | ( ~n6300 & n6555 ) ;
  assign n6557 = ( x69 & ~n6244 ) | ( x69 & n6556 ) | ( ~n6244 & n6556 ) ;
  assign n6558 = ( x70 & ~n6242 ) | ( x70 & n6557 ) | ( ~n6242 & n6557 ) ;
  assign n6559 = ( x71 & ~n6240 ) | ( x71 & n6558 ) | ( ~n6240 & n6558 ) ;
  assign n6560 = ( x72 & ~n6238 ) | ( x72 & n6559 ) | ( ~n6238 & n6559 ) ;
  assign n6561 = ( x73 & ~n6297 ) | ( x73 & n6560 ) | ( ~n6297 & n6560 ) ;
  assign n6562 = ( x74 & ~n6236 ) | ( x74 & n6561 ) | ( ~n6236 & n6561 ) ;
  assign n6563 = ( x75 & ~n6294 ) | ( x75 & n6562 ) | ( ~n6294 & n6562 ) ;
  assign n6564 = ( x76 & ~n6291 ) | ( x76 & n6563 ) | ( ~n6291 & n6563 ) ;
  assign n6565 = ( x77 & ~n6288 ) | ( x77 & n6564 ) | ( ~n6288 & n6564 ) ;
  assign n6566 = n6558 ^ n6240 ^ x71 ;
  assign n6567 = ( x78 & ~n6234 ) | ( x78 & n6565 ) | ( ~n6234 & n6565 ) ;
  assign n6568 = ( x79 & ~n6232 ) | ( x79 & n6567 ) | ( ~n6232 & n6567 ) ;
  assign n6569 = ( x80 & ~n6285 ) | ( x80 & n6568 ) | ( ~n6285 & n6568 ) ;
  assign n6570 = ( x81 & ~n6230 ) | ( x81 & n6569 ) | ( ~n6230 & n6569 ) ;
  assign n6571 = ( x82 & ~n6228 ) | ( x82 & n6570 ) | ( ~n6228 & n6570 ) ;
  assign n6572 = ( x83 & ~n6226 ) | ( x83 & n6571 ) | ( ~n6226 & n6571 ) ;
  assign n6573 = ( x84 & ~n6282 ) | ( x84 & n6572 ) | ( ~n6282 & n6572 ) ;
  assign n6574 = ( x85 & ~n6224 ) | ( x85 & n6573 ) | ( ~n6224 & n6573 ) ;
  assign n6575 = ( x86 & ~n6222 ) | ( x86 & n6574 ) | ( ~n6222 & n6574 ) ;
  assign n6576 = ( x87 & ~n6220 ) | ( x87 & n6575 ) | ( ~n6220 & n6575 ) ;
  assign n6577 = ( x88 & ~n6279 ) | ( x88 & n6576 ) | ( ~n6279 & n6576 ) ;
  assign n6578 = ( x89 & ~n6274 ) | ( x89 & n6577 ) | ( ~n6274 & n6577 ) ;
  assign n6579 = n6567 ^ n6232 ^ x79 ;
  assign n6580 = n6563 ^ n6291 ^ x76 ;
  assign n6581 = n6559 ^ n6238 ^ x72 ;
  assign n6582 = n6565 ^ n6234 ^ x78 ;
  assign n6583 = ( x90 & ~n6278 ) | ( x90 & n6578 ) | ( ~n6278 & n6578 ) ;
  assign n6584 = n6568 ^ n6285 ^ x80 ;
  assign n6585 = n6569 ^ n6230 ^ x81 ;
  assign n6586 = ( x91 & ~n6270 ) | ( x91 & n6583 ) | ( ~n6270 & n6583 ) ;
  assign n6587 = ( x92 & ~n6218 ) | ( x92 & n6586 ) | ( ~n6218 & n6586 ) ;
  assign n6588 = n6572 ^ n6282 ^ x84 ;
  assign n6589 = n6573 ^ n6224 ^ x85 ;
  assign n6590 = ( x93 & ~n6216 ) | ( x93 & n6587 ) | ( ~n6216 & n6587 ) ;
  assign n6591 = n6575 ^ n6220 ^ x87 ;
  assign n6592 = n6576 ^ n6279 ^ x88 ;
  assign n6593 = n6577 ^ n6274 ^ x89 ;
  assign n6594 = n6578 ^ n6278 ^ x90 ;
  assign n6595 = n6555 ^ n6300 ^ x68 ;
  assign n6596 = n5731 & n6252 ;
  assign n6597 = ( ~x114 & n182 ) | ( ~x114 & n6252 ) | ( n182 & n6252 ) ;
  assign n6598 = ( x94 & ~n6267 ) | ( x94 & n6590 ) | ( ~n6267 & n6590 ) ;
  assign n6599 = n6554 ^ n6246 ^ x67 ;
  assign n6600 = ( x95 & ~n6264 ) | ( x95 & n6598 ) | ( ~n6264 & n6598 ) ;
  assign n6601 = ( x96 & ~n6261 ) | ( x96 & n6600 ) | ( ~n6261 & n6600 ) ;
  assign n6602 = ( x97 & ~n6214 ) | ( x97 & n6601 ) | ( ~n6214 & n6601 ) ;
  assign n6603 = ( x98 & ~n6342 ) | ( x98 & n6602 ) | ( ~n6342 & n6602 ) ;
  assign n6604 = ( x99 & ~n6339 ) | ( x99 & n6603 ) | ( ~n6339 & n6603 ) ;
  assign n6605 = ( x100 & ~n6336 ) | ( x100 & n6604 ) | ( ~n6336 & n6604 ) ;
  assign n6606 = ( x101 & ~n6333 ) | ( x101 & n6605 ) | ( ~n6333 & n6605 ) ;
  assign n6607 = ( x102 & ~n6330 ) | ( x102 & n6606 ) | ( ~n6330 & n6606 ) ;
  assign n6608 = ( x103 & ~n6327 ) | ( x103 & n6607 ) | ( ~n6327 & n6607 ) ;
  assign n6609 = ( x104 & ~n6324 ) | ( x104 & n6608 ) | ( ~n6324 & n6608 ) ;
  assign n6610 = ( x105 & ~n6321 ) | ( x105 & n6609 ) | ( ~n6321 & n6609 ) ;
  assign n6611 = ( x106 & ~n6318 ) | ( x106 & n6610 ) | ( ~n6318 & n6610 ) ;
  assign n6612 = ( x107 & ~n6315 ) | ( x107 & n6611 ) | ( ~n6315 & n6611 ) ;
  assign n6613 = ( x108 & ~n6312 ) | ( x108 & n6612 ) | ( ~n6312 & n6612 ) ;
  assign n6614 = ( x109 & ~n6309 ) | ( x109 & n6613 ) | ( ~n6309 & n6613 ) ;
  assign n6615 = ( x110 & ~n6306 ) | ( x110 & n6614 ) | ( ~n6306 & n6614 ) ;
  assign n6616 = ( x111 & ~n6303 ) | ( x111 & n6615 ) | ( ~n6303 & n6615 ) ;
  assign n6617 = ( x112 & ~n6258 ) | ( x112 & n6616 ) | ( ~n6258 & n6616 ) ;
  assign n6618 = ( x113 & ~n6255 ) | ( x113 & n6617 ) | ( ~n6255 & n6617 ) ;
  assign n6619 = ( x114 & ~n6252 ) | ( x114 & n6618 ) | ( ~n6252 & n6618 ) ;
  assign n6620 = n6597 | n6619 ;
  assign n6621 = ( ~n6252 & n6596 ) | ( ~n6252 & n6620 ) | ( n6596 & n6620 ) ;
  assign n6622 = n6618 ^ n6252 ^ x114 ;
  assign n6623 = n6621 ^ n6230 ^ 1'b0 ;
  assign n6624 = ( n6230 & n6585 ) | ( n6230 & ~n6623 ) | ( n6585 & ~n6623 ) ;
  assign n6625 = n6621 ^ n6291 ^ 1'b0 ;
  assign n6626 = ( n6291 & n6580 ) | ( n6291 & ~n6625 ) | ( n6580 & ~n6625 ) ;
  assign n6627 = n6621 ^ n6279 ^ 1'b0 ;
  assign n6628 = n6621 ^ n6300 ^ 1'b0 ;
  assign n6629 = ( n6300 & n6595 ) | ( n6300 & ~n6628 ) | ( n6595 & ~n6628 ) ;
  assign n6630 = n6621 ^ n6278 ^ 1'b0 ;
  assign n6631 = n6621 ^ n6238 ^ 1'b0 ;
  assign n6632 = ( n6238 & n6581 ) | ( n6238 & ~n6631 ) | ( n6581 & ~n6631 ) ;
  assign n6633 = ( n6278 & n6594 ) | ( n6278 & ~n6630 ) | ( n6594 & ~n6630 ) ;
  assign n6634 = n6621 ^ n6551 ^ 1'b0 ;
  assign n6635 = ~n6621 & n6622 ;
  assign n6636 = ( n6550 & n6551 ) | ( n6550 & n6634 ) | ( n6551 & n6634 ) ;
  assign n6637 = n6621 ^ n6285 ^ 1'b0 ;
  assign n6638 = n6621 ^ n6267 ^ 1'b0 ;
  assign n6639 = n6621 ^ n6224 ^ 1'b0 ;
  assign n6640 = ( n6224 & n6589 ) | ( n6224 & ~n6639 ) | ( n6589 & ~n6639 ) ;
  assign n6641 = n6621 ^ n6240 ^ 1'b0 ;
  assign n6642 = ( n6240 & n6566 ) | ( n6240 & ~n6641 ) | ( n6566 & ~n6641 ) ;
  assign n6643 = n6621 ^ n6234 ^ 1'b0 ;
  assign n6644 = n6596 & ~n6620 ;
  assign n6645 = ( n6234 & n6582 ) | ( n6234 & ~n6643 ) | ( n6582 & ~n6643 ) ;
  assign n6646 = ( n6596 & n6635 ) | ( n6596 & ~n6644 ) | ( n6635 & ~n6644 ) ;
  assign n6647 = n6621 ^ n6274 ^ 1'b0 ;
  assign n6648 = n6590 ^ n6267 ^ x94 ;
  assign n6649 = ( n6274 & n6593 ) | ( n6274 & ~n6647 ) | ( n6593 & ~n6647 ) ;
  assign n6650 = n6621 ^ n6246 ^ 1'b0 ;
  assign n6651 = n6621 ^ n6220 ^ 1'b0 ;
  assign n6652 = ( n6246 & n6599 ) | ( n6246 & ~n6650 ) | ( n6599 & ~n6650 ) ;
  assign n6653 = n6621 ^ n6232 ^ 1'b0 ;
  assign n6654 = ( n6285 & n6584 ) | ( n6285 & ~n6637 ) | ( n6584 & ~n6637 ) ;
  assign n6655 = n6621 ^ n6282 ^ 1'b0 ;
  assign n6656 = ( n6220 & n6591 ) | ( n6220 & ~n6651 ) | ( n6591 & ~n6651 ) ;
  assign n6657 = ( n6279 & n6592 ) | ( n6279 & ~n6627 ) | ( n6592 & ~n6627 ) ;
  assign n6658 = ( n6282 & n6588 ) | ( n6282 & ~n6655 ) | ( n6588 & ~n6655 ) ;
  assign n6659 = ( n6232 & n6579 ) | ( n6232 & ~n6653 ) | ( n6579 & ~n6653 ) ;
  assign n6660 = ( n6267 & ~n6638 ) | ( n6267 & n6648 ) | ( ~n6638 & n6648 ) ;
  assign n6661 = n6617 ^ n6255 ^ x113 ;
  assign n6662 = n6621 ^ n6255 ^ 1'b0 ;
  assign n6663 = ( n6255 & n6661 ) | ( n6255 & ~n6662 ) | ( n6661 & ~n6662 ) ;
  assign n6664 = n6616 ^ n6258 ^ x112 ;
  assign n6665 = n6621 ^ n6258 ^ 1'b0 ;
  assign n6666 = ( n6258 & n6664 ) | ( n6258 & ~n6665 ) | ( n6664 & ~n6665 ) ;
  assign n6667 = n6601 ^ n6214 ^ x97 ;
  assign n6668 = n6621 ^ n6214 ^ 1'b0 ;
  assign n6669 = ( n6214 & n6667 ) | ( n6214 & ~n6668 ) | ( n6667 & ~n6668 ) ;
  assign n6670 = n6600 ^ n6261 ^ x96 ;
  assign n6671 = n6621 ^ n6261 ^ 1'b0 ;
  assign n6672 = ( n6261 & n6670 ) | ( n6261 & ~n6671 ) | ( n6670 & ~n6671 ) ;
  assign n6673 = n6598 ^ n6264 ^ x95 ;
  assign n6674 = n6621 ^ n6264 ^ 1'b0 ;
  assign n6675 = ( n6264 & n6673 ) | ( n6264 & ~n6674 ) | ( n6673 & ~n6674 ) ;
  assign n6676 = n6587 ^ n6216 ^ x93 ;
  assign n6677 = n6621 ^ n6216 ^ 1'b0 ;
  assign n6678 = ( n6216 & n6676 ) | ( n6216 & ~n6677 ) | ( n6676 & ~n6677 ) ;
  assign n6679 = n6586 ^ n6218 ^ x92 ;
  assign n6680 = n6621 ^ n6218 ^ 1'b0 ;
  assign n6681 = ( n6218 & n6679 ) | ( n6218 & ~n6680 ) | ( n6679 & ~n6680 ) ;
  assign n6682 = n6583 ^ n6270 ^ x91 ;
  assign n6683 = n6621 ^ n6270 ^ 1'b0 ;
  assign n6684 = ( n6270 & n6682 ) | ( n6270 & ~n6683 ) | ( n6682 & ~n6683 ) ;
  assign n6685 = n6574 ^ n6222 ^ x86 ;
  assign n6686 = n6621 ^ n6222 ^ 1'b0 ;
  assign n6687 = ( n6222 & n6685 ) | ( n6222 & ~n6686 ) | ( n6685 & ~n6686 ) ;
  assign n6688 = n6571 ^ n6226 ^ x83 ;
  assign n6689 = n6621 ^ n6226 ^ 1'b0 ;
  assign n6690 = ( n6226 & n6688 ) | ( n6226 & ~n6689 ) | ( n6688 & ~n6689 ) ;
  assign n6691 = n6570 ^ n6228 ^ x82 ;
  assign n6692 = n6621 ^ n6228 ^ 1'b0 ;
  assign n6693 = ( n6228 & n6691 ) | ( n6228 & ~n6692 ) | ( n6691 & ~n6692 ) ;
  assign n6694 = n6564 ^ n6288 ^ x77 ;
  assign n6695 = n6621 ^ n6288 ^ 1'b0 ;
  assign n6696 = ( n6288 & n6694 ) | ( n6288 & ~n6695 ) | ( n6694 & ~n6695 ) ;
  assign n6697 = n6562 ^ n6294 ^ x75 ;
  assign n6698 = n6621 ^ n6294 ^ 1'b0 ;
  assign n6699 = ( n6294 & n6697 ) | ( n6294 & ~n6698 ) | ( n6697 & ~n6698 ) ;
  assign n6700 = n6561 ^ n6236 ^ x74 ;
  assign n6701 = n6621 ^ n6236 ^ 1'b0 ;
  assign n6702 = ( n6236 & n6700 ) | ( n6236 & ~n6701 ) | ( n6700 & ~n6701 ) ;
  assign n6703 = n6560 ^ n6297 ^ x73 ;
  assign n6704 = n6621 ^ n6297 ^ 1'b0 ;
  assign n6705 = ( n6297 & n6703 ) | ( n6297 & ~n6704 ) | ( n6703 & ~n6704 ) ;
  assign n6706 = n6557 ^ n6242 ^ x70 ;
  assign n6707 = n6621 ^ n6242 ^ 1'b0 ;
  assign n6708 = ( n6242 & n6706 ) | ( n6242 & ~n6707 ) | ( n6706 & ~n6707 ) ;
  assign n6709 = n6556 ^ n6244 ^ x69 ;
  assign n6710 = n6621 ^ n6244 ^ 1'b0 ;
  assign n6711 = ( n6244 & n6709 ) | ( n6244 & ~n6710 ) | ( n6709 & ~n6710 ) ;
  assign n6712 = n6615 ^ n6303 ^ x111 ;
  assign n6713 = n6621 ^ n6303 ^ 1'b0 ;
  assign n6714 = ( n6303 & n6712 ) | ( n6303 & ~n6713 ) | ( n6712 & ~n6713 ) ;
  assign n6715 = n6614 ^ n6306 ^ x110 ;
  assign n6716 = n6613 ^ n6309 ^ x109 ;
  assign n6717 = n6621 ^ n6309 ^ 1'b0 ;
  assign n6718 = ( n6309 & n6716 ) | ( n6309 & ~n6717 ) | ( n6716 & ~n6717 ) ;
  assign n6719 = n6612 ^ n6312 ^ x108 ;
  assign n6720 = n6621 ^ n6312 ^ 1'b0 ;
  assign n6721 = ( n6312 & n6719 ) | ( n6312 & ~n6720 ) | ( n6719 & ~n6720 ) ;
  assign n6722 = n6611 ^ n6315 ^ x107 ;
  assign n6723 = n6621 ^ n6315 ^ 1'b0 ;
  assign n6724 = ( n6315 & n6722 ) | ( n6315 & ~n6723 ) | ( n6722 & ~n6723 ) ;
  assign n6725 = n6610 ^ n6318 ^ x106 ;
  assign n6726 = n6621 ^ n6318 ^ 1'b0 ;
  assign n6727 = n6609 ^ n6321 ^ x105 ;
  assign n6728 = n6621 ^ n6321 ^ 1'b0 ;
  assign n6729 = ( n6321 & n6727 ) | ( n6321 & ~n6728 ) | ( n6727 & ~n6728 ) ;
  assign n6730 = n6608 ^ n6324 ^ x104 ;
  assign n6731 = n6621 ^ n6324 ^ 1'b0 ;
  assign n6732 = ( n6324 & n6730 ) | ( n6324 & ~n6731 ) | ( n6730 & ~n6731 ) ;
  assign n6733 = n6607 ^ n6327 ^ x103 ;
  assign n6734 = n6621 ^ n6306 ^ 1'b0 ;
  assign n6735 = ( n6306 & n6715 ) | ( n6306 & ~n6734 ) | ( n6715 & ~n6734 ) ;
  assign n6736 = n6621 ^ n6327 ^ 1'b0 ;
  assign n6737 = ( n6327 & n6733 ) | ( n6327 & ~n6736 ) | ( n6733 & ~n6736 ) ;
  assign n6738 = n6606 ^ n6330 ^ x102 ;
  assign n6739 = n6621 ^ n6330 ^ 1'b0 ;
  assign n6740 = ( n6330 & n6738 ) | ( n6330 & ~n6739 ) | ( n6738 & ~n6739 ) ;
  assign n6741 = n6605 ^ n6333 ^ x101 ;
  assign n6742 = n6621 ^ n6333 ^ 1'b0 ;
  assign n6743 = ( n6333 & n6741 ) | ( n6333 & ~n6742 ) | ( n6741 & ~n6742 ) ;
  assign n6744 = n6604 ^ n6336 ^ x100 ;
  assign n6745 = n6621 ^ n6336 ^ 1'b0 ;
  assign n6746 = ( n6336 & n6744 ) | ( n6336 & ~n6745 ) | ( n6744 & ~n6745 ) ;
  assign n6747 = n6603 ^ n6339 ^ x99 ;
  assign n6748 = n6621 ^ n6339 ^ 1'b0 ;
  assign n6749 = ( n6339 & n6747 ) | ( n6339 & ~n6748 ) | ( n6747 & ~n6748 ) ;
  assign n6750 = n6602 ^ n6342 ^ x98 ;
  assign n6751 = n6621 ^ n6342 ^ 1'b0 ;
  assign n6752 = ( n6342 & n6750 ) | ( n6342 & ~n6751 ) | ( n6750 & ~n6751 ) ;
  assign n6753 = ( n6318 & n6725 ) | ( n6318 & ~n6726 ) | ( n6725 & ~n6726 ) ;
  assign n6754 = n6621 ^ n6553 ^ 1'b0 ;
  assign n6755 = ( n6248 & n6553 ) | ( n6248 & n6754 ) | ( n6553 & n6754 ) ;
  assign n6756 = x64 & n6621 ;
  assign n6757 = ~x12 & x64 ;
  assign n6758 = n6756 ^ x64 ^ x13 ;
  assign n6759 = n6758 ^ n6757 ^ x65 ;
  assign n6760 = ( x65 & n6757 ) | ( x65 & n6759 ) | ( n6757 & n6759 ) ;
  assign n6761 = n6760 ^ n6636 ^ x66 ;
  assign n6762 = ( x66 & n6760 ) | ( x66 & n6761 ) | ( n6760 & n6761 ) ;
  assign n6763 = ( x67 & ~n6755 ) | ( x67 & n6762 ) | ( ~n6755 & n6762 ) ;
  assign n6764 = ( x68 & ~n6652 ) | ( x68 & n6763 ) | ( ~n6652 & n6763 ) ;
  assign n6765 = ( x69 & ~n6629 ) | ( x69 & n6764 ) | ( ~n6629 & n6764 ) ;
  assign n6766 = ( x70 & ~n6711 ) | ( x70 & n6765 ) | ( ~n6711 & n6765 ) ;
  assign n6767 = ( x71 & ~n6708 ) | ( x71 & n6766 ) | ( ~n6708 & n6766 ) ;
  assign n6768 = ( x72 & ~n6642 ) | ( x72 & n6767 ) | ( ~n6642 & n6767 ) ;
  assign n6769 = n6766 ^ n6708 ^ x71 ;
  assign n6770 = ( x73 & ~n6632 ) | ( x73 & n6768 ) | ( ~n6632 & n6768 ) ;
  assign n6771 = ( x74 & ~n6705 ) | ( x74 & n6770 ) | ( ~n6705 & n6770 ) ;
  assign n6772 = ( x75 & ~n6702 ) | ( x75 & n6771 ) | ( ~n6702 & n6771 ) ;
  assign n6773 = ( x76 & ~n6699 ) | ( x76 & n6772 ) | ( ~n6699 & n6772 ) ;
  assign n6774 = ( x77 & ~n6626 ) | ( x77 & n6773 ) | ( ~n6626 & n6773 ) ;
  assign n6775 = ( x78 & ~n6696 ) | ( x78 & n6774 ) | ( ~n6696 & n6774 ) ;
  assign n6776 = ( x79 & ~n6645 ) | ( x79 & n6775 ) | ( ~n6645 & n6775 ) ;
  assign n6777 = ( x80 & ~n6659 ) | ( x80 & n6776 ) | ( ~n6659 & n6776 ) ;
  assign n6778 = ( x81 & ~n6654 ) | ( x81 & n6777 ) | ( ~n6654 & n6777 ) ;
  assign n6779 = ( x82 & ~n6624 ) | ( x82 & n6778 ) | ( ~n6624 & n6778 ) ;
  assign n6780 = ( x83 & ~n6693 ) | ( x83 & n6779 ) | ( ~n6693 & n6779 ) ;
  assign n6781 = ( x84 & ~n6690 ) | ( x84 & n6780 ) | ( ~n6690 & n6780 ) ;
  assign n6782 = ( x85 & ~n6658 ) | ( x85 & n6781 ) | ( ~n6658 & n6781 ) ;
  assign n6783 = ( x86 & ~n6640 ) | ( x86 & n6782 ) | ( ~n6640 & n6782 ) ;
  assign n6784 = ( x87 & ~n6687 ) | ( x87 & n6783 ) | ( ~n6687 & n6783 ) ;
  assign n6785 = ( x88 & ~n6656 ) | ( x88 & n6784 ) | ( ~n6656 & n6784 ) ;
  assign n6786 = ( x89 & ~n6657 ) | ( x89 & n6785 ) | ( ~n6657 & n6785 ) ;
  assign n6787 = ( x90 & ~n6649 ) | ( x90 & n6786 ) | ( ~n6649 & n6786 ) ;
  assign n6788 = ( x91 & ~n6633 ) | ( x91 & n6787 ) | ( ~n6633 & n6787 ) ;
  assign n6789 = ( x92 & ~n6684 ) | ( x92 & n6788 ) | ( ~n6684 & n6788 ) ;
  assign n6790 = n6789 ^ n6681 ^ x93 ;
  assign n6791 = n6768 ^ n6632 ^ x73 ;
  assign n6792 = n6776 ^ n6659 ^ x80 ;
  assign n6793 = n6777 ^ n6654 ^ x81 ;
  assign n6794 = n6778 ^ n6624 ^ x82 ;
  assign n6795 = n6762 ^ n6755 ^ x67 ;
  assign n6796 = n6780 ^ n6690 ^ x84 ;
  assign n6797 = n6781 ^ n6658 ^ x85 ;
  assign n6798 = ( x93 & ~n6681 ) | ( x93 & n6789 ) | ( ~n6681 & n6789 ) ;
  assign n6799 = n6783 ^ n6687 ^ x87 ;
  assign n6800 = n6784 ^ n6656 ^ x88 ;
  assign n6801 = n6763 ^ n6652 ^ x68 ;
  assign n6802 = n6785 ^ n6657 ^ x89 ;
  assign n6803 = n6771 ^ n6702 ^ x75 ;
  assign n6804 = n6773 ^ n6626 ^ x77 ;
  assign n6805 = n6774 ^ n6696 ^ x78 ;
  assign n6806 = n6767 ^ n6642 ^ x72 ;
  assign n6807 = ( x94 & ~n6678 ) | ( x94 & n6798 ) | ( ~n6678 & n6798 ) ;
  assign n6808 = ( x95 & ~n6660 ) | ( x95 & n6807 ) | ( ~n6660 & n6807 ) ;
  assign n6809 = ( x96 & ~n6675 ) | ( x96 & n6808 ) | ( ~n6675 & n6808 ) ;
  assign n6810 = ( x97 & ~n6672 ) | ( x97 & n6809 ) | ( ~n6672 & n6809 ) ;
  assign n6811 = ( x98 & ~n6669 ) | ( x98 & n6810 ) | ( ~n6669 & n6810 ) ;
  assign n6812 = ( x99 & ~n6752 ) | ( x99 & n6811 ) | ( ~n6752 & n6811 ) ;
  assign n6813 = ( x100 & ~n6749 ) | ( x100 & n6812 ) | ( ~n6749 & n6812 ) ;
  assign n6814 = ( x101 & ~n6746 ) | ( x101 & n6813 ) | ( ~n6746 & n6813 ) ;
  assign n6815 = ( x102 & ~n6743 ) | ( x102 & n6814 ) | ( ~n6743 & n6814 ) ;
  assign n6816 = ( x103 & ~n6740 ) | ( x103 & n6815 ) | ( ~n6740 & n6815 ) ;
  assign n6817 = ( x104 & ~n6737 ) | ( x104 & n6816 ) | ( ~n6737 & n6816 ) ;
  assign n6818 = ( x105 & ~n6732 ) | ( x105 & n6817 ) | ( ~n6732 & n6817 ) ;
  assign n6819 = ( x106 & ~n6729 ) | ( x106 & n6818 ) | ( ~n6729 & n6818 ) ;
  assign n6820 = ( x107 & ~n6753 ) | ( x107 & n6819 ) | ( ~n6753 & n6819 ) ;
  assign n6821 = ( x108 & ~n6724 ) | ( x108 & n6820 ) | ( ~n6724 & n6820 ) ;
  assign n6822 = ( x109 & ~n6721 ) | ( x109 & n6821 ) | ( ~n6721 & n6821 ) ;
  assign n6823 = ( x110 & ~n6718 ) | ( x110 & n6822 ) | ( ~n6718 & n6822 ) ;
  assign n6824 = ( x111 & ~n6735 ) | ( x111 & n6823 ) | ( ~n6735 & n6823 ) ;
  assign n6825 = ( x112 & ~n6714 ) | ( x112 & n6824 ) | ( ~n6714 & n6824 ) ;
  assign n6826 = ( x113 & ~n6666 ) | ( x113 & n6825 ) | ( ~n6666 & n6825 ) ;
  assign n6827 = ( x114 & ~n6663 ) | ( x114 & n6826 ) | ( ~n6663 & n6826 ) ;
  assign n6828 = ( x115 & ~n6646 ) | ( x115 & n6827 ) | ( ~n6646 & n6827 ) ;
  assign n6829 = n174 | n6828 ;
  assign n6830 = n6807 ^ n6660 ^ x95 ;
  assign n6831 = n6829 ^ n6660 ^ 1'b0 ;
  assign n6832 = ( n6660 & n6830 ) | ( n6660 & ~n6831 ) | ( n6830 & ~n6831 ) ;
  assign n6833 = n6829 ^ n6681 ^ 1'b0 ;
  assign n6834 = ( n6681 & n6790 ) | ( n6681 & ~n6833 ) | ( n6790 & ~n6833 ) ;
  assign n6835 = n6829 ^ n6657 ^ 1'b0 ;
  assign n6836 = ( n6657 & n6802 ) | ( n6657 & ~n6835 ) | ( n6802 & ~n6835 ) ;
  assign n6837 = n6829 ^ n6656 ^ 1'b0 ;
  assign n6838 = ( n6656 & n6800 ) | ( n6656 & ~n6837 ) | ( n6800 & ~n6837 ) ;
  assign n6839 = n6829 ^ n6687 ^ 1'b0 ;
  assign n6840 = ( n6687 & n6799 ) | ( n6687 & ~n6839 ) | ( n6799 & ~n6839 ) ;
  assign n6841 = n6829 ^ n6658 ^ 1'b0 ;
  assign n6842 = ( n6658 & n6797 ) | ( n6658 & ~n6841 ) | ( n6797 & ~n6841 ) ;
  assign n6843 = n6829 ^ n6690 ^ 1'b0 ;
  assign n6844 = ( n6690 & n6796 ) | ( n6690 & ~n6843 ) | ( n6796 & ~n6843 ) ;
  assign n6845 = n6829 ^ n6624 ^ 1'b0 ;
  assign n6846 = ( n6624 & n6794 ) | ( n6624 & ~n6845 ) | ( n6794 & ~n6845 ) ;
  assign n6847 = n6829 ^ n6654 ^ 1'b0 ;
  assign n6848 = ( n6654 & n6793 ) | ( n6654 & ~n6847 ) | ( n6793 & ~n6847 ) ;
  assign n6849 = n6829 ^ n6659 ^ 1'b0 ;
  assign n6850 = ( n6659 & n6792 ) | ( n6659 & ~n6849 ) | ( n6792 & ~n6849 ) ;
  assign n6851 = n6829 ^ n6696 ^ 1'b0 ;
  assign n6852 = ( n6696 & n6805 ) | ( n6696 & ~n6851 ) | ( n6805 & ~n6851 ) ;
  assign n6853 = n6829 ^ n6626 ^ 1'b0 ;
  assign n6854 = ( n6626 & n6804 ) | ( n6626 & ~n6853 ) | ( n6804 & ~n6853 ) ;
  assign n6855 = n6829 ^ n6702 ^ 1'b0 ;
  assign n6856 = ( n6702 & n6803 ) | ( n6702 & ~n6855 ) | ( n6803 & ~n6855 ) ;
  assign n6857 = n6829 ^ n6632 ^ 1'b0 ;
  assign n6858 = ( n6632 & n6791 ) | ( n6632 & ~n6857 ) | ( n6791 & ~n6857 ) ;
  assign n6859 = n6829 ^ n6642 ^ 1'b0 ;
  assign n6860 = ( n6642 & n6806 ) | ( n6642 & ~n6859 ) | ( n6806 & ~n6859 ) ;
  assign n6861 = n6829 ^ n6708 ^ 1'b0 ;
  assign n6862 = ( n6708 & n6769 ) | ( n6708 & ~n6861 ) | ( n6769 & ~n6861 ) ;
  assign n6863 = n6829 ^ n6652 ^ 1'b0 ;
  assign n6864 = ( n6652 & n6801 ) | ( n6652 & ~n6863 ) | ( n6801 & ~n6863 ) ;
  assign n6865 = n6829 ^ n6755 ^ 1'b0 ;
  assign n6866 = ( n6755 & n6795 ) | ( n6755 & ~n6865 ) | ( n6795 & ~n6865 ) ;
  assign n6867 = n6829 ^ n6759 ^ 1'b0 ;
  assign n6868 = ( n6758 & n6759 ) | ( n6758 & n6867 ) | ( n6759 & n6867 ) ;
  assign n6869 = n6824 ^ n6714 ^ x112 ;
  assign n6870 = n6829 ^ n6714 ^ 1'b0 ;
  assign n6871 = ( n6714 & n6869 ) | ( n6714 & ~n6870 ) | ( n6869 & ~n6870 ) ;
  assign n6872 = n6823 ^ n6735 ^ x111 ;
  assign n6873 = n6829 ^ n6735 ^ 1'b0 ;
  assign n6874 = ( n6735 & n6872 ) | ( n6735 & ~n6873 ) | ( n6872 & ~n6873 ) ;
  assign n6875 = n6821 ^ n6721 ^ x109 ;
  assign n6876 = n6829 ^ n6721 ^ 1'b0 ;
  assign n6877 = ( n6721 & n6875 ) | ( n6721 & ~n6876 ) | ( n6875 & ~n6876 ) ;
  assign n6878 = n6818 ^ n6729 ^ x106 ;
  assign n6879 = n6829 ^ n6729 ^ 1'b0 ;
  assign n6880 = ( n6729 & n6878 ) | ( n6729 & ~n6879 ) | ( n6878 & ~n6879 ) ;
  assign n6881 = n6817 ^ n6732 ^ x105 ;
  assign n6882 = n6829 ^ n6732 ^ 1'b0 ;
  assign n6883 = ( n6732 & n6881 ) | ( n6732 & ~n6882 ) | ( n6881 & ~n6882 ) ;
  assign n6884 = n6816 ^ n6737 ^ x104 ;
  assign n6885 = n6829 ^ n6737 ^ 1'b0 ;
  assign n6886 = ( n6737 & n6884 ) | ( n6737 & ~n6885 ) | ( n6884 & ~n6885 ) ;
  assign n6887 = n6815 ^ n6740 ^ x103 ;
  assign n6888 = n6829 ^ n6740 ^ 1'b0 ;
  assign n6889 = ( n6740 & n6887 ) | ( n6740 & ~n6888 ) | ( n6887 & ~n6888 ) ;
  assign n6890 = n6814 ^ n6743 ^ x102 ;
  assign n6891 = n6829 ^ n6743 ^ 1'b0 ;
  assign n6892 = ( n6743 & n6890 ) | ( n6743 & ~n6891 ) | ( n6890 & ~n6891 ) ;
  assign n6893 = n6809 ^ n6672 ^ x97 ;
  assign n6894 = n6829 ^ n6672 ^ 1'b0 ;
  assign n6895 = ( n6672 & n6893 ) | ( n6672 & ~n6894 ) | ( n6893 & ~n6894 ) ;
  assign n6896 = n6787 ^ n6633 ^ x91 ;
  assign n6897 = n6829 ^ n6633 ^ 1'b0 ;
  assign n6898 = ( n6633 & n6896 ) | ( n6633 & ~n6897 ) | ( n6896 & ~n6897 ) ;
  assign n6899 = n6786 ^ n6649 ^ x90 ;
  assign n6900 = n6829 ^ n6649 ^ 1'b0 ;
  assign n6901 = ( n6649 & n6899 ) | ( n6649 & ~n6900 ) | ( n6899 & ~n6900 ) ;
  assign n6902 = n6779 ^ n6693 ^ x83 ;
  assign n6903 = n6829 ^ n6693 ^ 1'b0 ;
  assign n6904 = ( n6693 & n6902 ) | ( n6693 & ~n6903 ) | ( n6902 & ~n6903 ) ;
  assign n6905 = n6775 ^ n6645 ^ x79 ;
  assign n6906 = n6829 ^ n6645 ^ 1'b0 ;
  assign n6907 = ( n6645 & n6905 ) | ( n6645 & ~n6906 ) | ( n6905 & ~n6906 ) ;
  assign n6908 = n6772 ^ n6699 ^ x76 ;
  assign n6909 = n6829 ^ n6699 ^ 1'b0 ;
  assign n6910 = ( n6699 & n6908 ) | ( n6699 & ~n6909 ) | ( n6908 & ~n6909 ) ;
  assign n6911 = n6770 ^ n6705 ^ x74 ;
  assign n6912 = n6829 ^ n6705 ^ 1'b0 ;
  assign n6913 = ( n6705 & n6911 ) | ( n6705 & ~n6912 ) | ( n6911 & ~n6912 ) ;
  assign n6914 = n6765 ^ n6711 ^ x70 ;
  assign n6915 = n6829 ^ n6711 ^ 1'b0 ;
  assign n6916 = ( n6711 & n6914 ) | ( n6711 & ~n6915 ) | ( n6914 & ~n6915 ) ;
  assign n6917 = n6764 ^ n6629 ^ x69 ;
  assign n6918 = n6829 ^ n6629 ^ 1'b0 ;
  assign n6919 = ( n6629 & n6917 ) | ( n6629 & ~n6918 ) | ( n6917 & ~n6918 ) ;
  assign n6920 = n6826 ^ n6663 ^ x114 ;
  assign n6921 = n6829 ^ n6663 ^ 1'b0 ;
  assign n6922 = ( n6663 & n6920 ) | ( n6663 & ~n6921 ) | ( n6920 & ~n6921 ) ;
  assign n6923 = n6825 ^ n6666 ^ x113 ;
  assign n6924 = n6829 ^ n6666 ^ 1'b0 ;
  assign n6925 = ( n6666 & n6923 ) | ( n6666 & ~n6924 ) | ( n6923 & ~n6924 ) ;
  assign n6926 = n6822 ^ n6718 ^ x110 ;
  assign n6927 = n6829 ^ n6718 ^ 1'b0 ;
  assign n6928 = ( n6718 & n6926 ) | ( n6718 & ~n6927 ) | ( n6926 & ~n6927 ) ;
  assign n6929 = n6820 ^ n6724 ^ x108 ;
  assign n6930 = n6829 ^ n6724 ^ 1'b0 ;
  assign n6931 = ( n6724 & n6929 ) | ( n6724 & ~n6930 ) | ( n6929 & ~n6930 ) ;
  assign n6932 = n6819 ^ n6753 ^ x107 ;
  assign n6933 = n6829 ^ n6753 ^ 1'b0 ;
  assign n6934 = ( n6753 & n6932 ) | ( n6753 & ~n6933 ) | ( n6932 & ~n6933 ) ;
  assign n6935 = n6813 ^ n6746 ^ x101 ;
  assign n6936 = n6829 ^ n6746 ^ 1'b0 ;
  assign n6937 = ( n6746 & n6935 ) | ( n6746 & ~n6936 ) | ( n6935 & ~n6936 ) ;
  assign n6938 = n6812 ^ n6749 ^ x100 ;
  assign n6939 = n6829 ^ n6749 ^ 1'b0 ;
  assign n6940 = ( n6749 & n6938 ) | ( n6749 & ~n6939 ) | ( n6938 & ~n6939 ) ;
  assign n6941 = n6811 ^ n6752 ^ x99 ;
  assign n6942 = n6829 ^ n6752 ^ 1'b0 ;
  assign n6943 = ( n6752 & n6941 ) | ( n6752 & ~n6942 ) | ( n6941 & ~n6942 ) ;
  assign n6944 = n6810 ^ n6669 ^ x98 ;
  assign n6945 = n6829 ^ n6669 ^ 1'b0 ;
  assign n6946 = ( n6669 & n6944 ) | ( n6669 & ~n6945 ) | ( n6944 & ~n6945 ) ;
  assign n6947 = n6808 ^ n6675 ^ x96 ;
  assign n6948 = n6829 ^ n6675 ^ 1'b0 ;
  assign n6949 = ( n6675 & n6947 ) | ( n6675 & ~n6948 ) | ( n6947 & ~n6948 ) ;
  assign n6950 = n6798 ^ n6678 ^ x94 ;
  assign n6951 = n6829 ^ n6678 ^ 1'b0 ;
  assign n6952 = ( n6678 & n6950 ) | ( n6678 & ~n6951 ) | ( n6950 & ~n6951 ) ;
  assign n6953 = n6788 ^ n6684 ^ x92 ;
  assign n6954 = n6829 ^ n6684 ^ 1'b0 ;
  assign n6955 = ( n6684 & n6953 ) | ( n6684 & ~n6954 ) | ( n6953 & ~n6954 ) ;
  assign n6956 = n6782 ^ n6640 ^ x86 ;
  assign n6957 = n6829 ^ n6640 ^ 1'b0 ;
  assign n6958 = ( n6640 & n6956 ) | ( n6640 & ~n6957 ) | ( n6956 & ~n6957 ) ;
  assign n6959 = n6829 ^ n6761 ^ 1'b0 ;
  assign n6960 = ( n6636 & n6761 ) | ( n6636 & n6959 ) | ( n6761 & n6959 ) ;
  assign n6961 = n6827 ^ n6646 ^ x115 ;
  assign n6962 = n6961 ^ n6829 ^ 1'b0 ;
  assign n6963 = ( n6646 & n6961 ) | ( n6646 & n6962 ) | ( n6961 & n6962 ) ;
  assign n6964 = n174 & n6646 ;
  assign n6965 = ~n174 & n6757 ;
  assign n6966 = ( x64 & x116 ) | ( x64 & ~n171 ) | ( x116 & ~n171 ) ;
  assign n6967 = ~x11 & x64 ;
  assign n6968 = n6828 | n6965 ;
  assign n6969 = ( x12 & ~n6828 ) | ( x12 & n6968 ) | ( ~n6828 & n6968 ) ;
  assign n6970 = ~x116 & n6966 ;
  assign n6971 = n6969 & ~n6970 ;
  assign n6972 = ( n6968 & n6969 ) | ( n6968 & n6971 ) | ( n6969 & n6971 ) ;
  assign n6973 = n6972 ^ n6967 ^ x65 ;
  assign n6974 = ( x65 & n6967 ) | ( x65 & n6973 ) | ( n6967 & n6973 ) ;
  assign n6975 = n6974 ^ n6868 ^ x66 ;
  assign n6976 = ( x66 & n6974 ) | ( x66 & n6975 ) | ( n6974 & n6975 ) ;
  assign n6977 = ( x67 & ~n6960 ) | ( x67 & n6976 ) | ( ~n6960 & n6976 ) ;
  assign n6978 = ( x68 & ~n6866 ) | ( x68 & n6977 ) | ( ~n6866 & n6977 ) ;
  assign n6979 = ( x69 & ~n6864 ) | ( x69 & n6978 ) | ( ~n6864 & n6978 ) ;
  assign n6980 = ( x70 & ~n6919 ) | ( x70 & n6979 ) | ( ~n6919 & n6979 ) ;
  assign n6981 = ( x71 & ~n6916 ) | ( x71 & n6980 ) | ( ~n6916 & n6980 ) ;
  assign n6982 = ( x72 & ~n6862 ) | ( x72 & n6981 ) | ( ~n6862 & n6981 ) ;
  assign n6983 = ( x73 & ~n6860 ) | ( x73 & n6982 ) | ( ~n6860 & n6982 ) ;
  assign n6984 = ( x74 & ~n6858 ) | ( x74 & n6983 ) | ( ~n6858 & n6983 ) ;
  assign n6985 = ( x75 & ~n6913 ) | ( x75 & n6984 ) | ( ~n6913 & n6984 ) ;
  assign n6986 = ( x76 & ~n6856 ) | ( x76 & n6985 ) | ( ~n6856 & n6985 ) ;
  assign n6987 = ( x77 & ~n6910 ) | ( x77 & n6986 ) | ( ~n6910 & n6986 ) ;
  assign n6988 = ( x78 & ~n6854 ) | ( x78 & n6987 ) | ( ~n6854 & n6987 ) ;
  assign n6989 = ( x79 & ~n6852 ) | ( x79 & n6988 ) | ( ~n6852 & n6988 ) ;
  assign n6990 = ( x80 & ~n6907 ) | ( x80 & n6989 ) | ( ~n6907 & n6989 ) ;
  assign n6991 = ( x81 & ~n6850 ) | ( x81 & n6990 ) | ( ~n6850 & n6990 ) ;
  assign n6992 = ( x82 & ~n6848 ) | ( x82 & n6991 ) | ( ~n6848 & n6991 ) ;
  assign n6993 = ( x83 & ~n6846 ) | ( x83 & n6992 ) | ( ~n6846 & n6992 ) ;
  assign n6994 = ( x84 & ~n6904 ) | ( x84 & n6993 ) | ( ~n6904 & n6993 ) ;
  assign n6995 = ( x85 & ~n6844 ) | ( x85 & n6994 ) | ( ~n6844 & n6994 ) ;
  assign n6996 = ( x86 & ~n6842 ) | ( x86 & n6995 ) | ( ~n6842 & n6995 ) ;
  assign n6997 = ( x87 & ~n6958 ) | ( x87 & n6996 ) | ( ~n6958 & n6996 ) ;
  assign n6998 = ( x88 & ~n6840 ) | ( x88 & n6997 ) | ( ~n6840 & n6997 ) ;
  assign n6999 = ( x89 & ~n6838 ) | ( x89 & n6998 ) | ( ~n6838 & n6998 ) ;
  assign n7000 = ( x90 & ~n6836 ) | ( x90 & n6999 ) | ( ~n6836 & n6999 ) ;
  assign n7001 = ( x91 & ~n6901 ) | ( x91 & n7000 ) | ( ~n6901 & n7000 ) ;
  assign n7002 = ( x92 & ~n6898 ) | ( x92 & n7001 ) | ( ~n6898 & n7001 ) ;
  assign n7003 = ( x93 & ~n6955 ) | ( x93 & n7002 ) | ( ~n6955 & n7002 ) ;
  assign n7004 = ( x94 & ~n6834 ) | ( x94 & n7003 ) | ( ~n6834 & n7003 ) ;
  assign n7005 = ( x95 & ~n6952 ) | ( x95 & n7004 ) | ( ~n6952 & n7004 ) ;
  assign n7006 = n6996 ^ n6958 ^ x87 ;
  assign n7007 = n6993 ^ n6904 ^ x84 ;
  assign n7008 = ( x96 & ~n6832 ) | ( x96 & n7005 ) | ( ~n6832 & n7005 ) ;
  assign n7009 = n7004 ^ n6952 ^ x95 ;
  assign n7010 = n7008 ^ n6949 ^ x97 ;
  assign n7011 = n7001 ^ n6898 ^ x92 ;
  assign n7012 = n6983 ^ n6858 ^ x74 ;
  assign n7013 = n6987 ^ n6854 ^ x78 ;
  assign n7014 = n6986 ^ n6910 ^ x77 ;
  assign n7015 = n6988 ^ n6852 ^ x79 ;
  assign n7016 = n6981 ^ n6862 ^ x72 ;
  assign n7017 = n6978 ^ n6864 ^ x69 ;
  assign n7018 = ( x97 & ~n6949 ) | ( x97 & n7008 ) | ( ~n6949 & n7008 ) ;
  assign n7019 = ( x98 & ~n6895 ) | ( x98 & n7018 ) | ( ~n6895 & n7018 ) ;
  assign n7020 = ( x99 & ~n6946 ) | ( x99 & n7019 ) | ( ~n6946 & n7019 ) ;
  assign n7021 = ( x100 & ~n6943 ) | ( x100 & n7020 ) | ( ~n6943 & n7020 ) ;
  assign n7022 = ( x101 & ~n6940 ) | ( x101 & n7021 ) | ( ~n6940 & n7021 ) ;
  assign n7023 = ( x102 & ~n6937 ) | ( x102 & n7022 ) | ( ~n6937 & n7022 ) ;
  assign n7024 = ( x103 & ~n6892 ) | ( x103 & n7023 ) | ( ~n6892 & n7023 ) ;
  assign n7025 = ( x116 & n171 ) | ( x116 & ~n6963 ) | ( n171 & ~n6963 ) ;
  assign n7026 = ( x104 & ~n6889 ) | ( x104 & n7024 ) | ( ~n6889 & n7024 ) ;
  assign n7027 = ( x105 & ~n6886 ) | ( x105 & n7026 ) | ( ~n6886 & n7026 ) ;
  assign n7028 = ( x106 & ~n6883 ) | ( x106 & n7027 ) | ( ~n6883 & n7027 ) ;
  assign n7029 = ( x107 & ~n6880 ) | ( x107 & n7028 ) | ( ~n6880 & n7028 ) ;
  assign n7030 = ( x108 & ~n6934 ) | ( x108 & n7029 ) | ( ~n6934 & n7029 ) ;
  assign n7031 = ( x109 & ~n6931 ) | ( x109 & n7030 ) | ( ~n6931 & n7030 ) ;
  assign n7032 = ( x110 & ~n6877 ) | ( x110 & n7031 ) | ( ~n6877 & n7031 ) ;
  assign n7033 = ( x111 & ~n6928 ) | ( x111 & n7032 ) | ( ~n6928 & n7032 ) ;
  assign n7034 = ( x112 & ~n6874 ) | ( x112 & n7033 ) | ( ~n6874 & n7033 ) ;
  assign n7035 = n7024 ^ n6889 ^ x104 ;
  assign n7036 = ( x113 & ~n6871 ) | ( x113 & n7034 ) | ( ~n6871 & n7034 ) ;
  assign n7037 = n7020 ^ n6943 ^ x100 ;
  assign n7038 = ( x114 & ~n6925 ) | ( x114 & n7036 ) | ( ~n6925 & n7036 ) ;
  assign n7039 = ( x115 & ~n6922 ) | ( x115 & n7038 ) | ( ~n6922 & n7038 ) ;
  assign n7040 = ( ~x116 & n6963 ) | ( ~x116 & n7039 ) | ( n6963 & n7039 ) ;
  assign n7041 = n7025 | n7040 ;
  assign n7042 = n174 & n6963 ;
  assign n7043 = n7039 ^ n6963 ^ x116 ;
  assign n7044 = ( ~n6963 & n7041 ) | ( ~n6963 & n7042 ) | ( n7041 & n7042 ) ;
  assign n7045 = n7043 & ~n7044 ;
  assign n7046 = n7044 ^ n6949 ^ 1'b0 ;
  assign n7047 = ( n6949 & n7010 ) | ( n6949 & ~n7046 ) | ( n7010 & ~n7046 ) ;
  assign n7048 = n7044 ^ n6910 ^ 1'b0 ;
  assign n7049 = n6964 & ~n7041 ;
  assign n7050 = n7044 ^ n6975 ^ 1'b0 ;
  assign n7051 = ( n6868 & n6975 ) | ( n6868 & n7050 ) | ( n6975 & n7050 ) ;
  assign n7052 = n7044 ^ n6858 ^ 1'b0 ;
  assign n7053 = ( n6858 & n7012 ) | ( n6858 & ~n7052 ) | ( n7012 & ~n7052 ) ;
  assign n7054 = n7044 ^ n6864 ^ 1'b0 ;
  assign n7055 = ( n6910 & n7014 ) | ( n6910 & ~n7048 ) | ( n7014 & ~n7048 ) ;
  assign n7056 = n7044 ^ n6973 ^ 1'b0 ;
  assign n7057 = ( n6864 & n7017 ) | ( n6864 & ~n7054 ) | ( n7017 & ~n7054 ) ;
  assign n7058 = ( n6972 & n6973 ) | ( n6972 & n7056 ) | ( n6973 & n7056 ) ;
  assign n7059 = n7044 ^ n6952 ^ 1'b0 ;
  assign n7060 = ( n6952 & n7009 ) | ( n6952 & ~n7059 ) | ( n7009 & ~n7059 ) ;
  assign n7061 = n7044 ^ n6862 ^ 1'b0 ;
  assign n7062 = ( n6862 & n7016 ) | ( n6862 & ~n7061 ) | ( n7016 & ~n7061 ) ;
  assign n7063 = n7044 ^ n6943 ^ 1'b0 ;
  assign n7064 = ( n6943 & n7037 ) | ( n6943 & ~n7063 ) | ( n7037 & ~n7063 ) ;
  assign n7065 = n7044 ^ n6904 ^ 1'b0 ;
  assign n7066 = n7044 ^ n6958 ^ 1'b0 ;
  assign n7067 = ( n6958 & n7006 ) | ( n6958 & ~n7066 ) | ( n7006 & ~n7066 ) ;
  assign n7068 = n7044 ^ n6852 ^ 1'b0 ;
  assign n7069 = n7044 ^ n6889 ^ 1'b0 ;
  assign n7070 = n7044 ^ n6892 ^ 1'b0 ;
  assign n7071 = ( n6904 & n7007 ) | ( n6904 & ~n7065 ) | ( n7007 & ~n7065 ) ;
  assign n7072 = ( n6889 & n7035 ) | ( n6889 & ~n7069 ) | ( n7035 & ~n7069 ) ;
  assign n7073 = n7023 ^ n6892 ^ x103 ;
  assign n7074 = n7044 ^ n6898 ^ 1'b0 ;
  assign n7075 = n7044 ^ n6854 ^ 1'b0 ;
  assign n7076 = ( n6854 & n7013 ) | ( n6854 & ~n7075 ) | ( n7013 & ~n7075 ) ;
  assign n7077 = ( n6892 & ~n7070 ) | ( n6892 & n7073 ) | ( ~n7070 & n7073 ) ;
  assign n7078 = ( n6898 & n7011 ) | ( n6898 & ~n7074 ) | ( n7011 & ~n7074 ) ;
  assign n7079 = ( n6852 & n7015 ) | ( n6852 & ~n7068 ) | ( n7015 & ~n7068 ) ;
  assign n7080 = ( n6964 & n7045 ) | ( n6964 & ~n7049 ) | ( n7045 & ~n7049 ) ;
  assign n7081 = n7038 ^ n6922 ^ x115 ;
  assign n7082 = n7044 ^ n6922 ^ 1'b0 ;
  assign n7083 = ( n6922 & n7081 ) | ( n6922 & ~n7082 ) | ( n7081 & ~n7082 ) ;
  assign n7084 = n7036 ^ n6925 ^ x114 ;
  assign n7085 = n7044 ^ n6925 ^ 1'b0 ;
  assign n7086 = ( n6925 & n7084 ) | ( n6925 & ~n7085 ) | ( n7084 & ~n7085 ) ;
  assign n7087 = n6998 ^ n6838 ^ x89 ;
  assign n7088 = n7044 ^ n6838 ^ 1'b0 ;
  assign n7089 = ( n6838 & n7087 ) | ( n6838 & ~n7088 ) | ( n7087 & ~n7088 ) ;
  assign n7090 = n6997 ^ n6840 ^ x88 ;
  assign n7091 = n7044 ^ n6840 ^ 1'b0 ;
  assign n7092 = ( n6840 & n7090 ) | ( n6840 & ~n7091 ) | ( n7090 & ~n7091 ) ;
  assign n7093 = n6995 ^ n6842 ^ x86 ;
  assign n7094 = n7044 ^ n6842 ^ 1'b0 ;
  assign n7095 = ( n6842 & n7093 ) | ( n6842 & ~n7094 ) | ( n7093 & ~n7094 ) ;
  assign n7096 = n6994 ^ n6844 ^ x85 ;
  assign n7097 = n7044 ^ n6844 ^ 1'b0 ;
  assign n7098 = ( n6844 & n7096 ) | ( n6844 & ~n7097 ) | ( n7096 & ~n7097 ) ;
  assign n7099 = n6992 ^ n6846 ^ x83 ;
  assign n7100 = n7044 ^ n6846 ^ 1'b0 ;
  assign n7101 = ( n6846 & n7099 ) | ( n6846 & ~n7100 ) | ( n7099 & ~n7100 ) ;
  assign n7102 = n6991 ^ n6848 ^ x82 ;
  assign n7103 = n7044 ^ n6848 ^ 1'b0 ;
  assign n7104 = ( n6848 & n7102 ) | ( n6848 & ~n7103 ) | ( n7102 & ~n7103 ) ;
  assign n7105 = n6990 ^ n6850 ^ x81 ;
  assign n7106 = n7044 ^ n6850 ^ 1'b0 ;
  assign n7107 = ( n6850 & n7105 ) | ( n6850 & ~n7106 ) | ( n7105 & ~n7106 ) ;
  assign n7108 = n6989 ^ n6907 ^ x80 ;
  assign n7109 = n7044 ^ n6907 ^ 1'b0 ;
  assign n7110 = ( n6907 & n7108 ) | ( n6907 & ~n7109 ) | ( n7108 & ~n7109 ) ;
  assign n7111 = n6985 ^ n6856 ^ x76 ;
  assign n7112 = n7044 ^ n6856 ^ 1'b0 ;
  assign n7113 = ( n6856 & n7111 ) | ( n6856 & ~n7112 ) | ( n7111 & ~n7112 ) ;
  assign n7114 = n6984 ^ n6913 ^ x75 ;
  assign n7115 = n7044 ^ n6913 ^ 1'b0 ;
  assign n7116 = ( n6913 & n7114 ) | ( n6913 & ~n7115 ) | ( n7114 & ~n7115 ) ;
  assign n7117 = n6982 ^ n6860 ^ x73 ;
  assign n7118 = n7044 ^ n6860 ^ 1'b0 ;
  assign n7119 = ( n6860 & n7117 ) | ( n6860 & ~n7118 ) | ( n7117 & ~n7118 ) ;
  assign n7120 = n6980 ^ n6916 ^ x71 ;
  assign n7121 = n7044 ^ n6916 ^ 1'b0 ;
  assign n7122 = ( n6916 & n7120 ) | ( n6916 & ~n7121 ) | ( n7120 & ~n7121 ) ;
  assign n7123 = n6979 ^ n6919 ^ x70 ;
  assign n7124 = n7044 ^ n6919 ^ 1'b0 ;
  assign n7125 = ( n6919 & n7123 ) | ( n6919 & ~n7124 ) | ( n7123 & ~n7124 ) ;
  assign n7126 = n6977 ^ n6866 ^ x68 ;
  assign n7127 = n7044 ^ n6866 ^ 1'b0 ;
  assign n7128 = ( n6866 & n7126 ) | ( n6866 & ~n7127 ) | ( n7126 & ~n7127 ) ;
  assign n7129 = n6976 ^ n6960 ^ x67 ;
  assign n7130 = n7044 ^ n6960 ^ 1'b0 ;
  assign n7131 = ( n6960 & n7129 ) | ( n6960 & ~n7130 ) | ( n7129 & ~n7130 ) ;
  assign n7132 = n7034 ^ n6871 ^ x113 ;
  assign n7133 = n7044 ^ n6871 ^ 1'b0 ;
  assign n7134 = ( n6871 & n7132 ) | ( n6871 & ~n7133 ) | ( n7132 & ~n7133 ) ;
  assign n7135 = n7030 ^ n6931 ^ x109 ;
  assign n7136 = n7044 ^ n6931 ^ 1'b0 ;
  assign n7137 = ( n6931 & n7135 ) | ( n6931 & ~n7136 ) | ( n7135 & ~n7136 ) ;
  assign n7138 = n7029 ^ n6934 ^ x108 ;
  assign n7139 = n7044 ^ n6934 ^ 1'b0 ;
  assign n7140 = ( n6934 & n7138 ) | ( n6934 & ~n7139 ) | ( n7138 & ~n7139 ) ;
  assign n7141 = n7028 ^ n6880 ^ x107 ;
  assign n7142 = n7044 ^ n6880 ^ 1'b0 ;
  assign n7143 = ( n6880 & n7141 ) | ( n6880 & ~n7142 ) | ( n7141 & ~n7142 ) ;
  assign n7144 = n7027 ^ n6883 ^ x106 ;
  assign n7145 = n7044 ^ n6883 ^ 1'b0 ;
  assign n7146 = ( n6883 & n7144 ) | ( n6883 & ~n7145 ) | ( n7144 & ~n7145 ) ;
  assign n7147 = n7026 ^ n6886 ^ x105 ;
  assign n7148 = n7044 ^ n6886 ^ 1'b0 ;
  assign n7149 = ( n6886 & n7147 ) | ( n6886 & ~n7148 ) | ( n7147 & ~n7148 ) ;
  assign n7150 = n7022 ^ n6937 ^ x102 ;
  assign n7151 = n7044 ^ n6937 ^ 1'b0 ;
  assign n7152 = ( n6937 & n7150 ) | ( n6937 & ~n7151 ) | ( n7150 & ~n7151 ) ;
  assign n7153 = n7021 ^ n6940 ^ x101 ;
  assign n7154 = n7044 ^ n6940 ^ 1'b0 ;
  assign n7155 = ( n6940 & n7153 ) | ( n6940 & ~n7154 ) | ( n7153 & ~n7154 ) ;
  assign n7156 = n7019 ^ n6946 ^ x99 ;
  assign n7157 = n7044 ^ n6946 ^ 1'b0 ;
  assign n7158 = ( n6946 & n7156 ) | ( n6946 & ~n7157 ) | ( n7156 & ~n7157 ) ;
  assign n7159 = n7018 ^ n6895 ^ x98 ;
  assign n7160 = n7044 ^ n6895 ^ 1'b0 ;
  assign n7161 = ( n6895 & n7159 ) | ( n6895 & ~n7160 ) | ( n7159 & ~n7160 ) ;
  assign n7162 = n7005 ^ n6832 ^ x96 ;
  assign n7163 = n7044 ^ n6832 ^ 1'b0 ;
  assign n7164 = ( n6832 & n7162 ) | ( n6832 & ~n7163 ) | ( n7162 & ~n7163 ) ;
  assign n7165 = n7003 ^ n6834 ^ x94 ;
  assign n7166 = n7044 ^ n6834 ^ 1'b0 ;
  assign n7167 = ( n6834 & n7165 ) | ( n6834 & ~n7166 ) | ( n7165 & ~n7166 ) ;
  assign n7168 = n7002 ^ n6955 ^ x93 ;
  assign n7169 = n7044 ^ n6955 ^ 1'b0 ;
  assign n7170 = ( n6955 & n7168 ) | ( n6955 & ~n7169 ) | ( n7168 & ~n7169 ) ;
  assign n7171 = n7000 ^ n6901 ^ x91 ;
  assign n7172 = n7044 ^ n6901 ^ 1'b0 ;
  assign n7173 = ( n6901 & n7171 ) | ( n6901 & ~n7172 ) | ( n7171 & ~n7172 ) ;
  assign n7174 = n6999 ^ n6836 ^ x90 ;
  assign n7175 = n7044 ^ n6836 ^ 1'b0 ;
  assign n7176 = ( n6836 & n7174 ) | ( n6836 & ~n7175 ) | ( n7174 & ~n7175 ) ;
  assign n7177 = x64 & n7044 ;
  assign n7178 = n7177 ^ x64 ^ x11 ;
  assign n7179 = ( ~x118 & x119 ) | ( ~x118 & n163 ) | ( x119 & n163 ) ;
  assign n7180 = ~x10 & x64 ;
  assign n7181 = n7180 ^ n7178 ^ x65 ;
  assign n7182 = ( x65 & n7180 ) | ( x65 & n7181 ) | ( n7180 & n7181 ) ;
  assign n7183 = n7182 ^ n7058 ^ x66 ;
  assign n7184 = ( x66 & n7182 ) | ( x66 & n7183 ) | ( n7182 & n7183 ) ;
  assign n7185 = ( x67 & ~n7051 ) | ( x67 & n7184 ) | ( ~n7051 & n7184 ) ;
  assign n7186 = ( x68 & ~n7131 ) | ( x68 & n7185 ) | ( ~n7131 & n7185 ) ;
  assign n7187 = x118 | n7179 ;
  assign n7188 = n7186 ^ n7128 ^ x69 ;
  assign n7189 = ( x69 & ~n7128 ) | ( x69 & n7186 ) | ( ~n7128 & n7186 ) ;
  assign n7190 = ( x70 & ~n7057 ) | ( x70 & n7189 ) | ( ~n7057 & n7189 ) ;
  assign n7191 = ( x71 & ~n7125 ) | ( x71 & n7190 ) | ( ~n7125 & n7190 ) ;
  assign n7192 = ( x72 & ~n7122 ) | ( x72 & n7191 ) | ( ~n7122 & n7191 ) ;
  assign n7193 = ( x73 & ~n7062 ) | ( x73 & n7192 ) | ( ~n7062 & n7192 ) ;
  assign n7194 = ( x74 & ~n7119 ) | ( x74 & n7193 ) | ( ~n7119 & n7193 ) ;
  assign n7195 = ( x75 & ~n7053 ) | ( x75 & n7194 ) | ( ~n7053 & n7194 ) ;
  assign n7196 = ( x76 & ~n7116 ) | ( x76 & n7195 ) | ( ~n7116 & n7195 ) ;
  assign n7197 = ( x77 & ~n7113 ) | ( x77 & n7196 ) | ( ~n7113 & n7196 ) ;
  assign n7198 = ( x78 & ~n7055 ) | ( x78 & n7197 ) | ( ~n7055 & n7197 ) ;
  assign n7199 = ( x79 & ~n7076 ) | ( x79 & n7198 ) | ( ~n7076 & n7198 ) ;
  assign n7200 = ( x80 & ~n7079 ) | ( x80 & n7199 ) | ( ~n7079 & n7199 ) ;
  assign n7201 = n7194 ^ n7053 ^ x75 ;
  assign n7202 = ( x81 & ~n7110 ) | ( x81 & n7200 ) | ( ~n7110 & n7200 ) ;
  assign n7203 = ( x82 & ~n7107 ) | ( x82 & n7202 ) | ( ~n7107 & n7202 ) ;
  assign n7204 = n7044 ^ n6928 ^ 1'b0 ;
  assign n7205 = n7198 ^ n7076 ^ x79 ;
  assign n7206 = ( x83 & ~n7104 ) | ( x83 & n7203 ) | ( ~n7104 & n7203 ) ;
  assign n7207 = n7031 ^ n6877 ^ x110 ;
  assign n7208 = n7032 ^ n6928 ^ x111 ;
  assign n7209 = n7202 ^ n7107 ^ x82 ;
  assign n7210 = n7203 ^ n7104 ^ x83 ;
  assign n7211 = n7033 ^ n6874 ^ x112 ;
  assign n7212 = n7044 ^ n6874 ^ 1'b0 ;
  assign n7213 = ( n6874 & n7211 ) | ( n6874 & ~n7212 ) | ( n7211 & ~n7212 ) ;
  assign n7214 = ( x84 & ~n7101 ) | ( x84 & n7206 ) | ( ~n7101 & n7206 ) ;
  assign n7215 = ( x85 & ~n7071 ) | ( x85 & n7214 ) | ( ~n7071 & n7214 ) ;
  assign n7216 = ( x86 & ~n7098 ) | ( x86 & n7215 ) | ( ~n7098 & n7215 ) ;
  assign n7217 = ( x87 & ~n7095 ) | ( x87 & n7216 ) | ( ~n7095 & n7216 ) ;
  assign n7218 = ( x88 & ~n7067 ) | ( x88 & n7217 ) | ( ~n7067 & n7217 ) ;
  assign n7219 = n7216 ^ n7095 ^ x87 ;
  assign n7220 = ( n6928 & ~n7204 ) | ( n6928 & n7208 ) | ( ~n7204 & n7208 ) ;
  assign n7221 = ( x89 & ~n7092 ) | ( x89 & n7218 ) | ( ~n7092 & n7218 ) ;
  assign n7222 = n7044 ^ n6877 ^ 1'b0 ;
  assign n7223 = ( n6877 & n7207 ) | ( n6877 & ~n7222 ) | ( n7207 & ~n7222 ) ;
  assign n7224 = ( x90 & ~n7089 ) | ( x90 & n7221 ) | ( ~n7089 & n7221 ) ;
  assign n7225 = ( x91 & ~n7176 ) | ( x91 & n7224 ) | ( ~n7176 & n7224 ) ;
  assign n7226 = n7225 ^ n7173 ^ x92 ;
  assign n7227 = ( x92 & ~n7173 ) | ( x92 & n7225 ) | ( ~n7173 & n7225 ) ;
  assign n7228 = ( x93 & ~n7078 ) | ( x93 & n7227 ) | ( ~n7078 & n7227 ) ;
  assign n7229 = ( x94 & ~n7170 ) | ( x94 & n7228 ) | ( ~n7170 & n7228 ) ;
  assign n7230 = ( x95 & ~n7167 ) | ( x95 & n7229 ) | ( ~n7167 & n7229 ) ;
  assign n7231 = ( x96 & ~n7060 ) | ( x96 & n7230 ) | ( ~n7060 & n7230 ) ;
  assign n7232 = ( x97 & ~n7164 ) | ( x97 & n7231 ) | ( ~n7164 & n7231 ) ;
  assign n7233 = ( x98 & ~n7047 ) | ( x98 & n7232 ) | ( ~n7047 & n7232 ) ;
  assign n7234 = ( x99 & ~n7161 ) | ( x99 & n7233 ) | ( ~n7161 & n7233 ) ;
  assign n7235 = ( x100 & ~n7158 ) | ( x100 & n7234 ) | ( ~n7158 & n7234 ) ;
  assign n7236 = ( x101 & ~n7064 ) | ( x101 & n7235 ) | ( ~n7064 & n7235 ) ;
  assign n7237 = ( x102 & ~n7155 ) | ( x102 & n7236 ) | ( ~n7155 & n7236 ) ;
  assign n7238 = ( x103 & ~n7152 ) | ( x103 & n7237 ) | ( ~n7152 & n7237 ) ;
  assign n7239 = ( x104 & ~n7077 ) | ( x104 & n7238 ) | ( ~n7077 & n7238 ) ;
  assign n7240 = ( ~x117 & n7080 ) | ( ~x117 & n7187 ) | ( n7080 & n7187 ) ;
  assign n7241 = ( x105 & ~n7072 ) | ( x105 & n7239 ) | ( ~n7072 & n7239 ) ;
  assign n7242 = n7229 ^ n7167 ^ x95 ;
  assign n7243 = ( x106 & ~n7149 ) | ( x106 & n7241 ) | ( ~n7149 & n7241 ) ;
  assign n7244 = ( x107 & ~n7146 ) | ( x107 & n7243 ) | ( ~n7146 & n7243 ) ;
  assign n7245 = ( x108 & ~n7143 ) | ( x108 & n7244 ) | ( ~n7143 & n7244 ) ;
  assign n7246 = ( x109 & ~n7140 ) | ( x109 & n7245 ) | ( ~n7140 & n7245 ) ;
  assign n7247 = ( x110 & ~n7137 ) | ( x110 & n7246 ) | ( ~n7137 & n7246 ) ;
  assign n7248 = ( x111 & ~n7223 ) | ( x111 & n7247 ) | ( ~n7223 & n7247 ) ;
  assign n7249 = ( x112 & ~n7220 ) | ( x112 & n7248 ) | ( ~n7220 & n7248 ) ;
  assign n7250 = ( x113 & ~n7213 ) | ( x113 & n7249 ) | ( ~n7213 & n7249 ) ;
  assign n7251 = ( x114 & ~n7134 ) | ( x114 & n7250 ) | ( ~n7134 & n7250 ) ;
  assign n7252 = ( x115 & ~n7086 ) | ( x115 & n7251 ) | ( ~n7086 & n7251 ) ;
  assign n7253 = ( x116 & ~n7083 ) | ( x116 & n7252 ) | ( ~n7083 & n7252 ) ;
  assign n7254 = ( x117 & ~n7080 ) | ( x117 & n7253 ) | ( ~n7080 & n7253 ) ;
  assign n7255 = n7240 | n7254 ;
  assign n7256 = n7253 ^ n7080 ^ x117 ;
  assign n7257 = n171 & n7080 ;
  assign n7258 = ( ~n7080 & n7255 ) | ( ~n7080 & n7257 ) | ( n7255 & n7257 ) ;
  assign n7259 = n7256 & ~n7258 ;
  assign n7260 = ~n7255 & n7257 ;
  assign n7261 = n7246 ^ n7137 ^ x110 ;
  assign n7262 = ( n7257 & n7259 ) | ( n7257 & ~n7260 ) | ( n7259 & ~n7260 ) ;
  assign n7263 = n7258 ^ n7053 ^ 1'b0 ;
  assign n7264 = n7258 ^ n7167 ^ 1'b0 ;
  assign n7265 = ( n7053 & n7201 ) | ( n7053 & ~n7263 ) | ( n7201 & ~n7263 ) ;
  assign n7266 = ( n7167 & n7242 ) | ( n7167 & ~n7264 ) | ( n7242 & ~n7264 ) ;
  assign n7267 = n7230 ^ n7060 ^ x96 ;
  assign n7268 = n7258 ^ n7104 ^ 1'b0 ;
  assign n7269 = n7258 ^ n7107 ^ 1'b0 ;
  assign n7270 = n7258 ^ n7183 ^ 1'b0 ;
  assign n7271 = n7258 ^ n7128 ^ 1'b0 ;
  assign n7272 = ( n7128 & n7188 ) | ( n7128 & ~n7271 ) | ( n7188 & ~n7271 ) ;
  assign n7273 = ( n7107 & n7209 ) | ( n7107 & ~n7269 ) | ( n7209 & ~n7269 ) ;
  assign n7274 = n7258 ^ n7060 ^ 1'b0 ;
  assign n7275 = n7258 ^ n7076 ^ 1'b0 ;
  assign n7276 = ( n7104 & n7210 ) | ( n7104 & ~n7268 ) | ( n7210 & ~n7268 ) ;
  assign n7277 = n7258 ^ n7095 ^ 1'b0 ;
  assign n7278 = ( n7076 & n7205 ) | ( n7076 & ~n7275 ) | ( n7205 & ~n7275 ) ;
  assign n7279 = n7258 ^ n7181 ^ 1'b0 ;
  assign n7280 = ( n7060 & n7267 ) | ( n7060 & ~n7274 ) | ( n7267 & ~n7274 ) ;
  assign n7281 = ( n7095 & n7219 ) | ( n7095 & ~n7277 ) | ( n7219 & ~n7277 ) ;
  assign n7282 = n7258 ^ n7137 ^ 1'b0 ;
  assign n7283 = ( n7137 & n7261 ) | ( n7137 & ~n7282 ) | ( n7261 & ~n7282 ) ;
  assign n7284 = ( n7178 & n7181 ) | ( n7178 & n7279 ) | ( n7181 & n7279 ) ;
  assign n7285 = ( n7058 & n7183 ) | ( n7058 & n7270 ) | ( n7183 & n7270 ) ;
  assign n7286 = n7258 ^ n7173 ^ 1'b0 ;
  assign n7287 = ( n7173 & n7226 ) | ( n7173 & ~n7286 ) | ( n7226 & ~n7286 ) ;
  assign n7288 = n7252 ^ n7083 ^ x116 ;
  assign n7289 = n7258 ^ n7083 ^ 1'b0 ;
  assign n7290 = ( n7083 & n7288 ) | ( n7083 & ~n7289 ) | ( n7288 & ~n7289 ) ;
  assign n7291 = n7251 ^ n7086 ^ x115 ;
  assign n7292 = n7258 ^ n7086 ^ 1'b0 ;
  assign n7293 = ( n7086 & n7291 ) | ( n7086 & ~n7292 ) | ( n7291 & ~n7292 ) ;
  assign n7294 = n7250 ^ n7134 ^ x114 ;
  assign n7295 = n7258 ^ n7134 ^ 1'b0 ;
  assign n7296 = ( n7134 & n7294 ) | ( n7134 & ~n7295 ) | ( n7294 & ~n7295 ) ;
  assign n7297 = n7214 ^ n7071 ^ x85 ;
  assign n7298 = n7258 ^ n7071 ^ 1'b0 ;
  assign n7299 = ( n7071 & n7297 ) | ( n7071 & ~n7298 ) | ( n7297 & ~n7298 ) ;
  assign n7300 = n7206 ^ n7101 ^ x84 ;
  assign n7301 = n7258 ^ n7101 ^ 1'b0 ;
  assign n7302 = ( n7101 & n7300 ) | ( n7101 & ~n7301 ) | ( n7300 & ~n7301 ) ;
  assign n7303 = n7200 ^ n7110 ^ x81 ;
  assign n7304 = n7258 ^ n7110 ^ 1'b0 ;
  assign n7305 = ( n7110 & n7303 ) | ( n7110 & ~n7304 ) | ( n7303 & ~n7304 ) ;
  assign n7306 = n7199 ^ n7079 ^ x80 ;
  assign n7307 = n7258 ^ n7079 ^ 1'b0 ;
  assign n7308 = ( n7079 & n7306 ) | ( n7079 & ~n7307 ) | ( n7306 & ~n7307 ) ;
  assign n7309 = n7197 ^ n7055 ^ x78 ;
  assign n7310 = n7258 ^ n7055 ^ 1'b0 ;
  assign n7311 = ( n7055 & n7309 ) | ( n7055 & ~n7310 ) | ( n7309 & ~n7310 ) ;
  assign n7312 = n7196 ^ n7113 ^ x77 ;
  assign n7313 = n7258 ^ n7113 ^ 1'b0 ;
  assign n7314 = ( n7113 & n7312 ) | ( n7113 & ~n7313 ) | ( n7312 & ~n7313 ) ;
  assign n7315 = n7195 ^ n7116 ^ x76 ;
  assign n7316 = n7258 ^ n7116 ^ 1'b0 ;
  assign n7317 = ( n7116 & n7315 ) | ( n7116 & ~n7316 ) | ( n7315 & ~n7316 ) ;
  assign n7318 = n7193 ^ n7119 ^ x74 ;
  assign n7319 = n7258 ^ n7119 ^ 1'b0 ;
  assign n7320 = ( n7119 & n7318 ) | ( n7119 & ~n7319 ) | ( n7318 & ~n7319 ) ;
  assign n7321 = n7192 ^ n7062 ^ x73 ;
  assign n7322 = n7258 ^ n7062 ^ 1'b0 ;
  assign n7323 = ( n7062 & n7321 ) | ( n7062 & ~n7322 ) | ( n7321 & ~n7322 ) ;
  assign n7324 = n7191 ^ n7122 ^ x72 ;
  assign n7325 = n7258 ^ n7122 ^ 1'b0 ;
  assign n7326 = ( n7122 & n7324 ) | ( n7122 & ~n7325 ) | ( n7324 & ~n7325 ) ;
  assign n7327 = n7190 ^ n7125 ^ x71 ;
  assign n7328 = n7258 ^ n7125 ^ 1'b0 ;
  assign n7329 = ( n7125 & n7327 ) | ( n7125 & ~n7328 ) | ( n7327 & ~n7328 ) ;
  assign n7330 = n7189 ^ n7057 ^ x70 ;
  assign n7331 = n7258 ^ n7057 ^ 1'b0 ;
  assign n7332 = ( n7057 & n7330 ) | ( n7057 & ~n7331 ) | ( n7330 & ~n7331 ) ;
  assign n7333 = n7185 ^ n7131 ^ x68 ;
  assign n7334 = n7258 ^ n7131 ^ 1'b0 ;
  assign n7335 = ( n7131 & n7333 ) | ( n7131 & ~n7334 ) | ( n7333 & ~n7334 ) ;
  assign n7336 = n7184 ^ n7051 ^ x67 ;
  assign n7337 = n7258 ^ n7051 ^ 1'b0 ;
  assign n7338 = ( n7051 & n7336 ) | ( n7051 & ~n7337 ) | ( n7336 & ~n7337 ) ;
  assign n7339 = n7249 ^ n7213 ^ x113 ;
  assign n7340 = n7258 ^ n7213 ^ 1'b0 ;
  assign n7341 = ( n7213 & n7339 ) | ( n7213 & ~n7340 ) | ( n7339 & ~n7340 ) ;
  assign n7342 = n7248 ^ n7220 ^ x112 ;
  assign n7343 = n7258 ^ n7220 ^ 1'b0 ;
  assign n7344 = ( n7220 & n7342 ) | ( n7220 & ~n7343 ) | ( n7342 & ~n7343 ) ;
  assign n7345 = n7247 ^ n7223 ^ x111 ;
  assign n7346 = n7258 ^ n7223 ^ 1'b0 ;
  assign n7347 = ( n7223 & n7345 ) | ( n7223 & ~n7346 ) | ( n7345 & ~n7346 ) ;
  assign n7348 = n7245 ^ n7140 ^ x109 ;
  assign n7349 = n7258 ^ n7140 ^ 1'b0 ;
  assign n7350 = ( n7140 & n7348 ) | ( n7140 & ~n7349 ) | ( n7348 & ~n7349 ) ;
  assign n7351 = n7244 ^ n7143 ^ x108 ;
  assign n7352 = n7258 ^ n7143 ^ 1'b0 ;
  assign n7353 = ( n7143 & n7351 ) | ( n7143 & ~n7352 ) | ( n7351 & ~n7352 ) ;
  assign n7354 = n7243 ^ n7146 ^ x107 ;
  assign n7355 = n7258 ^ n7146 ^ 1'b0 ;
  assign n7356 = ( n7146 & n7354 ) | ( n7146 & ~n7355 ) | ( n7354 & ~n7355 ) ;
  assign n7357 = n7231 ^ n7164 ^ x97 ;
  assign n7358 = n7258 ^ n7164 ^ 1'b0 ;
  assign n7359 = ( n7164 & n7357 ) | ( n7164 & ~n7358 ) | ( n7357 & ~n7358 ) ;
  assign n7360 = n7228 ^ n7170 ^ x94 ;
  assign n7361 = n7258 ^ n7170 ^ 1'b0 ;
  assign n7362 = ( n7170 & n7360 ) | ( n7170 & ~n7361 ) | ( n7360 & ~n7361 ) ;
  assign n7363 = n7227 ^ n7078 ^ x93 ;
  assign n7364 = n7258 ^ n7078 ^ 1'b0 ;
  assign n7365 = ( n7078 & n7363 ) | ( n7078 & ~n7364 ) | ( n7363 & ~n7364 ) ;
  assign n7366 = n7224 ^ n7176 ^ x91 ;
  assign n7367 = n7258 ^ n7176 ^ 1'b0 ;
  assign n7368 = ( n7176 & n7366 ) | ( n7176 & ~n7367 ) | ( n7366 & ~n7367 ) ;
  assign n7369 = n7221 ^ n7089 ^ x90 ;
  assign n7370 = n7258 ^ n7089 ^ 1'b0 ;
  assign n7371 = ( n7089 & n7369 ) | ( n7089 & ~n7370 ) | ( n7369 & ~n7370 ) ;
  assign n7372 = n7218 ^ n7092 ^ x89 ;
  assign n7373 = n7258 ^ n7092 ^ 1'b0 ;
  assign n7374 = ( n7092 & n7372 ) | ( n7092 & ~n7373 ) | ( n7372 & ~n7373 ) ;
  assign n7375 = n7217 ^ n7067 ^ x88 ;
  assign n7376 = n7258 ^ n7067 ^ 1'b0 ;
  assign n7377 = ( n7067 & n7375 ) | ( n7067 & ~n7376 ) | ( n7375 & ~n7376 ) ;
  assign n7378 = n7215 ^ n7098 ^ x86 ;
  assign n7379 = n7258 ^ n7098 ^ 1'b0 ;
  assign n7380 = ( n7098 & n7378 ) | ( n7098 & ~n7379 ) | ( n7378 & ~n7379 ) ;
  assign n7381 = ~x9 & x64 ;
  assign n7382 = x64 & n7258 ;
  assign n7383 = n7382 ^ x64 ^ x10 ;
  assign n7384 = n7383 ^ n7381 ^ x65 ;
  assign n7385 = ( x65 & n7381 ) | ( x65 & n7384 ) | ( n7381 & n7384 ) ;
  assign n7386 = n7385 ^ n7284 ^ x66 ;
  assign n7387 = ( x66 & n7385 ) | ( x66 & n7386 ) | ( n7385 & n7386 ) ;
  assign n7388 = ( x67 & ~n7285 ) | ( x67 & n7387 ) | ( ~n7285 & n7387 ) ;
  assign n7389 = ( x68 & ~n7338 ) | ( x68 & n7388 ) | ( ~n7338 & n7388 ) ;
  assign n7390 = ( x69 & ~n7335 ) | ( x69 & n7389 ) | ( ~n7335 & n7389 ) ;
  assign n7391 = ( x70 & ~n7272 ) | ( x70 & n7390 ) | ( ~n7272 & n7390 ) ;
  assign n7392 = ( x71 & ~n7332 ) | ( x71 & n7391 ) | ( ~n7332 & n7391 ) ;
  assign n7393 = ( x72 & ~n7329 ) | ( x72 & n7392 ) | ( ~n7329 & n7392 ) ;
  assign n7394 = ( x73 & ~n7326 ) | ( x73 & n7393 ) | ( ~n7326 & n7393 ) ;
  assign n7395 = ( x74 & ~n7323 ) | ( x74 & n7394 ) | ( ~n7323 & n7394 ) ;
  assign n7396 = ( x75 & ~n7320 ) | ( x75 & n7395 ) | ( ~n7320 & n7395 ) ;
  assign n7397 = ( x76 & ~n7265 ) | ( x76 & n7396 ) | ( ~n7265 & n7396 ) ;
  assign n7398 = ( x77 & ~n7317 ) | ( x77 & n7397 ) | ( ~n7317 & n7397 ) ;
  assign n7399 = ( x78 & ~n7314 ) | ( x78 & n7398 ) | ( ~n7314 & n7398 ) ;
  assign n7400 = n7398 ^ n7314 ^ x78 ;
  assign n7401 = ( x79 & ~n7311 ) | ( x79 & n7399 ) | ( ~n7311 & n7399 ) ;
  assign n7402 = ( x80 & ~n7278 ) | ( x80 & n7401 ) | ( ~n7278 & n7401 ) ;
  assign n7403 = ( x81 & ~n7308 ) | ( x81 & n7402 ) | ( ~n7308 & n7402 ) ;
  assign n7404 = ( x82 & ~n7305 ) | ( x82 & n7403 ) | ( ~n7305 & n7403 ) ;
  assign n7405 = ( x83 & ~n7273 ) | ( x83 & n7404 ) | ( ~n7273 & n7404 ) ;
  assign n7406 = ( x84 & ~n7276 ) | ( x84 & n7405 ) | ( ~n7276 & n7405 ) ;
  assign n7407 = ( x85 & ~n7302 ) | ( x85 & n7406 ) | ( ~n7302 & n7406 ) ;
  assign n7408 = ( x86 & ~n7299 ) | ( x86 & n7407 ) | ( ~n7299 & n7407 ) ;
  assign n7409 = n7258 ^ n7155 ^ 1'b0 ;
  assign n7410 = n7236 ^ n7155 ^ x102 ;
  assign n7411 = ( n7155 & ~n7409 ) | ( n7155 & n7410 ) | ( ~n7409 & n7410 ) ;
  assign n7412 = n7258 ^ n7072 ^ 1'b0 ;
  assign n7413 = n7258 ^ n7064 ^ 1'b0 ;
  assign n7414 = n7235 ^ n7064 ^ x101 ;
  assign n7415 = ( n7064 & ~n7413 ) | ( n7064 & n7414 ) | ( ~n7413 & n7414 ) ;
  assign n7416 = n7239 ^ n7072 ^ x105 ;
  assign n7417 = n7258 ^ n7158 ^ 1'b0 ;
  assign n7418 = ( n7072 & ~n7412 ) | ( n7072 & n7416 ) | ( ~n7412 & n7416 ) ;
  assign n7419 = ( x87 & ~n7380 ) | ( x87 & n7408 ) | ( ~n7380 & n7408 ) ;
  assign n7420 = ( x88 & ~n7281 ) | ( x88 & n7419 ) | ( ~n7281 & n7419 ) ;
  assign n7421 = n7419 ^ n7281 ^ x88 ;
  assign n7422 = n7258 ^ n7047 ^ 1'b0 ;
  assign n7423 = n7234 ^ n7158 ^ x100 ;
  assign n7424 = n7232 ^ n7047 ^ x98 ;
  assign n7425 = ( n7158 & ~n7417 ) | ( n7158 & n7423 ) | ( ~n7417 & n7423 ) ;
  assign n7426 = n7237 ^ n7152 ^ x103 ;
  assign n7427 = ( x89 & ~n7377 ) | ( x89 & n7420 ) | ( ~n7377 & n7420 ) ;
  assign n7428 = ( x90 & ~n7374 ) | ( x90 & n7427 ) | ( ~n7374 & n7427 ) ;
  assign n7429 = n7258 ^ n7149 ^ 1'b0 ;
  assign n7430 = n7388 ^ n7338 ^ x68 ;
  assign n7431 = ( n7047 & ~n7422 ) | ( n7047 & n7424 ) | ( ~n7422 & n7424 ) ;
  assign n7432 = ( x91 & ~n7371 ) | ( x91 & n7428 ) | ( ~n7371 & n7428 ) ;
  assign n7433 = n7427 ^ n7374 ^ x90 ;
  assign n7434 = n7241 ^ n7149 ^ x106 ;
  assign n7435 = n7238 ^ n7077 ^ x104 ;
  assign n7436 = n7395 ^ n7320 ^ x75 ;
  assign n7437 = n7393 ^ n7326 ^ x73 ;
  assign n7438 = n7258 ^ n7152 ^ 1'b0 ;
  assign n7439 = ( n7152 & n7426 ) | ( n7152 & ~n7438 ) | ( n7426 & ~n7438 ) ;
  assign n7440 = n7233 ^ n7161 ^ x99 ;
  assign n7441 = n7258 ^ n7077 ^ 1'b0 ;
  assign n7442 = n7258 ^ n7161 ^ 1'b0 ;
  assign n7443 = ( n7161 & n7440 ) | ( n7161 & ~n7442 ) | ( n7440 & ~n7442 ) ;
  assign n7444 = ( x92 & ~n7368 ) | ( x92 & n7432 ) | ( ~n7368 & n7432 ) ;
  assign n7445 = ( x93 & ~n7287 ) | ( x93 & n7444 ) | ( ~n7287 & n7444 ) ;
  assign n7446 = ( n7149 & ~n7429 ) | ( n7149 & n7434 ) | ( ~n7429 & n7434 ) ;
  assign n7447 = ( x94 & ~n7365 ) | ( x94 & n7445 ) | ( ~n7365 & n7445 ) ;
  assign n7448 = ( x95 & ~n7362 ) | ( x95 & n7447 ) | ( ~n7362 & n7447 ) ;
  assign n7449 = n7447 ^ n7362 ^ x95 ;
  assign n7450 = n7404 ^ n7273 ^ x83 ;
  assign n7451 = n7391 ^ n7332 ^ x71 ;
  assign n7452 = ( n7077 & n7435 ) | ( n7077 & ~n7441 ) | ( n7435 & ~n7441 ) ;
  assign n7453 = n7448 ^ n7266 ^ x96 ;
  assign n7454 = n7445 ^ n7365 ^ x94 ;
  assign n7455 = ( x96 & ~n7266 ) | ( x96 & n7448 ) | ( ~n7266 & n7448 ) ;
  assign n7456 = n7396 ^ n7265 ^ x76 ;
  assign n7457 = ( x97 & ~n7280 ) | ( x97 & n7455 ) | ( ~n7280 & n7455 ) ;
  assign n7458 = n7392 ^ n7329 ^ x72 ;
  assign n7459 = ( x98 & ~n7359 ) | ( x98 & n7457 ) | ( ~n7359 & n7457 ) ;
  assign n7460 = ( x99 & ~n7431 ) | ( x99 & n7459 ) | ( ~n7431 & n7459 ) ;
  assign n7461 = ( x100 & ~n7443 ) | ( x100 & n7460 ) | ( ~n7443 & n7460 ) ;
  assign n7462 = ( x101 & ~n7425 ) | ( x101 & n7461 ) | ( ~n7425 & n7461 ) ;
  assign n7463 = ( x102 & ~n7415 ) | ( x102 & n7462 ) | ( ~n7415 & n7462 ) ;
  assign n7464 = ( x103 & ~n7411 ) | ( x103 & n7463 ) | ( ~n7411 & n7463 ) ;
  assign n7465 = ( x104 & ~n7439 ) | ( x104 & n7464 ) | ( ~n7439 & n7464 ) ;
  assign n7466 = ( x105 & ~n7452 ) | ( x105 & n7465 ) | ( ~n7452 & n7465 ) ;
  assign n7467 = ( x106 & ~n7418 ) | ( x106 & n7466 ) | ( ~n7418 & n7466 ) ;
  assign n7468 = ( x107 & ~n7446 ) | ( x107 & n7467 ) | ( ~n7446 & n7467 ) ;
  assign n7469 = ( x108 & ~n7356 ) | ( x108 & n7468 ) | ( ~n7356 & n7468 ) ;
  assign n7470 = ( x109 & ~n7353 ) | ( x109 & n7469 ) | ( ~n7353 & n7469 ) ;
  assign n7471 = ( x110 & ~n7350 ) | ( x110 & n7470 ) | ( ~n7350 & n7470 ) ;
  assign n7472 = ( x111 & ~n7283 ) | ( x111 & n7471 ) | ( ~n7283 & n7471 ) ;
  assign n7473 = ( x112 & ~n7347 ) | ( x112 & n7472 ) | ( ~n7347 & n7472 ) ;
  assign n7474 = ( x113 & ~n7344 ) | ( x113 & n7473 ) | ( ~n7344 & n7473 ) ;
  assign n7475 = ( x114 & ~n7341 ) | ( x114 & n7474 ) | ( ~n7341 & n7474 ) ;
  assign n7476 = ( x115 & ~n7296 ) | ( x115 & n7475 ) | ( ~n7296 & n7475 ) ;
  assign n7477 = ( x116 & ~n7293 ) | ( x116 & n7476 ) | ( ~n7293 & n7476 ) ;
  assign n7478 = ( x117 & ~n7290 ) | ( x117 & n7477 ) | ( ~n7290 & n7477 ) ;
  assign n7479 = ( x118 & ~n7262 ) | ( x118 & n7478 ) | ( ~n7262 & n7478 ) ;
  assign n7480 = n1296 | n7479 ;
  assign n7481 = n7480 ^ n7453 ^ 1'b0 ;
  assign n7482 = ( n7266 & n7453 ) | ( n7266 & n7481 ) | ( n7453 & n7481 ) ;
  assign n7483 = n7480 ^ n7449 ^ 1'b0 ;
  assign n7484 = ( n7362 & n7449 ) | ( n7362 & n7483 ) | ( n7449 & n7483 ) ;
  assign n7485 = n7480 ^ n7454 ^ 1'b0 ;
  assign n7486 = ( n7365 & n7454 ) | ( n7365 & n7485 ) | ( n7454 & n7485 ) ;
  assign n7487 = n7480 ^ n7421 ^ 1'b0 ;
  assign n7488 = n7480 ^ n7450 ^ 1'b0 ;
  assign n7489 = ( n7273 & n7450 ) | ( n7273 & n7488 ) | ( n7450 & n7488 ) ;
  assign n7490 = n7480 ^ n7400 ^ 1'b0 ;
  assign n7491 = ( n7314 & n7400 ) | ( n7314 & n7490 ) | ( n7400 & n7490 ) ;
  assign n7492 = n7480 ^ n7456 ^ 1'b0 ;
  assign n7493 = ( n7265 & n7456 ) | ( n7265 & n7492 ) | ( n7456 & n7492 ) ;
  assign n7494 = n7480 ^ n7436 ^ 1'b0 ;
  assign n7495 = ( n7320 & n7436 ) | ( n7320 & n7494 ) | ( n7436 & n7494 ) ;
  assign n7496 = n7480 ^ n7437 ^ 1'b0 ;
  assign n7497 = ( n7326 & n7437 ) | ( n7326 & n7496 ) | ( n7437 & n7496 ) ;
  assign n7498 = n7480 ^ n7458 ^ 1'b0 ;
  assign n7499 = ( n7281 & n7421 ) | ( n7281 & n7487 ) | ( n7421 & n7487 ) ;
  assign n7500 = ( n7329 & n7458 ) | ( n7329 & n7498 ) | ( n7458 & n7498 ) ;
  assign n7501 = n7480 ^ n7451 ^ 1'b0 ;
  assign n7502 = ( n7332 & n7451 ) | ( n7332 & n7501 ) | ( n7451 & n7501 ) ;
  assign n7503 = n7480 ^ n7430 ^ 1'b0 ;
  assign n7504 = ( n7338 & n7430 ) | ( n7338 & n7503 ) | ( n7430 & n7503 ) ;
  assign n7505 = n7480 ^ n7284 ^ 1'b0 ;
  assign n7506 = ( n7284 & n7386 ) | ( n7284 & ~n7505 ) | ( n7386 & ~n7505 ) ;
  assign n7507 = n7480 ^ n7383 ^ 1'b0 ;
  assign n7508 = ( n7383 & n7384 ) | ( n7383 & ~n7507 ) | ( n7384 & ~n7507 ) ;
  assign n7509 = n7477 ^ n7290 ^ x117 ;
  assign n7510 = n7509 ^ n7480 ^ 1'b0 ;
  assign n7511 = ( n7290 & n7509 ) | ( n7290 & n7510 ) | ( n7509 & n7510 ) ;
  assign n7512 = n7476 ^ n7293 ^ x116 ;
  assign n7513 = n7512 ^ n7480 ^ 1'b0 ;
  assign n7514 = ( n7293 & n7512 ) | ( n7293 & n7513 ) | ( n7512 & n7513 ) ;
  assign n7515 = n7475 ^ n7296 ^ x115 ;
  assign n7516 = n7515 ^ n7480 ^ 1'b0 ;
  assign n7517 = ( n7296 & n7515 ) | ( n7296 & n7516 ) | ( n7515 & n7516 ) ;
  assign n7518 = n7474 ^ n7341 ^ x114 ;
  assign n7519 = n7518 ^ n7480 ^ 1'b0 ;
  assign n7520 = ( n7341 & n7518 ) | ( n7341 & n7519 ) | ( n7518 & n7519 ) ;
  assign n7521 = n7473 ^ n7344 ^ x113 ;
  assign n7522 = n7521 ^ n7480 ^ 1'b0 ;
  assign n7523 = ( n7344 & n7521 ) | ( n7344 & n7522 ) | ( n7521 & n7522 ) ;
  assign n7524 = n7472 ^ n7347 ^ x112 ;
  assign n7525 = n7524 ^ n7480 ^ 1'b0 ;
  assign n7526 = ( n7347 & n7524 ) | ( n7347 & n7525 ) | ( n7524 & n7525 ) ;
  assign n7527 = n7471 ^ n7283 ^ x111 ;
  assign n7528 = n7527 ^ n7480 ^ 1'b0 ;
  assign n7529 = ( n7283 & n7527 ) | ( n7283 & n7528 ) | ( n7527 & n7528 ) ;
  assign n7530 = n7470 ^ n7350 ^ x110 ;
  assign n7531 = n7530 ^ n7480 ^ 1'b0 ;
  assign n7532 = ( n7350 & n7530 ) | ( n7350 & n7531 ) | ( n7530 & n7531 ) ;
  assign n7533 = n7469 ^ n7353 ^ x109 ;
  assign n7534 = n7533 ^ n7480 ^ 1'b0 ;
  assign n7535 = ( n7353 & n7533 ) | ( n7353 & n7534 ) | ( n7533 & n7534 ) ;
  assign n7536 = n7468 ^ n7356 ^ x108 ;
  assign n7537 = n7536 ^ n7480 ^ 1'b0 ;
  assign n7538 = ( n7356 & n7536 ) | ( n7356 & n7537 ) | ( n7536 & n7537 ) ;
  assign n7539 = n7467 ^ n7446 ^ x107 ;
  assign n7540 = n7539 ^ n7480 ^ 1'b0 ;
  assign n7541 = ( n7446 & n7539 ) | ( n7446 & n7540 ) | ( n7539 & n7540 ) ;
  assign n7542 = n7466 ^ n7418 ^ x106 ;
  assign n7543 = n7542 ^ n7480 ^ 1'b0 ;
  assign n7544 = ( n7418 & n7542 ) | ( n7418 & n7543 ) | ( n7542 & n7543 ) ;
  assign n7545 = n7459 ^ n7431 ^ x99 ;
  assign n7546 = n7545 ^ n7480 ^ 1'b0 ;
  assign n7547 = ( n7431 & n7545 ) | ( n7431 & n7546 ) | ( n7545 & n7546 ) ;
  assign n7548 = n7457 ^ n7359 ^ x98 ;
  assign n7549 = n7548 ^ n7480 ^ 1'b0 ;
  assign n7550 = ( n7359 & n7548 ) | ( n7359 & n7549 ) | ( n7548 & n7549 ) ;
  assign n7551 = n7480 ^ n7433 ^ 1'b0 ;
  assign n7552 = ( n7374 & n7433 ) | ( n7374 & n7551 ) | ( n7433 & n7551 ) ;
  assign n7553 = n7465 ^ n7452 ^ x105 ;
  assign n7554 = n7553 ^ n7480 ^ 1'b0 ;
  assign n7555 = ( n7452 & n7553 ) | ( n7452 & n7554 ) | ( n7553 & n7554 ) ;
  assign n7556 = n7464 ^ n7439 ^ x104 ;
  assign n7557 = n7556 ^ n7480 ^ 1'b0 ;
  assign n7558 = ( n7439 & n7556 ) | ( n7439 & n7557 ) | ( n7556 & n7557 ) ;
  assign n7559 = n7463 ^ n7411 ^ x103 ;
  assign n7560 = n7559 ^ n7480 ^ 1'b0 ;
  assign n7561 = ( n7411 & n7559 ) | ( n7411 & n7560 ) | ( n7559 & n7560 ) ;
  assign n7562 = n7462 ^ n7415 ^ x102 ;
  assign n7563 = n7562 ^ n7480 ^ 1'b0 ;
  assign n7564 = ( n7415 & n7562 ) | ( n7415 & n7563 ) | ( n7562 & n7563 ) ;
  assign n7565 = n7461 ^ n7425 ^ x101 ;
  assign n7566 = n7565 ^ n7480 ^ 1'b0 ;
  assign n7567 = ( n7425 & n7565 ) | ( n7425 & n7566 ) | ( n7565 & n7566 ) ;
  assign n7568 = n7460 ^ n7443 ^ x100 ;
  assign n7569 = n7568 ^ n7480 ^ 1'b0 ;
  assign n7570 = ( n7443 & n7568 ) | ( n7443 & n7569 ) | ( n7568 & n7569 ) ;
  assign n7571 = n7455 ^ n7280 ^ x97 ;
  assign n7572 = n7571 ^ n7480 ^ 1'b0 ;
  assign n7573 = ( n7280 & n7571 ) | ( n7280 & n7572 ) | ( n7571 & n7572 ) ;
  assign n7574 = n7444 ^ n7287 ^ x93 ;
  assign n7575 = n7574 ^ n7480 ^ 1'b0 ;
  assign n7576 = ( n7287 & n7574 ) | ( n7287 & n7575 ) | ( n7574 & n7575 ) ;
  assign n7577 = n7432 ^ n7368 ^ x92 ;
  assign n7578 = n7577 ^ n7480 ^ 1'b0 ;
  assign n7579 = ( n7368 & n7577 ) | ( n7368 & n7578 ) | ( n7577 & n7578 ) ;
  assign n7580 = n7428 ^ n7371 ^ x91 ;
  assign n7581 = n7580 ^ n7480 ^ 1'b0 ;
  assign n7582 = ( n7371 & n7580 ) | ( n7371 & n7581 ) | ( n7580 & n7581 ) ;
  assign n7583 = n7420 ^ n7377 ^ x89 ;
  assign n7584 = n7583 ^ n7480 ^ 1'b0 ;
  assign n7585 = ( n7377 & n7583 ) | ( n7377 & n7584 ) | ( n7583 & n7584 ) ;
  assign n7586 = n7408 ^ n7380 ^ x87 ;
  assign n7587 = n7586 ^ n7480 ^ 1'b0 ;
  assign n7588 = ( n7380 & n7586 ) | ( n7380 & n7587 ) | ( n7586 & n7587 ) ;
  assign n7589 = n7407 ^ n7299 ^ x86 ;
  assign n7590 = n7589 ^ n7480 ^ 1'b0 ;
  assign n7591 = ( n7299 & n7589 ) | ( n7299 & n7590 ) | ( n7589 & n7590 ) ;
  assign n7592 = n7406 ^ n7302 ^ x85 ;
  assign n7593 = n7592 ^ n7480 ^ 1'b0 ;
  assign n7594 = ( n7302 & n7592 ) | ( n7302 & n7593 ) | ( n7592 & n7593 ) ;
  assign n7595 = n7405 ^ n7276 ^ x84 ;
  assign n7596 = n7595 ^ n7480 ^ 1'b0 ;
  assign n7597 = ( n7276 & n7595 ) | ( n7276 & n7596 ) | ( n7595 & n7596 ) ;
  assign n7598 = n7403 ^ n7305 ^ x82 ;
  assign n7599 = n7598 ^ n7480 ^ 1'b0 ;
  assign n7600 = ( n7305 & n7598 ) | ( n7305 & n7599 ) | ( n7598 & n7599 ) ;
  assign n7601 = n7402 ^ n7308 ^ x81 ;
  assign n7602 = n7601 ^ n7480 ^ 1'b0 ;
  assign n7603 = ( n7308 & n7601 ) | ( n7308 & n7602 ) | ( n7601 & n7602 ) ;
  assign n7604 = n7401 ^ n7278 ^ x80 ;
  assign n7605 = n7604 ^ n7480 ^ 1'b0 ;
  assign n7606 = ( n7278 & n7604 ) | ( n7278 & n7605 ) | ( n7604 & n7605 ) ;
  assign n7607 = n7399 ^ n7311 ^ x79 ;
  assign n7608 = n7607 ^ n7480 ^ 1'b0 ;
  assign n7609 = ( n7311 & n7607 ) | ( n7311 & n7608 ) | ( n7607 & n7608 ) ;
  assign n7610 = n7397 ^ n7317 ^ x77 ;
  assign n7611 = n7610 ^ n7480 ^ 1'b0 ;
  assign n7612 = ( n7317 & n7610 ) | ( n7317 & n7611 ) | ( n7610 & n7611 ) ;
  assign n7613 = n7394 ^ n7323 ^ x74 ;
  assign n7614 = n7613 ^ n7480 ^ 1'b0 ;
  assign n7615 = ( n7323 & n7613 ) | ( n7323 & n7614 ) | ( n7613 & n7614 ) ;
  assign n7616 = n7390 ^ n7272 ^ x70 ;
  assign n7617 = n7616 ^ n7480 ^ 1'b0 ;
  assign n7618 = ( n7272 & n7616 ) | ( n7272 & n7617 ) | ( n7616 & n7617 ) ;
  assign n7619 = n7389 ^ n7335 ^ x69 ;
  assign n7620 = n7619 ^ n7480 ^ 1'b0 ;
  assign n7621 = ( n7335 & n7619 ) | ( n7335 & n7620 ) | ( n7619 & n7620 ) ;
  assign n7622 = n7387 ^ n7285 ^ x67 ;
  assign n7623 = n7622 ^ n7480 ^ 1'b0 ;
  assign n7624 = ( n7285 & n7622 ) | ( n7285 & n7623 ) | ( n7622 & n7623 ) ;
  assign n7625 = n7478 ^ n7262 ^ x118 ;
  assign n7626 = n7625 ^ n7480 ^ 1'b0 ;
  assign n7627 = ( n7262 & n7625 ) | ( n7262 & n7626 ) | ( n7625 & n7626 ) ;
  assign n7628 = n1296 & n7262 ;
  assign n7629 = ~x8 & x64 ;
  assign n7630 = ( x64 & x119 ) | ( x64 & ~n163 ) | ( x119 & ~n163 ) ;
  assign n7631 = ~x119 & n7630 ;
  assign n7632 = ~n1296 & n7381 ;
  assign n7633 = n7479 | n7632 ;
  assign n7634 = ( x9 & ~n7479 ) | ( x9 & n7633 ) | ( ~n7479 & n7633 ) ;
  assign n7635 = ~n7631 & n7634 ;
  assign n7636 = ( n7633 & n7634 ) | ( n7633 & n7635 ) | ( n7634 & n7635 ) ;
  assign n7637 = n7636 ^ n7629 ^ x65 ;
  assign n7638 = ( x65 & n7629 ) | ( x65 & n7637 ) | ( n7629 & n7637 ) ;
  assign n7639 = n7638 ^ n7508 ^ x66 ;
  assign n7640 = ( x66 & n7638 ) | ( x66 & n7639 ) | ( n7638 & n7639 ) ;
  assign n7641 = ( x67 & ~n7506 ) | ( x67 & n7640 ) | ( ~n7506 & n7640 ) ;
  assign n7642 = ( x68 & ~n7624 ) | ( x68 & n7641 ) | ( ~n7624 & n7641 ) ;
  assign n7643 = n7642 ^ n7504 ^ x69 ;
  assign n7644 = n7640 ^ n7506 ^ x67 ;
  assign n7645 = ( x69 & ~n7504 ) | ( x69 & n7642 ) | ( ~n7504 & n7642 ) ;
  assign n7646 = ( x70 & ~n7621 ) | ( x70 & n7645 ) | ( ~n7621 & n7645 ) ;
  assign n7647 = n7645 ^ n7621 ^ x70 ;
  assign n7648 = ( x71 & ~n7618 ) | ( x71 & n7646 ) | ( ~n7618 & n7646 ) ;
  assign n7649 = ( x72 & ~n7502 ) | ( x72 & n7648 ) | ( ~n7502 & n7648 ) ;
  assign n7650 = ( x73 & ~n7500 ) | ( x73 & n7649 ) | ( ~n7500 & n7649 ) ;
  assign n7651 = ( x74 & ~n7497 ) | ( x74 & n7650 ) | ( ~n7497 & n7650 ) ;
  assign n7652 = ( x75 & ~n7615 ) | ( x75 & n7651 ) | ( ~n7615 & n7651 ) ;
  assign n7653 = ( x76 & ~n7495 ) | ( x76 & n7652 ) | ( ~n7495 & n7652 ) ;
  assign n7654 = n7646 ^ n7618 ^ x71 ;
  assign n7655 = ( x77 & ~n7493 ) | ( x77 & n7653 ) | ( ~n7493 & n7653 ) ;
  assign n7656 = n7655 ^ n7612 ^ x78 ;
  assign n7657 = ( x78 & ~n7612 ) | ( x78 & n7655 ) | ( ~n7612 & n7655 ) ;
  assign n7658 = n7649 ^ n7500 ^ x73 ;
  assign n7659 = n7641 ^ n7624 ^ x68 ;
  assign n7660 = n7653 ^ n7493 ^ x77 ;
  assign n7661 = n7648 ^ n7502 ^ x72 ;
  assign n7662 = ( x79 & ~n7491 ) | ( x79 & n7657 ) | ( ~n7491 & n7657 ) ;
  assign n7663 = ( x80 & ~n7609 ) | ( x80 & n7662 ) | ( ~n7609 & n7662 ) ;
  assign n7664 = ( x81 & ~n7606 ) | ( x81 & n7663 ) | ( ~n7606 & n7663 ) ;
  assign n7665 = ( x82 & ~n7603 ) | ( x82 & n7664 ) | ( ~n7603 & n7664 ) ;
  assign n7666 = ( x83 & ~n7600 ) | ( x83 & n7665 ) | ( ~n7600 & n7665 ) ;
  assign n7667 = n7666 ^ n7489 ^ x84 ;
  assign n7668 = n7663 ^ n7606 ^ x81 ;
  assign n7669 = n7664 ^ n7603 ^ x82 ;
  assign n7670 = n7665 ^ n7600 ^ x83 ;
  assign n7671 = n7650 ^ n7497 ^ x74 ;
  assign n7672 = ( x84 & ~n7489 ) | ( x84 & n7666 ) | ( ~n7489 & n7666 ) ;
  assign n7673 = ( x85 & ~n7597 ) | ( x85 & n7672 ) | ( ~n7597 & n7672 ) ;
  assign n7674 = ( x86 & ~n7594 ) | ( x86 & n7673 ) | ( ~n7594 & n7673 ) ;
  assign n7675 = ( x87 & ~n7591 ) | ( x87 & n7674 ) | ( ~n7591 & n7674 ) ;
  assign n7676 = n7675 ^ n7588 ^ x88 ;
  assign n7677 = n7651 ^ n7615 ^ x75 ;
  assign n7678 = n7662 ^ n7609 ^ x80 ;
  assign n7679 = n7673 ^ n7594 ^ x86 ;
  assign n7680 = n7674 ^ n7591 ^ x87 ;
  assign n7681 = n7652 ^ n7495 ^ x76 ;
  assign n7682 = ( x88 & ~n7588 ) | ( x88 & n7675 ) | ( ~n7588 & n7675 ) ;
  assign n7683 = ( x89 & ~n7499 ) | ( x89 & n7682 ) | ( ~n7499 & n7682 ) ;
  assign n7684 = n7683 ^ n7585 ^ x90 ;
  assign n7685 = n7657 ^ n7491 ^ x79 ;
  assign n7686 = ( x90 & ~n7585 ) | ( x90 & n7683 ) | ( ~n7585 & n7683 ) ;
  assign n7687 = ( x91 & ~n7552 ) | ( x91 & n7686 ) | ( ~n7552 & n7686 ) ;
  assign n7688 = ( x92 & ~n7582 ) | ( x92 & n7687 ) | ( ~n7582 & n7687 ) ;
  assign n7689 = n7687 ^ n7582 ^ x92 ;
  assign n7690 = n7672 ^ n7597 ^ x85 ;
  assign n7691 = n7686 ^ n7552 ^ x91 ;
  assign n7692 = n7682 ^ n7499 ^ x89 ;
  assign n7693 = ( x93 & ~n7579 ) | ( x93 & n7688 ) | ( ~n7579 & n7688 ) ;
  assign n7694 = ( x94 & ~n7576 ) | ( x94 & n7693 ) | ( ~n7576 & n7693 ) ;
  assign n7695 = ( x95 & ~n7486 ) | ( x95 & n7694 ) | ( ~n7486 & n7694 ) ;
  assign n7696 = ( x96 & ~n7484 ) | ( x96 & n7695 ) | ( ~n7484 & n7695 ) ;
  assign n7697 = ( x97 & ~n7482 ) | ( x97 & n7696 ) | ( ~n7482 & n7696 ) ;
  assign n7698 = ( x98 & ~n7573 ) | ( x98 & n7697 ) | ( ~n7573 & n7697 ) ;
  assign n7699 = ( x99 & ~n7550 ) | ( x99 & n7698 ) | ( ~n7550 & n7698 ) ;
  assign n7700 = ( x100 & ~n7547 ) | ( x100 & n7699 ) | ( ~n7547 & n7699 ) ;
  assign n7701 = ( x101 & ~n7570 ) | ( x101 & n7700 ) | ( ~n7570 & n7700 ) ;
  assign n7702 = ( x102 & ~n7567 ) | ( x102 & n7701 ) | ( ~n7567 & n7701 ) ;
  assign n7703 = ( x103 & ~n7564 ) | ( x103 & n7702 ) | ( ~n7564 & n7702 ) ;
  assign n7704 = ( x104 & ~n7561 ) | ( x104 & n7703 ) | ( ~n7561 & n7703 ) ;
  assign n7705 = ( x105 & ~n7558 ) | ( x105 & n7704 ) | ( ~n7558 & n7704 ) ;
  assign n7706 = ( x106 & ~n7555 ) | ( x106 & n7705 ) | ( ~n7555 & n7705 ) ;
  assign n7707 = ( x107 & ~n7544 ) | ( x107 & n7706 ) | ( ~n7544 & n7706 ) ;
  assign n7708 = ( x108 & ~n7541 ) | ( x108 & n7707 ) | ( ~n7541 & n7707 ) ;
  assign n7709 = ( x109 & ~n7538 ) | ( x109 & n7708 ) | ( ~n7538 & n7708 ) ;
  assign n7710 = ( x110 & ~n7535 ) | ( x110 & n7709 ) | ( ~n7535 & n7709 ) ;
  assign n7711 = ( x111 & ~n7532 ) | ( x111 & n7710 ) | ( ~n7532 & n7710 ) ;
  assign n7712 = ( x119 & n163 ) | ( x119 & ~n7627 ) | ( n163 & ~n7627 ) ;
  assign n7713 = ( x112 & ~n7529 ) | ( x112 & n7711 ) | ( ~n7529 & n7711 ) ;
  assign n7714 = ( x113 & ~n7526 ) | ( x113 & n7713 ) | ( ~n7526 & n7713 ) ;
  assign n7715 = ( x114 & ~n7523 ) | ( x114 & n7714 ) | ( ~n7523 & n7714 ) ;
  assign n7716 = ( x115 & ~n7520 ) | ( x115 & n7715 ) | ( ~n7520 & n7715 ) ;
  assign n7717 = ( x116 & ~n7517 ) | ( x116 & n7716 ) | ( ~n7517 & n7716 ) ;
  assign n7718 = ( x117 & ~n7514 ) | ( x117 & n7717 ) | ( ~n7514 & n7717 ) ;
  assign n7719 = ( x118 & ~n7511 ) | ( x118 & n7718 ) | ( ~n7511 & n7718 ) ;
  assign n7720 = ( ~x119 & n7627 ) | ( ~x119 & n7719 ) | ( n7627 & n7719 ) ;
  assign n7721 = n7712 | n7720 ;
  assign n7722 = n1296 & n7627 ;
  assign n7723 = ( ~n7627 & n7721 ) | ( ~n7627 & n7722 ) | ( n7721 & n7722 ) ;
  assign n7724 = n7719 ^ n7627 ^ x119 ;
  assign n7725 = ~n7723 & n7724 ;
  assign n7726 = n7723 ^ n7600 ^ 1'b0 ;
  assign n7727 = ( n7600 & n7670 ) | ( n7600 & ~n7726 ) | ( n7670 & ~n7726 ) ;
  assign n7728 = n7723 ^ n7497 ^ 1'b0 ;
  assign n7729 = ( n7497 & n7671 ) | ( n7497 & ~n7728 ) | ( n7671 & ~n7728 ) ;
  assign n7730 = n7723 ^ n7585 ^ 1'b0 ;
  assign n7731 = n7723 ^ n7624 ^ 1'b0 ;
  assign n7732 = ( n7624 & n7659 ) | ( n7624 & ~n7731 ) | ( n7659 & ~n7731 ) ;
  assign n7733 = n7723 ^ n7495 ^ 1'b0 ;
  assign n7734 = n7628 & ~n7721 ;
  assign n7735 = n7723 ^ n7582 ^ 1'b0 ;
  assign n7736 = n7723 ^ n7552 ^ 1'b0 ;
  assign n7737 = ( n7495 & n7681 ) | ( n7495 & ~n7733 ) | ( n7681 & ~n7733 ) ;
  assign n7738 = ( n7628 & n7725 ) | ( n7628 & ~n7734 ) | ( n7725 & ~n7734 ) ;
  assign n7739 = ( n7552 & n7691 ) | ( n7552 & ~n7736 ) | ( n7691 & ~n7736 ) ;
  assign n7740 = ( n7582 & n7689 ) | ( n7582 & ~n7735 ) | ( n7689 & ~n7735 ) ;
  assign n7741 = ( n7585 & n7684 ) | ( n7585 & ~n7730 ) | ( n7684 & ~n7730 ) ;
  assign n7742 = n7723 ^ n7499 ^ 1'b0 ;
  assign n7743 = ( n7499 & n7692 ) | ( n7499 & ~n7742 ) | ( n7692 & ~n7742 ) ;
  assign n7744 = n7723 ^ n7588 ^ 1'b0 ;
  assign n7745 = ( n7588 & n7676 ) | ( n7588 & ~n7744 ) | ( n7676 & ~n7744 ) ;
  assign n7746 = n7723 ^ n7591 ^ 1'b0 ;
  assign n7747 = ( n7591 & n7680 ) | ( n7591 & ~n7746 ) | ( n7680 & ~n7746 ) ;
  assign n7748 = n7723 ^ n7594 ^ 1'b0 ;
  assign n7749 = ( n7594 & n7679 ) | ( n7594 & ~n7748 ) | ( n7679 & ~n7748 ) ;
  assign n7750 = n7723 ^ n7597 ^ 1'b0 ;
  assign n7751 = ( n7597 & n7690 ) | ( n7597 & ~n7750 ) | ( n7690 & ~n7750 ) ;
  assign n7752 = n7723 ^ n7489 ^ 1'b0 ;
  assign n7753 = ( n7489 & n7667 ) | ( n7489 & ~n7752 ) | ( n7667 & ~n7752 ) ;
  assign n7754 = n7723 ^ n7603 ^ 1'b0 ;
  assign n7755 = ( n7603 & n7669 ) | ( n7603 & ~n7754 ) | ( n7669 & ~n7754 ) ;
  assign n7756 = n7723 ^ n7606 ^ 1'b0 ;
  assign n7757 = ( n7606 & n7668 ) | ( n7606 & ~n7756 ) | ( n7668 & ~n7756 ) ;
  assign n7758 = n7723 ^ n7609 ^ 1'b0 ;
  assign n7759 = ( n7609 & n7678 ) | ( n7609 & ~n7758 ) | ( n7678 & ~n7758 ) ;
  assign n7760 = n7723 ^ n7491 ^ 1'b0 ;
  assign n7761 = ( n7491 & n7685 ) | ( n7491 & ~n7760 ) | ( n7685 & ~n7760 ) ;
  assign n7762 = n7723 ^ n7612 ^ 1'b0 ;
  assign n7763 = ( n7612 & n7656 ) | ( n7612 & ~n7762 ) | ( n7656 & ~n7762 ) ;
  assign n7764 = n7723 ^ n7493 ^ 1'b0 ;
  assign n7765 = ( n7493 & n7660 ) | ( n7493 & ~n7764 ) | ( n7660 & ~n7764 ) ;
  assign n7766 = n7723 ^ n7615 ^ 1'b0 ;
  assign n7767 = ( n7615 & n7677 ) | ( n7615 & ~n7766 ) | ( n7677 & ~n7766 ) ;
  assign n7768 = n7723 ^ n7500 ^ 1'b0 ;
  assign n7769 = ( n7500 & n7658 ) | ( n7500 & ~n7768 ) | ( n7658 & ~n7768 ) ;
  assign n7770 = n7723 ^ n7502 ^ 1'b0 ;
  assign n7771 = ( n7502 & n7661 ) | ( n7502 & ~n7770 ) | ( n7661 & ~n7770 ) ;
  assign n7772 = n7723 ^ n7618 ^ 1'b0 ;
  assign n7773 = ( n7618 & n7654 ) | ( n7618 & ~n7772 ) | ( n7654 & ~n7772 ) ;
  assign n7774 = n7723 ^ n7621 ^ 1'b0 ;
  assign n7775 = ( n7621 & n7647 ) | ( n7621 & ~n7774 ) | ( n7647 & ~n7774 ) ;
  assign n7776 = n7723 ^ n7504 ^ 1'b0 ;
  assign n7777 = ( n7504 & n7643 ) | ( n7504 & ~n7776 ) | ( n7643 & ~n7776 ) ;
  assign n7778 = n7723 ^ n7506 ^ 1'b0 ;
  assign n7779 = ( n7506 & n7644 ) | ( n7506 & ~n7778 ) | ( n7644 & ~n7778 ) ;
  assign n7780 = n7723 ^ n7639 ^ 1'b0 ;
  assign n7781 = ( n7508 & n7639 ) | ( n7508 & n7780 ) | ( n7639 & n7780 ) ;
  assign n7782 = n7723 ^ n7637 ^ 1'b0 ;
  assign n7783 = ( n7636 & n7637 ) | ( n7636 & n7782 ) | ( n7637 & n7782 ) ;
  assign n7784 = n7718 ^ n7511 ^ x118 ;
  assign n7785 = n7723 ^ n7511 ^ 1'b0 ;
  assign n7786 = ( n7511 & n7784 ) | ( n7511 & ~n7785 ) | ( n7784 & ~n7785 ) ;
  assign n7787 = n7717 ^ n7514 ^ x117 ;
  assign n7788 = n7723 ^ n7514 ^ 1'b0 ;
  assign n7789 = ( n7514 & n7787 ) | ( n7514 & ~n7788 ) | ( n7787 & ~n7788 ) ;
  assign n7790 = n7716 ^ n7517 ^ x116 ;
  assign n7791 = n7723 ^ n7517 ^ 1'b0 ;
  assign n7792 = ( n7517 & n7790 ) | ( n7517 & ~n7791 ) | ( n7790 & ~n7791 ) ;
  assign n7793 = n7715 ^ n7520 ^ x115 ;
  assign n7794 = n7723 ^ n7520 ^ 1'b0 ;
  assign n7795 = ( n7520 & n7793 ) | ( n7520 & ~n7794 ) | ( n7793 & ~n7794 ) ;
  assign n7796 = n7714 ^ n7523 ^ x114 ;
  assign n7797 = n7723 ^ n7523 ^ 1'b0 ;
  assign n7798 = ( n7523 & n7796 ) | ( n7523 & ~n7797 ) | ( n7796 & ~n7797 ) ;
  assign n7799 = n7713 ^ n7526 ^ x113 ;
  assign n7800 = n7723 ^ n7526 ^ 1'b0 ;
  assign n7801 = ( n7526 & n7799 ) | ( n7526 & ~n7800 ) | ( n7799 & ~n7800 ) ;
  assign n7802 = n7711 ^ n7529 ^ x112 ;
  assign n7803 = n7723 ^ n7529 ^ 1'b0 ;
  assign n7804 = ( n7529 & n7802 ) | ( n7529 & ~n7803 ) | ( n7802 & ~n7803 ) ;
  assign n7805 = n7710 ^ n7532 ^ x111 ;
  assign n7806 = n7723 ^ n7532 ^ 1'b0 ;
  assign n7807 = ( n7532 & n7805 ) | ( n7532 & ~n7806 ) | ( n7805 & ~n7806 ) ;
  assign n7808 = n7709 ^ n7535 ^ x110 ;
  assign n7809 = n7723 ^ n7535 ^ 1'b0 ;
  assign n7810 = ( n7535 & n7808 ) | ( n7535 & ~n7809 ) | ( n7808 & ~n7809 ) ;
  assign n7811 = n7708 ^ n7538 ^ x109 ;
  assign n7812 = n7723 ^ n7538 ^ 1'b0 ;
  assign n7813 = ( n7538 & n7811 ) | ( n7538 & ~n7812 ) | ( n7811 & ~n7812 ) ;
  assign n7814 = n7707 ^ n7541 ^ x108 ;
  assign n7815 = n7723 ^ n7541 ^ 1'b0 ;
  assign n7816 = ( n7541 & n7814 ) | ( n7541 & ~n7815 ) | ( n7814 & ~n7815 ) ;
  assign n7817 = n7706 ^ n7544 ^ x107 ;
  assign n7818 = n7723 ^ n7544 ^ 1'b0 ;
  assign n7819 = ( n7544 & n7817 ) | ( n7544 & ~n7818 ) | ( n7817 & ~n7818 ) ;
  assign n7820 = n7705 ^ n7555 ^ x106 ;
  assign n7821 = n7723 ^ n7555 ^ 1'b0 ;
  assign n7822 = ( n7555 & n7820 ) | ( n7555 & ~n7821 ) | ( n7820 & ~n7821 ) ;
  assign n7823 = n7704 ^ n7558 ^ x105 ;
  assign n7824 = n7723 ^ n7558 ^ 1'b0 ;
  assign n7825 = ( n7558 & n7823 ) | ( n7558 & ~n7824 ) | ( n7823 & ~n7824 ) ;
  assign n7826 = n7703 ^ n7561 ^ x104 ;
  assign n7827 = n7723 ^ n7561 ^ 1'b0 ;
  assign n7828 = ( n7561 & n7826 ) | ( n7561 & ~n7827 ) | ( n7826 & ~n7827 ) ;
  assign n7829 = n7702 ^ n7564 ^ x103 ;
  assign n7830 = n7723 ^ n7564 ^ 1'b0 ;
  assign n7831 = ( n7564 & n7829 ) | ( n7564 & ~n7830 ) | ( n7829 & ~n7830 ) ;
  assign n7832 = n7701 ^ n7567 ^ x102 ;
  assign n7833 = n7723 ^ n7567 ^ 1'b0 ;
  assign n7834 = ( n7567 & n7832 ) | ( n7567 & ~n7833 ) | ( n7832 & ~n7833 ) ;
  assign n7835 = n7700 ^ n7570 ^ x101 ;
  assign n7836 = n7723 ^ n7570 ^ 1'b0 ;
  assign n7837 = ( n7570 & n7835 ) | ( n7570 & ~n7836 ) | ( n7835 & ~n7836 ) ;
  assign n7838 = n7699 ^ n7547 ^ x100 ;
  assign n7839 = n7723 ^ n7547 ^ 1'b0 ;
  assign n7840 = ( n7547 & n7838 ) | ( n7547 & ~n7839 ) | ( n7838 & ~n7839 ) ;
  assign n7841 = n7698 ^ n7550 ^ x99 ;
  assign n7842 = n7723 ^ n7550 ^ 1'b0 ;
  assign n7843 = ( n7550 & n7841 ) | ( n7550 & ~n7842 ) | ( n7841 & ~n7842 ) ;
  assign n7844 = n7697 ^ n7573 ^ x98 ;
  assign n7845 = n7723 ^ n7573 ^ 1'b0 ;
  assign n7846 = ( n7573 & n7844 ) | ( n7573 & ~n7845 ) | ( n7844 & ~n7845 ) ;
  assign n7847 = n7696 ^ n7482 ^ x97 ;
  assign n7848 = n7723 ^ n7482 ^ 1'b0 ;
  assign n7849 = ( n7482 & n7847 ) | ( n7482 & ~n7848 ) | ( n7847 & ~n7848 ) ;
  assign n7850 = n7695 ^ n7484 ^ x96 ;
  assign n7851 = n7723 ^ n7484 ^ 1'b0 ;
  assign n7852 = ( n7484 & n7850 ) | ( n7484 & ~n7851 ) | ( n7850 & ~n7851 ) ;
  assign n7853 = n7694 ^ n7486 ^ x95 ;
  assign n7854 = n7723 ^ n7486 ^ 1'b0 ;
  assign n7855 = ( n7486 & n7853 ) | ( n7486 & ~n7854 ) | ( n7853 & ~n7854 ) ;
  assign n7856 = n7693 ^ n7576 ^ x94 ;
  assign n7857 = n7723 ^ n7576 ^ 1'b0 ;
  assign n7858 = ( n7576 & n7856 ) | ( n7576 & ~n7857 ) | ( n7856 & ~n7857 ) ;
  assign n7859 = n7688 ^ n7579 ^ x93 ;
  assign n7860 = n7723 ^ n7579 ^ 1'b0 ;
  assign n7861 = ( n7579 & n7859 ) | ( n7579 & ~n7860 ) | ( n7859 & ~n7860 ) ;
  assign n7862 = x64 & n7723 ;
  assign n7863 = ~x7 & x64 ;
  assign n7864 = n7862 ^ x64 ^ x8 ;
  assign n7865 = n7864 ^ n7863 ^ x65 ;
  assign n7866 = ( x65 & n7863 ) | ( x65 & n7865 ) | ( n7863 & n7865 ) ;
  assign n7867 = n7866 ^ n7783 ^ x66 ;
  assign n7868 = ( x66 & n7866 ) | ( x66 & n7867 ) | ( n7866 & n7867 ) ;
  assign n7869 = ( x67 & ~n7781 ) | ( x67 & n7868 ) | ( ~n7781 & n7868 ) ;
  assign n7870 = ( x68 & ~n7779 ) | ( x68 & n7869 ) | ( ~n7779 & n7869 ) ;
  assign n7871 = ( x69 & ~n7732 ) | ( x69 & n7870 ) | ( ~n7732 & n7870 ) ;
  assign n7872 = ( x70 & ~n7777 ) | ( x70 & n7871 ) | ( ~n7777 & n7871 ) ;
  assign n7873 = ( x71 & ~n7775 ) | ( x71 & n7872 ) | ( ~n7775 & n7872 ) ;
  assign n7874 = ( x72 & ~n7773 ) | ( x72 & n7873 ) | ( ~n7773 & n7873 ) ;
  assign n7875 = ( x73 & ~n7771 ) | ( x73 & n7874 ) | ( ~n7771 & n7874 ) ;
  assign n7876 = ( x74 & ~n7769 ) | ( x74 & n7875 ) | ( ~n7769 & n7875 ) ;
  assign n7877 = ( x75 & ~n7729 ) | ( x75 & n7876 ) | ( ~n7729 & n7876 ) ;
  assign n7878 = ( x76 & ~n7767 ) | ( x76 & n7877 ) | ( ~n7767 & n7877 ) ;
  assign n7879 = ( x77 & ~n7737 ) | ( x77 & n7878 ) | ( ~n7737 & n7878 ) ;
  assign n7880 = ( x78 & ~n7765 ) | ( x78 & n7879 ) | ( ~n7765 & n7879 ) ;
  assign n7881 = ( x79 & ~n7763 ) | ( x79 & n7880 ) | ( ~n7763 & n7880 ) ;
  assign n7882 = ( x80 & ~n7761 ) | ( x80 & n7881 ) | ( ~n7761 & n7881 ) ;
  assign n7883 = ( x81 & ~n7759 ) | ( x81 & n7882 ) | ( ~n7759 & n7882 ) ;
  assign n7884 = ( x82 & ~n7757 ) | ( x82 & n7883 ) | ( ~n7757 & n7883 ) ;
  assign n7885 = ( x83 & ~n7755 ) | ( x83 & n7884 ) | ( ~n7755 & n7884 ) ;
  assign n7886 = ( x84 & ~n7727 ) | ( x84 & n7885 ) | ( ~n7727 & n7885 ) ;
  assign n7887 = ( x85 & ~n7753 ) | ( x85 & n7886 ) | ( ~n7753 & n7886 ) ;
  assign n7888 = ( x86 & ~n7751 ) | ( x86 & n7887 ) | ( ~n7751 & n7887 ) ;
  assign n7889 = ( x87 & ~n7749 ) | ( x87 & n7888 ) | ( ~n7749 & n7888 ) ;
  assign n7890 = ( x88 & ~n7747 ) | ( x88 & n7889 ) | ( ~n7747 & n7889 ) ;
  assign n7891 = n7872 ^ n7775 ^ x71 ;
  assign n7892 = ( x89 & ~n7745 ) | ( x89 & n7890 ) | ( ~n7745 & n7890 ) ;
  assign n7893 = n7871 ^ n7777 ^ x70 ;
  assign n7894 = n7875 ^ n7769 ^ x74 ;
  assign n7895 = n7876 ^ n7729 ^ x75 ;
  assign n7896 = ( x90 & ~n7743 ) | ( x90 & n7892 ) | ( ~n7743 & n7892 ) ;
  assign n7897 = n7878 ^ n7737 ^ x77 ;
  assign n7898 = n7879 ^ n7765 ^ x78 ;
  assign n7899 = ( x91 & ~n7741 ) | ( x91 & n7896 ) | ( ~n7741 & n7896 ) ;
  assign n7900 = n7881 ^ n7761 ^ x80 ;
  assign n7901 = n7882 ^ n7759 ^ x81 ;
  assign n7902 = n7883 ^ n7757 ^ x82 ;
  assign n7903 = n7884 ^ n7755 ^ x83 ;
  assign n7904 = n7885 ^ n7727 ^ x84 ;
  assign n7905 = n7886 ^ n7753 ^ x85 ;
  assign n7906 = n7887 ^ n7751 ^ x86 ;
  assign n7907 = n7888 ^ n7749 ^ x87 ;
  assign n7908 = ( x92 & ~n7739 ) | ( x92 & n7899 ) | ( ~n7739 & n7899 ) ;
  assign n7909 = ( x93 & ~n7740 ) | ( x93 & n7908 ) | ( ~n7740 & n7908 ) ;
  assign n7910 = ( x94 & ~n7861 ) | ( x94 & n7909 ) | ( ~n7861 & n7909 ) ;
  assign n7911 = ( x95 & ~n7858 ) | ( x95 & n7910 ) | ( ~n7858 & n7910 ) ;
  assign n7912 = ( x96 & ~n7855 ) | ( x96 & n7911 ) | ( ~n7855 & n7911 ) ;
  assign n7913 = ( x97 & ~n7852 ) | ( x97 & n7912 ) | ( ~n7852 & n7912 ) ;
  assign n7914 = ( x98 & ~n7849 ) | ( x98 & n7913 ) | ( ~n7849 & n7913 ) ;
  assign n7915 = n163 & n7738 ;
  assign n7916 = n7892 ^ n7743 ^ x90 ;
  assign n7917 = n7874 ^ n7771 ^ x73 ;
  assign n7918 = n7869 ^ n7779 ^ x68 ;
  assign n7919 = n7868 ^ n7781 ^ x67 ;
  assign n7920 = ( x99 & ~n7846 ) | ( x99 & n7914 ) | ( ~n7846 & n7914 ) ;
  assign n7921 = ( x100 & ~n7843 ) | ( x100 & n7920 ) | ( ~n7843 & n7920 ) ;
  assign n7922 = ( x101 & ~n7840 ) | ( x101 & n7921 ) | ( ~n7840 & n7921 ) ;
  assign n7923 = ( x102 & ~n7837 ) | ( x102 & n7922 ) | ( ~n7837 & n7922 ) ;
  assign n7924 = ( x103 & ~n7834 ) | ( x103 & n7923 ) | ( ~n7834 & n7923 ) ;
  assign n7925 = ( x104 & ~n7831 ) | ( x104 & n7924 ) | ( ~n7831 & n7924 ) ;
  assign n7926 = ( x105 & ~n7828 ) | ( x105 & n7925 ) | ( ~n7828 & n7925 ) ;
  assign n7927 = ( x106 & ~n7825 ) | ( x106 & n7926 ) | ( ~n7825 & n7926 ) ;
  assign n7928 = ( x107 & ~n7822 ) | ( x107 & n7927 ) | ( ~n7822 & n7927 ) ;
  assign n7929 = ( x108 & ~n7819 ) | ( x108 & n7928 ) | ( ~n7819 & n7928 ) ;
  assign n7930 = ( x109 & ~n7816 ) | ( x109 & n7929 ) | ( ~n7816 & n7929 ) ;
  assign n7931 = ( x110 & ~n7813 ) | ( x110 & n7930 ) | ( ~n7813 & n7930 ) ;
  assign n7932 = ( x111 & ~n7810 ) | ( x111 & n7931 ) | ( ~n7810 & n7931 ) ;
  assign n7933 = ( x112 & ~n7807 ) | ( x112 & n7932 ) | ( ~n7807 & n7932 ) ;
  assign n7934 = ( x113 & ~n7804 ) | ( x113 & n7933 ) | ( ~n7804 & n7933 ) ;
  assign n7935 = ( x114 & ~n7801 ) | ( x114 & n7934 ) | ( ~n7801 & n7934 ) ;
  assign n7936 = ( x115 & ~n7798 ) | ( x115 & n7935 ) | ( ~n7798 & n7935 ) ;
  assign n7937 = ( x116 & ~n7795 ) | ( x116 & n7936 ) | ( ~n7795 & n7936 ) ;
  assign n7938 = ( x117 & ~n7792 ) | ( x117 & n7937 ) | ( ~n7792 & n7937 ) ;
  assign n7939 = ( x118 & ~n7789 ) | ( x118 & n7938 ) | ( ~n7789 & n7938 ) ;
  assign n7940 = ( x119 & ~n7786 ) | ( x119 & n7939 ) | ( ~n7786 & n7939 ) ;
  assign n7941 = ( x120 & n156 ) | ( x120 & ~n7738 ) | ( n156 & ~n7738 ) ;
  assign n7942 = ( ~x120 & n7738 ) | ( ~x120 & n7940 ) | ( n7738 & n7940 ) ;
  assign n7943 = n7941 | n7942 ;
  assign n7944 = ( ~n7738 & n7915 ) | ( ~n7738 & n7943 ) | ( n7915 & n7943 ) ;
  assign n7945 = n7940 ^ n7738 ^ x120 ;
  assign n7946 = n7944 ^ n7777 ^ 1'b0 ;
  assign n7947 = ( n7777 & n7893 ) | ( n7777 & ~n7946 ) | ( n7893 & ~n7946 ) ;
  assign n7948 = n7944 ^ n7769 ^ 1'b0 ;
  assign n7949 = n7944 ^ n7867 ^ 1'b0 ;
  assign n7950 = n7915 & ~n7943 ;
  assign n7951 = ( n7769 & n7894 ) | ( n7769 & ~n7948 ) | ( n7894 & ~n7948 ) ;
  assign n7952 = n7944 ^ n7765 ^ 1'b0 ;
  assign n7953 = n7944 ^ n7779 ^ 1'b0 ;
  assign n7954 = ( n7783 & n7867 ) | ( n7783 & n7949 ) | ( n7867 & n7949 ) ;
  assign n7955 = ( n7765 & n7898 ) | ( n7765 & ~n7952 ) | ( n7898 & ~n7952 ) ;
  assign n7956 = n7944 ^ n7865 ^ 1'b0 ;
  assign n7957 = n7944 ^ n7775 ^ 1'b0 ;
  assign n7958 = n7944 ^ n7737 ^ 1'b0 ;
  assign n7959 = ( n7864 & n7865 ) | ( n7864 & n7956 ) | ( n7865 & n7956 ) ;
  assign n7960 = n7944 ^ n7743 ^ 1'b0 ;
  assign n7961 = n7944 ^ n7761 ^ 1'b0 ;
  assign n7962 = n7944 ^ n7755 ^ 1'b0 ;
  assign n7963 = ( n7755 & n7903 ) | ( n7755 & ~n7962 ) | ( n7903 & ~n7962 ) ;
  assign n7964 = ( n7743 & n7916 ) | ( n7743 & ~n7960 ) | ( n7916 & ~n7960 ) ;
  assign n7965 = ~n7944 & n7945 ;
  assign n7966 = ( n7779 & n7918 ) | ( n7779 & ~n7953 ) | ( n7918 & ~n7953 ) ;
  assign n7967 = ( n7915 & ~n7950 ) | ( n7915 & n7965 ) | ( ~n7950 & n7965 ) ;
  assign n7968 = ( n7761 & n7900 ) | ( n7761 & ~n7961 ) | ( n7900 & ~n7961 ) ;
  assign n7969 = ( n7737 & n7897 ) | ( n7737 & ~n7958 ) | ( n7897 & ~n7958 ) ;
  assign n7970 = ( n7775 & n7891 ) | ( n7775 & ~n7957 ) | ( n7891 & ~n7957 ) ;
  assign n7971 = n7944 ^ n7727 ^ 1'b0 ;
  assign n7972 = n7944 ^ n7757 ^ 1'b0 ;
  assign n7973 = n7944 ^ n7751 ^ 1'b0 ;
  assign n7974 = n7944 ^ n7781 ^ 1'b0 ;
  assign n7975 = n7944 ^ n7759 ^ 1'b0 ;
  assign n7976 = ( n7757 & n7902 ) | ( n7757 & ~n7972 ) | ( n7902 & ~n7972 ) ;
  assign n7977 = ( n7759 & n7901 ) | ( n7759 & ~n7975 ) | ( n7901 & ~n7975 ) ;
  assign n7978 = n7944 ^ n7771 ^ 1'b0 ;
  assign n7979 = n7944 ^ n7753 ^ 1'b0 ;
  assign n7980 = ( n7753 & n7905 ) | ( n7753 & ~n7979 ) | ( n7905 & ~n7979 ) ;
  assign n7981 = n7944 ^ n7749 ^ 1'b0 ;
  assign n7982 = ( n7749 & n7907 ) | ( n7749 & ~n7981 ) | ( n7907 & ~n7981 ) ;
  assign n7983 = n7944 ^ n7729 ^ 1'b0 ;
  assign n7984 = ( n7729 & n7895 ) | ( n7729 & ~n7983 ) | ( n7895 & ~n7983 ) ;
  assign n7985 = ( n7751 & n7906 ) | ( n7751 & ~n7973 ) | ( n7906 & ~n7973 ) ;
  assign n7986 = ( n7781 & n7919 ) | ( n7781 & ~n7974 ) | ( n7919 & ~n7974 ) ;
  assign n7987 = ( n7771 & n7917 ) | ( n7771 & ~n7978 ) | ( n7917 & ~n7978 ) ;
  assign n7988 = ( n7727 & n7904 ) | ( n7727 & ~n7971 ) | ( n7904 & ~n7971 ) ;
  assign n7989 = n7939 ^ n7786 ^ x119 ;
  assign n7990 = n7944 ^ n7786 ^ 1'b0 ;
  assign n7991 = ( n7786 & n7989 ) | ( n7786 & ~n7990 ) | ( n7989 & ~n7990 ) ;
  assign n7992 = n7938 ^ n7789 ^ x118 ;
  assign n7993 = n7944 ^ n7789 ^ 1'b0 ;
  assign n7994 = ( n7789 & n7992 ) | ( n7789 & ~n7993 ) | ( n7992 & ~n7993 ) ;
  assign n7995 = n7937 ^ n7792 ^ x117 ;
  assign n7996 = n7944 ^ n7792 ^ 1'b0 ;
  assign n7997 = ( n7792 & n7995 ) | ( n7792 & ~n7996 ) | ( n7995 & ~n7996 ) ;
  assign n7998 = n7920 ^ n7843 ^ x100 ;
  assign n7999 = n7944 ^ n7843 ^ 1'b0 ;
  assign n8000 = ( n7843 & n7998 ) | ( n7843 & ~n7999 ) | ( n7998 & ~n7999 ) ;
  assign n8001 = n7914 ^ n7846 ^ x99 ;
  assign n8002 = n7944 ^ n7846 ^ 1'b0 ;
  assign n8003 = ( n7846 & n8001 ) | ( n7846 & ~n8002 ) | ( n8001 & ~n8002 ) ;
  assign n8004 = n7913 ^ n7849 ^ x98 ;
  assign n8005 = n7944 ^ n7849 ^ 1'b0 ;
  assign n8006 = n7912 ^ n7852 ^ x97 ;
  assign n8007 = n7944 ^ n7852 ^ 1'b0 ;
  assign n8008 = ( n7852 & n8006 ) | ( n7852 & ~n8007 ) | ( n8006 & ~n8007 ) ;
  assign n8009 = n7911 ^ n7855 ^ x96 ;
  assign n8010 = n7944 ^ n7855 ^ 1'b0 ;
  assign n8011 = ( n7855 & n8009 ) | ( n7855 & ~n8010 ) | ( n8009 & ~n8010 ) ;
  assign n8012 = n7910 ^ n7858 ^ x95 ;
  assign n8013 = n7944 ^ n7858 ^ 1'b0 ;
  assign n8014 = ( n7858 & n8012 ) | ( n7858 & ~n8013 ) | ( n8012 & ~n8013 ) ;
  assign n8015 = n7909 ^ n7861 ^ x94 ;
  assign n8016 = n7944 ^ n7861 ^ 1'b0 ;
  assign n8017 = ( n7861 & n8015 ) | ( n7861 & ~n8016 ) | ( n8015 & ~n8016 ) ;
  assign n8018 = n7908 ^ n7740 ^ x93 ;
  assign n8019 = n7944 ^ n7740 ^ 1'b0 ;
  assign n8020 = ( n7740 & n8018 ) | ( n7740 & ~n8019 ) | ( n8018 & ~n8019 ) ;
  assign n8021 = n7899 ^ n7739 ^ x92 ;
  assign n8022 = n7944 ^ n7739 ^ 1'b0 ;
  assign n8023 = ( n7739 & n8021 ) | ( n7739 & ~n8022 ) | ( n8021 & ~n8022 ) ;
  assign n8024 = n7896 ^ n7741 ^ x91 ;
  assign n8025 = n7944 ^ n7741 ^ 1'b0 ;
  assign n8026 = ( n7741 & n8024 ) | ( n7741 & ~n8025 ) | ( n8024 & ~n8025 ) ;
  assign n8027 = n7890 ^ n7745 ^ x89 ;
  assign n8028 = n7944 ^ n7745 ^ 1'b0 ;
  assign n8029 = ( n7745 & n8027 ) | ( n7745 & ~n8028 ) | ( n8027 & ~n8028 ) ;
  assign n8030 = n7889 ^ n7747 ^ x88 ;
  assign n8031 = n7944 ^ n7747 ^ 1'b0 ;
  assign n8032 = ( n7747 & n8030 ) | ( n7747 & ~n8031 ) | ( n8030 & ~n8031 ) ;
  assign n8033 = n7880 ^ n7763 ^ x79 ;
  assign n8034 = n7944 ^ n7763 ^ 1'b0 ;
  assign n8035 = ( n7763 & n8033 ) | ( n7763 & ~n8034 ) | ( n8033 & ~n8034 ) ;
  assign n8036 = n7877 ^ n7767 ^ x76 ;
  assign n8037 = n7944 ^ n7767 ^ 1'b0 ;
  assign n8038 = ( n7767 & n8036 ) | ( n7767 & ~n8037 ) | ( n8036 & ~n8037 ) ;
  assign n8039 = n7873 ^ n7773 ^ x72 ;
  assign n8040 = n7944 ^ n7773 ^ 1'b0 ;
  assign n8041 = ( n7773 & n8039 ) | ( n7773 & ~n8040 ) | ( n8039 & ~n8040 ) ;
  assign n8042 = n7870 ^ n7732 ^ x69 ;
  assign n8043 = n7944 ^ n7732 ^ 1'b0 ;
  assign n8044 = ( n7732 & n8042 ) | ( n7732 & ~n8043 ) | ( n8042 & ~n8043 ) ;
  assign n8045 = ( n7849 & n8004 ) | ( n7849 & ~n8005 ) | ( n8004 & ~n8005 ) ;
  assign n8046 = n7936 ^ n7795 ^ x116 ;
  assign n8047 = n7944 ^ n7795 ^ 1'b0 ;
  assign n8048 = ( n7795 & n8046 ) | ( n7795 & ~n8047 ) | ( n8046 & ~n8047 ) ;
  assign n8049 = n7935 ^ n7798 ^ x115 ;
  assign n8050 = n7944 ^ n7798 ^ 1'b0 ;
  assign n8051 = ( n7798 & n8049 ) | ( n7798 & ~n8050 ) | ( n8049 & ~n8050 ) ;
  assign n8052 = n7934 ^ n7801 ^ x114 ;
  assign n8053 = n7944 ^ n7801 ^ 1'b0 ;
  assign n8054 = ( n7801 & n8052 ) | ( n7801 & ~n8053 ) | ( n8052 & ~n8053 ) ;
  assign n8055 = n7933 ^ n7804 ^ x113 ;
  assign n8056 = n7944 ^ n7804 ^ 1'b0 ;
  assign n8057 = ( n7804 & n8055 ) | ( n7804 & ~n8056 ) | ( n8055 & ~n8056 ) ;
  assign n8058 = n7932 ^ n7807 ^ x112 ;
  assign n8059 = n7944 ^ n7807 ^ 1'b0 ;
  assign n8060 = ( n7807 & n8058 ) | ( n7807 & ~n8059 ) | ( n8058 & ~n8059 ) ;
  assign n8061 = n7931 ^ n7810 ^ x111 ;
  assign n8062 = n7944 ^ n7810 ^ 1'b0 ;
  assign n8063 = ( n7810 & n8061 ) | ( n7810 & ~n8062 ) | ( n8061 & ~n8062 ) ;
  assign n8064 = n7944 ^ n7813 ^ 1'b0 ;
  assign n8065 = n7929 ^ n7816 ^ x109 ;
  assign n8066 = n7944 ^ n7816 ^ 1'b0 ;
  assign n8067 = ( n7816 & n8065 ) | ( n7816 & ~n8066 ) | ( n8065 & ~n8066 ) ;
  assign n8068 = n7928 ^ n7819 ^ x108 ;
  assign n8069 = n7944 ^ n7819 ^ 1'b0 ;
  assign n8070 = n7930 ^ n7813 ^ x110 ;
  assign n8071 = ( n7813 & ~n8064 ) | ( n7813 & n8070 ) | ( ~n8064 & n8070 ) ;
  assign n8072 = ( n7819 & n8068 ) | ( n7819 & ~n8069 ) | ( n8068 & ~n8069 ) ;
  assign n8073 = n7927 ^ n7822 ^ x107 ;
  assign n8074 = n7944 ^ n7822 ^ 1'b0 ;
  assign n8075 = ( n7822 & n8073 ) | ( n7822 & ~n8074 ) | ( n8073 & ~n8074 ) ;
  assign n8076 = n7926 ^ n7825 ^ x106 ;
  assign n8077 = n7944 ^ n7825 ^ 1'b0 ;
  assign n8078 = ( n7825 & n8076 ) | ( n7825 & ~n8077 ) | ( n8076 & ~n8077 ) ;
  assign n8079 = n7925 ^ n7828 ^ x105 ;
  assign n8080 = n7944 ^ n7828 ^ 1'b0 ;
  assign n8081 = ( n7828 & n8079 ) | ( n7828 & ~n8080 ) | ( n8079 & ~n8080 ) ;
  assign n8082 = n7924 ^ n7831 ^ x104 ;
  assign n8083 = n7944 ^ n7831 ^ 1'b0 ;
  assign n8084 = ( n7831 & n8082 ) | ( n7831 & ~n8083 ) | ( n8082 & ~n8083 ) ;
  assign n8085 = n7923 ^ n7834 ^ x103 ;
  assign n8086 = n7944 ^ n7834 ^ 1'b0 ;
  assign n8087 = ( n7834 & n8085 ) | ( n7834 & ~n8086 ) | ( n8085 & ~n8086 ) ;
  assign n8088 = n7922 ^ n7837 ^ x102 ;
  assign n8089 = n7944 ^ n7837 ^ 1'b0 ;
  assign n8090 = ( n7837 & n8088 ) | ( n7837 & ~n8089 ) | ( n8088 & ~n8089 ) ;
  assign n8091 = n7921 ^ n7840 ^ x101 ;
  assign n8092 = n7944 ^ n7840 ^ 1'b0 ;
  assign n8093 = ( n7840 & n8091 ) | ( n7840 & ~n8092 ) | ( n8091 & ~n8092 ) ;
  assign n8094 = x64 & n7944 ;
  assign n8095 = n8094 ^ x64 ^ x7 ;
  assign n8096 = ~x6 & x64 ;
  assign n8097 = n8096 ^ n8095 ^ x65 ;
  assign n8098 = ( x65 & n8096 ) | ( x65 & n8097 ) | ( n8096 & n8097 ) ;
  assign n8099 = n8098 ^ n7959 ^ x66 ;
  assign n8100 = ( x66 & n8098 ) | ( x66 & n8099 ) | ( n8098 & n8099 ) ;
  assign n8101 = ( x67 & ~n7954 ) | ( x67 & n8100 ) | ( ~n7954 & n8100 ) ;
  assign n8102 = ( x68 & ~n7986 ) | ( x68 & n8101 ) | ( ~n7986 & n8101 ) ;
  assign n8103 = ( x69 & ~n7966 ) | ( x69 & n8102 ) | ( ~n7966 & n8102 ) ;
  assign n8104 = ( x70 & ~n8044 ) | ( x70 & n8103 ) | ( ~n8044 & n8103 ) ;
  assign n8105 = ( x71 & ~n7947 ) | ( x71 & n8104 ) | ( ~n7947 & n8104 ) ;
  assign n8106 = ( x72 & ~n7970 ) | ( x72 & n8105 ) | ( ~n7970 & n8105 ) ;
  assign n8107 = ( x73 & ~n8041 ) | ( x73 & n8106 ) | ( ~n8041 & n8106 ) ;
  assign n8108 = ( x74 & ~n7987 ) | ( x74 & n8107 ) | ( ~n7987 & n8107 ) ;
  assign n8109 = ( x75 & ~n7951 ) | ( x75 & n8108 ) | ( ~n7951 & n8108 ) ;
  assign n8110 = ( x76 & ~n7984 ) | ( x76 & n8109 ) | ( ~n7984 & n8109 ) ;
  assign n8111 = ( x77 & ~n8038 ) | ( x77 & n8110 ) | ( ~n8038 & n8110 ) ;
  assign n8112 = ( x78 & ~n7969 ) | ( x78 & n8111 ) | ( ~n7969 & n8111 ) ;
  assign n8113 = ( x79 & ~n7955 ) | ( x79 & n8112 ) | ( ~n7955 & n8112 ) ;
  assign n8114 = ( x80 & ~n8035 ) | ( x80 & n8113 ) | ( ~n8035 & n8113 ) ;
  assign n8115 = ( x81 & ~n7968 ) | ( x81 & n8114 ) | ( ~n7968 & n8114 ) ;
  assign n8116 = ( x82 & ~n7977 ) | ( x82 & n8115 ) | ( ~n7977 & n8115 ) ;
  assign n8117 = ( x83 & ~n7976 ) | ( x83 & n8116 ) | ( ~n7976 & n8116 ) ;
  assign n8118 = ( x84 & ~n7963 ) | ( x84 & n8117 ) | ( ~n7963 & n8117 ) ;
  assign n8119 = ( x85 & ~n7988 ) | ( x85 & n8118 ) | ( ~n7988 & n8118 ) ;
  assign n8120 = ( x86 & ~n7980 ) | ( x86 & n8119 ) | ( ~n7980 & n8119 ) ;
  assign n8121 = ( x87 & ~n7985 ) | ( x87 & n8120 ) | ( ~n7985 & n8120 ) ;
  assign n8122 = ( x88 & ~n7982 ) | ( x88 & n8121 ) | ( ~n7982 & n8121 ) ;
  assign n8123 = ( x89 & ~n8032 ) | ( x89 & n8122 ) | ( ~n8032 & n8122 ) ;
  assign n8124 = ( x90 & ~n8029 ) | ( x90 & n8123 ) | ( ~n8029 & n8123 ) ;
  assign n8125 = ( x91 & ~n7964 ) | ( x91 & n8124 ) | ( ~n7964 & n8124 ) ;
  assign n8126 = ( x92 & ~n8026 ) | ( x92 & n8125 ) | ( ~n8026 & n8125 ) ;
  assign n8127 = ( x93 & ~n8023 ) | ( x93 & n8126 ) | ( ~n8023 & n8126 ) ;
  assign n8128 = ( x94 & ~n8020 ) | ( x94 & n8127 ) | ( ~n8020 & n8127 ) ;
  assign n8129 = ( x95 & ~n8017 ) | ( x95 & n8128 ) | ( ~n8017 & n8128 ) ;
  assign n8130 = ( x96 & ~n8014 ) | ( x96 & n8129 ) | ( ~n8014 & n8129 ) ;
  assign n8131 = ( x97 & ~n8011 ) | ( x97 & n8130 ) | ( ~n8011 & n8130 ) ;
  assign n8132 = ( x98 & ~n8008 ) | ( x98 & n8131 ) | ( ~n8008 & n8131 ) ;
  assign n8133 = ( x99 & ~n8045 ) | ( x99 & n8132 ) | ( ~n8045 & n8132 ) ;
  assign n8134 = ( x100 & ~n8003 ) | ( x100 & n8133 ) | ( ~n8003 & n8133 ) ;
  assign n8135 = n8119 ^ n7980 ^ x86 ;
  assign n8136 = n8120 ^ n7985 ^ x87 ;
  assign n8137 = n8121 ^ n7982 ^ x88 ;
  assign n8138 = n8117 ^ n7963 ^ x84 ;
  assign n8139 = n8116 ^ n7976 ^ x83 ;
  assign n8140 = n8113 ^ n8035 ^ x80 ;
  assign n8141 = n8125 ^ n8026 ^ x92 ;
  assign n8142 = n8126 ^ n8023 ^ x93 ;
  assign n8143 = n8134 ^ n8000 ^ x101 ;
  assign n8144 = ( x101 & ~n8000 ) | ( x101 & n8134 ) | ( ~n8000 & n8134 ) ;
  assign n8145 = n8131 ^ n8008 ^ x98 ;
  assign n8146 = n8111 ^ n7969 ^ x78 ;
  assign n8147 = n8110 ^ n8038 ^ x77 ;
  assign n8148 = n8108 ^ n7951 ^ x75 ;
  assign n8149 = n8106 ^ n8041 ^ x73 ;
  assign n8150 = n8101 ^ n7986 ^ x68 ;
  assign n8151 = n8100 ^ n7954 ^ x67 ;
  assign n8152 = ( x102 & ~n8093 ) | ( x102 & n8144 ) | ( ~n8093 & n8144 ) ;
  assign n8153 = ( x103 & ~n8090 ) | ( x103 & n8152 ) | ( ~n8090 & n8152 ) ;
  assign n8154 = ( x104 & ~n8087 ) | ( x104 & n8153 ) | ( ~n8087 & n8153 ) ;
  assign n8155 = ( x105 & ~n8084 ) | ( x105 & n8154 ) | ( ~n8084 & n8154 ) ;
  assign n8156 = ( x106 & ~n8081 ) | ( x106 & n8155 ) | ( ~n8081 & n8155 ) ;
  assign n8157 = ( x107 & ~n8078 ) | ( x107 & n8156 ) | ( ~n8078 & n8156 ) ;
  assign n8158 = ( x108 & ~n8075 ) | ( x108 & n8157 ) | ( ~n8075 & n8157 ) ;
  assign n8159 = ( x109 & ~n8072 ) | ( x109 & n8158 ) | ( ~n8072 & n8158 ) ;
  assign n8160 = ( x110 & ~n8067 ) | ( x110 & n8159 ) | ( ~n8067 & n8159 ) ;
  assign n8161 = ( x111 & ~n8071 ) | ( x111 & n8160 ) | ( ~n8071 & n8160 ) ;
  assign n8162 = ( x112 & ~n8063 ) | ( x112 & n8161 ) | ( ~n8063 & n8161 ) ;
  assign n8163 = ( x113 & ~n8060 ) | ( x113 & n8162 ) | ( ~n8060 & n8162 ) ;
  assign n8164 = ( x114 & ~n8057 ) | ( x114 & n8163 ) | ( ~n8057 & n8163 ) ;
  assign n8165 = ( x115 & ~n8054 ) | ( x115 & n8164 ) | ( ~n8054 & n8164 ) ;
  assign n8166 = ( x116 & ~n8051 ) | ( x116 & n8165 ) | ( ~n8051 & n8165 ) ;
  assign n8167 = ( x117 & ~n8048 ) | ( x117 & n8166 ) | ( ~n8048 & n8166 ) ;
  assign n8168 = ( x118 & ~n7997 ) | ( x118 & n8167 ) | ( ~n7997 & n8167 ) ;
  assign n8169 = ( x119 & ~n7994 ) | ( x119 & n8168 ) | ( ~n7994 & n8168 ) ;
  assign n8170 = ( x120 & ~n7991 ) | ( x120 & n8169 ) | ( ~n7991 & n8169 ) ;
  assign n8171 = ( x121 & ~n7967 ) | ( x121 & n8170 ) | ( ~n7967 & n8170 ) ;
  assign n8172 = n155 | n8171 ;
  assign n8173 = n8156 ^ n8078 ^ x107 ;
  assign n8174 = n8172 ^ n8145 ^ 1'b0 ;
  assign n8175 = ( n8008 & n8145 ) | ( n8008 & n8174 ) | ( n8145 & n8174 ) ;
  assign n8176 = n8172 ^ n7959 ^ 1'b0 ;
  assign n8177 = n8172 ^ n8146 ^ 1'b0 ;
  assign n8178 = ( n7959 & n8099 ) | ( n7959 & ~n8176 ) | ( n8099 & ~n8176 ) ;
  assign n8179 = n8172 ^ n8149 ^ 1'b0 ;
  assign n8180 = n8172 ^ n8148 ^ 1'b0 ;
  assign n8181 = ( n7969 & n8146 ) | ( n7969 & n8177 ) | ( n8146 & n8177 ) ;
  assign n8182 = ( n8041 & n8149 ) | ( n8041 & n8179 ) | ( n8149 & n8179 ) ;
  assign n8183 = n8172 ^ n8150 ^ 1'b0 ;
  assign n8184 = n8172 ^ n8142 ^ 1'b0 ;
  assign n8185 = n8172 ^ n8137 ^ 1'b0 ;
  assign n8186 = ( n7982 & n8137 ) | ( n7982 & n8185 ) | ( n8137 & n8185 ) ;
  assign n8187 = n8173 ^ n8172 ^ 1'b0 ;
  assign n8188 = n8155 ^ n8081 ^ x106 ;
  assign n8189 = n8172 ^ n8140 ^ 1'b0 ;
  assign n8190 = ( n8035 & n8140 ) | ( n8035 & n8189 ) | ( n8140 & n8189 ) ;
  assign n8191 = n8172 ^ n8151 ^ 1'b0 ;
  assign n8192 = ( n7954 & n8151 ) | ( n7954 & n8191 ) | ( n8151 & n8191 ) ;
  assign n8193 = n8154 ^ n8084 ^ x105 ;
  assign n8194 = n8172 ^ n8139 ^ 1'b0 ;
  assign n8195 = ( n8023 & n8142 ) | ( n8023 & n8184 ) | ( n8142 & n8184 ) ;
  assign n8196 = ( n7976 & n8139 ) | ( n7976 & n8194 ) | ( n8139 & n8194 ) ;
  assign n8197 = n8193 ^ n8172 ^ 1'b0 ;
  assign n8198 = ( n7986 & n8150 ) | ( n7986 & n8183 ) | ( n8150 & n8183 ) ;
  assign n8199 = n8172 ^ n8095 ^ 1'b0 ;
  assign n8200 = n8172 ^ n8147 ^ 1'b0 ;
  assign n8201 = ( n8095 & n8097 ) | ( n8095 & ~n8199 ) | ( n8097 & ~n8199 ) ;
  assign n8202 = ( n8084 & n8193 ) | ( n8084 & n8197 ) | ( n8193 & n8197 ) ;
  assign n8203 = ( n8038 & n8147 ) | ( n8038 & n8200 ) | ( n8147 & n8200 ) ;
  assign n8204 = n8157 ^ n8075 ^ x108 ;
  assign n8205 = ( n7951 & n8148 ) | ( n7951 & n8180 ) | ( n8148 & n8180 ) ;
  assign n8206 = n8188 ^ n8172 ^ 1'b0 ;
  assign n8207 = n8172 ^ n8143 ^ 1'b0 ;
  assign n8208 = n8172 ^ n8138 ^ 1'b0 ;
  assign n8209 = ( n7963 & n8138 ) | ( n7963 & n8208 ) | ( n8138 & n8208 ) ;
  assign n8210 = n8204 ^ n8172 ^ 1'b0 ;
  assign n8211 = n8172 ^ n8135 ^ 1'b0 ;
  assign n8212 = n8172 ^ n8141 ^ 1'b0 ;
  assign n8213 = ( n8075 & n8204 ) | ( n8075 & n8210 ) | ( n8204 & n8210 ) ;
  assign n8214 = ( n8081 & n8188 ) | ( n8081 & n8206 ) | ( n8188 & n8206 ) ;
  assign n8215 = n8172 ^ n8136 ^ 1'b0 ;
  assign n8216 = ( n8000 & n8143 ) | ( n8000 & n8207 ) | ( n8143 & n8207 ) ;
  assign n8217 = ( n7980 & n8135 ) | ( n7980 & n8211 ) | ( n8135 & n8211 ) ;
  assign n8218 = ( n8078 & n8173 ) | ( n8078 & n8187 ) | ( n8173 & n8187 ) ;
  assign n8219 = ( n7985 & n8136 ) | ( n7985 & n8215 ) | ( n8136 & n8215 ) ;
  assign n8220 = ( n8026 & n8141 ) | ( n8026 & n8212 ) | ( n8141 & n8212 ) ;
  assign n8221 = n8169 ^ n7991 ^ x120 ;
  assign n8222 = n8221 ^ n8172 ^ 1'b0 ;
  assign n8223 = ( n7991 & n8221 ) | ( n7991 & n8222 ) | ( n8221 & n8222 ) ;
  assign n8224 = n8167 ^ n7997 ^ x118 ;
  assign n8225 = n8224 ^ n8172 ^ 1'b0 ;
  assign n8226 = ( n7997 & n8224 ) | ( n7997 & n8225 ) | ( n8224 & n8225 ) ;
  assign n8227 = n8165 ^ n8051 ^ x116 ;
  assign n8228 = n8227 ^ n8172 ^ 1'b0 ;
  assign n8229 = ( n8051 & n8227 ) | ( n8051 & n8228 ) | ( n8227 & n8228 ) ;
  assign n8230 = n8164 ^ n8054 ^ x115 ;
  assign n8231 = n8230 ^ n8172 ^ 1'b0 ;
  assign n8232 = ( n8054 & n8230 ) | ( n8054 & n8231 ) | ( n8230 & n8231 ) ;
  assign n8233 = n8163 ^ n8057 ^ x114 ;
  assign n8234 = n8233 ^ n8172 ^ 1'b0 ;
  assign n8235 = ( n8057 & n8233 ) | ( n8057 & n8234 ) | ( n8233 & n8234 ) ;
  assign n8236 = n8162 ^ n8060 ^ x113 ;
  assign n8237 = n8236 ^ n8172 ^ 1'b0 ;
  assign n8238 = ( n8060 & n8236 ) | ( n8060 & n8237 ) | ( n8236 & n8237 ) ;
  assign n8239 = n8161 ^ n8063 ^ x112 ;
  assign n8240 = n8239 ^ n8172 ^ 1'b0 ;
  assign n8241 = ( n8063 & n8239 ) | ( n8063 & n8240 ) | ( n8239 & n8240 ) ;
  assign n8242 = n8160 ^ n8071 ^ x111 ;
  assign n8243 = n8242 ^ n8172 ^ 1'b0 ;
  assign n8244 = ( n8071 & n8242 ) | ( n8071 & n8243 ) | ( n8242 & n8243 ) ;
  assign n8245 = n8159 ^ n8067 ^ x110 ;
  assign n8246 = n8158 ^ n8072 ^ x109 ;
  assign n8247 = n8246 ^ n8172 ^ 1'b0 ;
  assign n8248 = ( n8072 & n8246 ) | ( n8072 & n8247 ) | ( n8246 & n8247 ) ;
  assign n8249 = n8153 ^ n8087 ^ x104 ;
  assign n8250 = n8249 ^ n8172 ^ 1'b0 ;
  assign n8251 = ( n8087 & n8249 ) | ( n8087 & n8250 ) | ( n8249 & n8250 ) ;
  assign n8252 = n8144 ^ n8093 ^ x102 ;
  assign n8253 = n8252 ^ n8172 ^ 1'b0 ;
  assign n8254 = ( n8093 & n8252 ) | ( n8093 & n8253 ) | ( n8252 & n8253 ) ;
  assign n8255 = n8132 ^ n8045 ^ x99 ;
  assign n8256 = n8255 ^ n8172 ^ 1'b0 ;
  assign n8257 = ( n8045 & n8255 ) | ( n8045 & n8256 ) | ( n8255 & n8256 ) ;
  assign n8258 = n8129 ^ n8014 ^ x96 ;
  assign n8259 = n8258 ^ n8172 ^ 1'b0 ;
  assign n8260 = ( n8014 & n8258 ) | ( n8014 & n8259 ) | ( n8258 & n8259 ) ;
  assign n8261 = n8245 ^ n8172 ^ 1'b0 ;
  assign n8262 = ( n8067 & n8245 ) | ( n8067 & n8261 ) | ( n8245 & n8261 ) ;
  assign n8263 = n8124 ^ n7964 ^ x91 ;
  assign n8264 = n8263 ^ n8172 ^ 1'b0 ;
  assign n8265 = ( n7964 & n8263 ) | ( n7964 & n8264 ) | ( n8263 & n8264 ) ;
  assign n8266 = n8122 ^ n8032 ^ x89 ;
  assign n8267 = n8266 ^ n8172 ^ 1'b0 ;
  assign n8268 = ( n8032 & n8266 ) | ( n8032 & n8267 ) | ( n8266 & n8267 ) ;
  assign n8269 = n8112 ^ n7955 ^ x79 ;
  assign n8270 = n8269 ^ n8172 ^ 1'b0 ;
  assign n8271 = ( n7955 & n8269 ) | ( n7955 & n8270 ) | ( n8269 & n8270 ) ;
  assign n8272 = n8109 ^ n7984 ^ x76 ;
  assign n8273 = n8272 ^ n8172 ^ 1'b0 ;
  assign n8274 = ( n7984 & n8272 ) | ( n7984 & n8273 ) | ( n8272 & n8273 ) ;
  assign n8275 = n8107 ^ n7987 ^ x74 ;
  assign n8276 = n8275 ^ n8172 ^ 1'b0 ;
  assign n8277 = ( n7987 & n8275 ) | ( n7987 & n8276 ) | ( n8275 & n8276 ) ;
  assign n8278 = n8168 ^ n7994 ^ x119 ;
  assign n8279 = n8278 ^ n8172 ^ 1'b0 ;
  assign n8280 = ( n7994 & n8278 ) | ( n7994 & n8279 ) | ( n8278 & n8279 ) ;
  assign n8281 = n8166 ^ n8048 ^ x117 ;
  assign n8282 = n8281 ^ n8172 ^ 1'b0 ;
  assign n8283 = ( n8048 & n8281 ) | ( n8048 & n8282 ) | ( n8281 & n8282 ) ;
  assign n8284 = n8152 ^ n8090 ^ x103 ;
  assign n8285 = n8284 ^ n8172 ^ 1'b0 ;
  assign n8286 = ( n8090 & n8284 ) | ( n8090 & n8285 ) | ( n8284 & n8285 ) ;
  assign n8287 = n8133 ^ n8003 ^ x100 ;
  assign n8288 = n8287 ^ n8172 ^ 1'b0 ;
  assign n8289 = ( n8003 & n8287 ) | ( n8003 & n8288 ) | ( n8287 & n8288 ) ;
  assign n8290 = n8130 ^ n8011 ^ x97 ;
  assign n8291 = n8290 ^ n8172 ^ 1'b0 ;
  assign n8292 = ( n8011 & n8290 ) | ( n8011 & n8291 ) | ( n8290 & n8291 ) ;
  assign n8293 = n8128 ^ n8017 ^ x95 ;
  assign n8294 = n8293 ^ n8172 ^ 1'b0 ;
  assign n8295 = ( n8017 & n8293 ) | ( n8017 & n8294 ) | ( n8293 & n8294 ) ;
  assign n8296 = n8127 ^ n8020 ^ x94 ;
  assign n8297 = n8296 ^ n8172 ^ 1'b0 ;
  assign n8298 = ( n8020 & n8296 ) | ( n8020 & n8297 ) | ( n8296 & n8297 ) ;
  assign n8299 = n8123 ^ n8029 ^ x90 ;
  assign n8300 = n8299 ^ n8172 ^ 1'b0 ;
  assign n8301 = ( n8029 & n8299 ) | ( n8029 & n8300 ) | ( n8299 & n8300 ) ;
  assign n8302 = n8118 ^ n7988 ^ x85 ;
  assign n8303 = n8302 ^ n8172 ^ 1'b0 ;
  assign n8304 = ( n7988 & n8302 ) | ( n7988 & n8303 ) | ( n8302 & n8303 ) ;
  assign n8305 = n8115 ^ n7977 ^ x82 ;
  assign n8306 = n8305 ^ n8172 ^ 1'b0 ;
  assign n8307 = ( n7977 & n8305 ) | ( n7977 & n8306 ) | ( n8305 & n8306 ) ;
  assign n8308 = n8114 ^ n7968 ^ x81 ;
  assign n8309 = n8308 ^ n8172 ^ 1'b0 ;
  assign n8310 = ( n7968 & n8308 ) | ( n7968 & n8309 ) | ( n8308 & n8309 ) ;
  assign n8311 = n8105 ^ n7970 ^ x72 ;
  assign n8312 = n8311 ^ n8172 ^ 1'b0 ;
  assign n8313 = ( n7970 & n8311 ) | ( n7970 & n8312 ) | ( n8311 & n8312 ) ;
  assign n8314 = n8104 ^ n7947 ^ x71 ;
  assign n8315 = n8314 ^ n8172 ^ 1'b0 ;
  assign n8316 = ( n7947 & n8314 ) | ( n7947 & n8315 ) | ( n8314 & n8315 ) ;
  assign n8317 = n8103 ^ n8044 ^ x70 ;
  assign n8318 = n8317 ^ n8172 ^ 1'b0 ;
  assign n8319 = ( n8044 & n8317 ) | ( n8044 & n8318 ) | ( n8317 & n8318 ) ;
  assign n8320 = n8102 ^ n7966 ^ x69 ;
  assign n8321 = n8320 ^ n8172 ^ 1'b0 ;
  assign n8322 = ( n7966 & n8320 ) | ( n7966 & n8321 ) | ( n8320 & n8321 ) ;
  assign n8323 = n8170 ^ n7967 ^ x121 ;
  assign n8324 = n8323 ^ n8172 ^ 1'b0 ;
  assign n8325 = ( n7967 & n8323 ) | ( n7967 & n8324 ) | ( n8323 & n8324 ) ;
  assign n8326 = ~x5 & x64 ;
  assign n8327 = ~n155 & n8096 ;
  assign n8328 = n8171 | n8327 ;
  assign n8329 = ( x6 & ~n8171 ) | ( x6 & n8328 ) | ( ~n8171 & n8328 ) ;
  assign n8330 = x123 | n154 ;
  assign n8331 = x64 & ~x122 ;
  assign n8332 = ~n8330 & n8331 ;
  assign n8333 = n8329 & ~n8332 ;
  assign n8334 = ( n8328 & n8329 ) | ( n8328 & n8333 ) | ( n8329 & n8333 ) ;
  assign n8335 = n8334 ^ n8326 ^ x65 ;
  assign n8336 = ( x65 & n8326 ) | ( x65 & n8335 ) | ( n8326 & n8335 ) ;
  assign n8337 = n8336 ^ n8201 ^ x66 ;
  assign n8338 = ( x66 & n8336 ) | ( x66 & n8337 ) | ( n8336 & n8337 ) ;
  assign n8339 = ( x67 & ~n8178 ) | ( x67 & n8338 ) | ( ~n8178 & n8338 ) ;
  assign n8340 = ( x68 & ~n8192 ) | ( x68 & n8339 ) | ( ~n8192 & n8339 ) ;
  assign n8341 = ( x69 & ~n8198 ) | ( x69 & n8340 ) | ( ~n8198 & n8340 ) ;
  assign n8342 = ( x70 & ~n8322 ) | ( x70 & n8341 ) | ( ~n8322 & n8341 ) ;
  assign n8343 = ( x71 & ~n8319 ) | ( x71 & n8342 ) | ( ~n8319 & n8342 ) ;
  assign n8344 = ( x72 & ~n8316 ) | ( x72 & n8343 ) | ( ~n8316 & n8343 ) ;
  assign n8345 = ( x73 & ~n8313 ) | ( x73 & n8344 ) | ( ~n8313 & n8344 ) ;
  assign n8346 = ( x74 & ~n8182 ) | ( x74 & n8345 ) | ( ~n8182 & n8345 ) ;
  assign n8347 = ( x75 & ~n8277 ) | ( x75 & n8346 ) | ( ~n8277 & n8346 ) ;
  assign n8348 = ( x76 & ~n8205 ) | ( x76 & n8347 ) | ( ~n8205 & n8347 ) ;
  assign n8349 = ( x77 & ~n8274 ) | ( x77 & n8348 ) | ( ~n8274 & n8348 ) ;
  assign n8350 = ( x78 & ~n8203 ) | ( x78 & n8349 ) | ( ~n8203 & n8349 ) ;
  assign n8351 = ( x79 & ~n8181 ) | ( x79 & n8350 ) | ( ~n8181 & n8350 ) ;
  assign n8352 = ( x80 & ~n8271 ) | ( x80 & n8351 ) | ( ~n8271 & n8351 ) ;
  assign n8353 = ( x81 & ~n8190 ) | ( x81 & n8352 ) | ( ~n8190 & n8352 ) ;
  assign n8354 = ( x82 & ~n8310 ) | ( x82 & n8353 ) | ( ~n8310 & n8353 ) ;
  assign n8355 = ( x83 & ~n8307 ) | ( x83 & n8354 ) | ( ~n8307 & n8354 ) ;
  assign n8356 = ( x84 & ~n8196 ) | ( x84 & n8355 ) | ( ~n8196 & n8355 ) ;
  assign n8357 = ( x85 & ~n8209 ) | ( x85 & n8356 ) | ( ~n8209 & n8356 ) ;
  assign n8358 = ( x86 & ~n8304 ) | ( x86 & n8357 ) | ( ~n8304 & n8357 ) ;
  assign n8359 = n8346 ^ n8277 ^ x75 ;
  assign n8360 = n8347 ^ n8205 ^ x76 ;
  assign n8361 = n8348 ^ n8274 ^ x77 ;
  assign n8362 = n8349 ^ n8203 ^ x78 ;
  assign n8363 = n8350 ^ n8181 ^ x79 ;
  assign n8364 = ( x87 & ~n8217 ) | ( x87 & n8358 ) | ( ~n8217 & n8358 ) ;
  assign n8365 = n8352 ^ n8190 ^ x81 ;
  assign n8366 = n8353 ^ n8310 ^ x82 ;
  assign n8367 = n8354 ^ n8307 ^ x83 ;
  assign n8368 = n8355 ^ n8196 ^ x84 ;
  assign n8369 = n8356 ^ n8209 ^ x85 ;
  assign n8370 = ( x88 & ~n8219 ) | ( x88 & n8364 ) | ( ~n8219 & n8364 ) ;
  assign n8371 = ( x89 & ~n8186 ) | ( x89 & n8370 ) | ( ~n8186 & n8370 ) ;
  assign n8372 = ( x90 & ~n8268 ) | ( x90 & n8371 ) | ( ~n8268 & n8371 ) ;
  assign n8373 = ( x91 & ~n8301 ) | ( x91 & n8372 ) | ( ~n8301 & n8372 ) ;
  assign n8374 = ( x92 & ~n8265 ) | ( x92 & n8373 ) | ( ~n8265 & n8373 ) ;
  assign n8375 = ( x93 & ~n8220 ) | ( x93 & n8374 ) | ( ~n8220 & n8374 ) ;
  assign n8376 = ( x94 & ~n8195 ) | ( x94 & n8375 ) | ( ~n8195 & n8375 ) ;
  assign n8377 = ( x95 & ~n8298 ) | ( x95 & n8376 ) | ( ~n8298 & n8376 ) ;
  assign n8378 = ( x96 & ~n8295 ) | ( x96 & n8377 ) | ( ~n8295 & n8377 ) ;
  assign n8379 = ( x97 & ~n8260 ) | ( x97 & n8378 ) | ( ~n8260 & n8378 ) ;
  assign n8380 = ( x98 & ~n8292 ) | ( x98 & n8379 ) | ( ~n8292 & n8379 ) ;
  assign n8381 = ( x99 & ~n8175 ) | ( x99 & n8380 ) | ( ~n8175 & n8380 ) ;
  assign n8382 = ( x100 & ~n8257 ) | ( x100 & n8381 ) | ( ~n8257 & n8381 ) ;
  assign n8383 = n155 & n8325 ;
  assign n8384 = n8357 ^ n8304 ^ x86 ;
  assign n8385 = n155 & n7967 ;
  assign n8386 = ( x101 & ~n8289 ) | ( x101 & n8382 ) | ( ~n8289 & n8382 ) ;
  assign n8387 = ( x102 & ~n8216 ) | ( x102 & n8386 ) | ( ~n8216 & n8386 ) ;
  assign n8388 = ( x103 & ~n8254 ) | ( x103 & n8387 ) | ( ~n8254 & n8387 ) ;
  assign n8389 = ( x104 & ~n8286 ) | ( x104 & n8388 ) | ( ~n8286 & n8388 ) ;
  assign n8390 = ( x105 & ~n8251 ) | ( x105 & n8389 ) | ( ~n8251 & n8389 ) ;
  assign n8391 = ( x106 & ~n8202 ) | ( x106 & n8390 ) | ( ~n8202 & n8390 ) ;
  assign n8392 = ( x107 & ~n8214 ) | ( x107 & n8391 ) | ( ~n8214 & n8391 ) ;
  assign n8393 = ( x108 & ~n8218 ) | ( x108 & n8392 ) | ( ~n8218 & n8392 ) ;
  assign n8394 = ( x109 & ~n8213 ) | ( x109 & n8393 ) | ( ~n8213 & n8393 ) ;
  assign n8395 = ( x110 & ~n8248 ) | ( x110 & n8394 ) | ( ~n8248 & n8394 ) ;
  assign n8396 = ( x111 & ~n8262 ) | ( x111 & n8395 ) | ( ~n8262 & n8395 ) ;
  assign n8397 = ( x112 & ~n8244 ) | ( x112 & n8396 ) | ( ~n8244 & n8396 ) ;
  assign n8398 = ( x113 & ~n8241 ) | ( x113 & n8397 ) | ( ~n8241 & n8397 ) ;
  assign n8399 = ( x114 & ~n8238 ) | ( x114 & n8398 ) | ( ~n8238 & n8398 ) ;
  assign n8400 = ( x115 & ~n8235 ) | ( x115 & n8399 ) | ( ~n8235 & n8399 ) ;
  assign n8401 = ( x116 & ~n8232 ) | ( x116 & n8400 ) | ( ~n8232 & n8400 ) ;
  assign n8402 = ( x117 & ~n8229 ) | ( x117 & n8401 ) | ( ~n8229 & n8401 ) ;
  assign n8403 = ( x118 & ~n8283 ) | ( x118 & n8402 ) | ( ~n8283 & n8402 ) ;
  assign n8404 = ( x119 & ~n8226 ) | ( x119 & n8403 ) | ( ~n8226 & n8403 ) ;
  assign n8405 = ( x120 & ~n8280 ) | ( x120 & n8404 ) | ( ~n8280 & n8404 ) ;
  assign n8406 = ( x122 & ~n8325 ) | ( x122 & n8330 ) | ( ~n8325 & n8330 ) ;
  assign n8407 = ( x121 & ~n8223 ) | ( x121 & n8405 ) | ( ~n8223 & n8405 ) ;
  assign n8408 = ( ~x122 & n8325 ) | ( ~x122 & n8407 ) | ( n8325 & n8407 ) ;
  assign n8409 = n8406 | n8408 ;
  assign n8410 = ( ~n8325 & n8383 ) | ( ~n8325 & n8409 ) | ( n8383 & n8409 ) ;
  assign n8411 = n8404 ^ n8280 ^ x120 ;
  assign n8412 = n8410 ^ n8280 ^ 1'b0 ;
  assign n8413 = ( n8280 & n8411 ) | ( n8280 & ~n8412 ) | ( n8411 & ~n8412 ) ;
  assign n8414 = n8403 ^ n8226 ^ x119 ;
  assign n8415 = n8410 ^ n8226 ^ 1'b0 ;
  assign n8416 = ( n8226 & n8414 ) | ( n8226 & ~n8415 ) | ( n8414 & ~n8415 ) ;
  assign n8417 = n8402 ^ n8283 ^ x118 ;
  assign n8418 = n8410 ^ n8283 ^ 1'b0 ;
  assign n8419 = ( n8283 & n8417 ) | ( n8283 & ~n8418 ) | ( n8417 & ~n8418 ) ;
  assign n8420 = n8410 ^ n8229 ^ 1'b0 ;
  assign n8421 = n8400 ^ n8232 ^ x116 ;
  assign n8422 = n8410 ^ n8232 ^ 1'b0 ;
  assign n8423 = n8401 ^ n8229 ^ x117 ;
  assign n8424 = ( n8229 & ~n8420 ) | ( n8229 & n8423 ) | ( ~n8420 & n8423 ) ;
  assign n8425 = ( n8232 & n8421 ) | ( n8232 & ~n8422 ) | ( n8421 & ~n8422 ) ;
  assign n8426 = n8399 ^ n8235 ^ x115 ;
  assign n8427 = n8410 ^ n8235 ^ 1'b0 ;
  assign n8428 = ( n8235 & n8426 ) | ( n8235 & ~n8427 ) | ( n8426 & ~n8427 ) ;
  assign n8429 = n8410 ^ n8304 ^ 1'b0 ;
  assign n8430 = ( n8304 & n8384 ) | ( n8304 & ~n8429 ) | ( n8384 & ~n8429 ) ;
  assign n8431 = n8410 ^ n8209 ^ 1'b0 ;
  assign n8432 = ( n8209 & n8369 ) | ( n8209 & ~n8431 ) | ( n8369 & ~n8431 ) ;
  assign n8433 = n8410 ^ n8196 ^ 1'b0 ;
  assign n8434 = ( n8196 & n8368 ) | ( n8196 & ~n8433 ) | ( n8368 & ~n8433 ) ;
  assign n8435 = n8410 ^ n8307 ^ 1'b0 ;
  assign n8436 = ( n8307 & n8367 ) | ( n8307 & ~n8435 ) | ( n8367 & ~n8435 ) ;
  assign n8437 = n8410 ^ n8310 ^ 1'b0 ;
  assign n8438 = ( n8310 & n8366 ) | ( n8310 & ~n8437 ) | ( n8366 & ~n8437 ) ;
  assign n8439 = n8410 ^ n8190 ^ 1'b0 ;
  assign n8440 = ( n8190 & n8365 ) | ( n8190 & ~n8439 ) | ( n8365 & ~n8439 ) ;
  assign n8441 = n8410 ^ n8181 ^ 1'b0 ;
  assign n8442 = ( n8181 & n8363 ) | ( n8181 & ~n8441 ) | ( n8363 & ~n8441 ) ;
  assign n8443 = n8410 ^ n8203 ^ 1'b0 ;
  assign n8444 = ( n8203 & n8362 ) | ( n8203 & ~n8443 ) | ( n8362 & ~n8443 ) ;
  assign n8445 = n8410 ^ n8274 ^ 1'b0 ;
  assign n8446 = ( n8274 & n8361 ) | ( n8274 & ~n8445 ) | ( n8361 & ~n8445 ) ;
  assign n8447 = n8410 ^ n8205 ^ 1'b0 ;
  assign n8448 = ( n8205 & n8360 ) | ( n8205 & ~n8447 ) | ( n8360 & ~n8447 ) ;
  assign n8449 = n8410 ^ n8277 ^ 1'b0 ;
  assign n8450 = ( n8277 & n8359 ) | ( n8277 & ~n8449 ) | ( n8359 & ~n8449 ) ;
  assign n8451 = n8410 ^ n8337 ^ 1'b0 ;
  assign n8452 = ( n8201 & n8337 ) | ( n8201 & n8451 ) | ( n8337 & n8451 ) ;
  assign n8453 = n8410 ^ n8335 ^ 1'b0 ;
  assign n8454 = ( n8334 & n8335 ) | ( n8334 & n8453 ) | ( n8335 & n8453 ) ;
  assign n8455 = n8407 ^ n8325 ^ x122 ;
  assign n8456 = ~n8410 & n8455 ;
  assign n8457 = n8385 & ~n8409 ;
  assign n8458 = ( n8385 & n8456 ) | ( n8385 & ~n8457 ) | ( n8456 & ~n8457 ) ;
  assign n8459 = n8405 ^ n8223 ^ x121 ;
  assign n8460 = n8410 ^ n8223 ^ 1'b0 ;
  assign n8461 = ( n8223 & n8459 ) | ( n8223 & ~n8460 ) | ( n8459 & ~n8460 ) ;
  assign n8462 = n8398 ^ n8238 ^ x114 ;
  assign n8463 = n8410 ^ n8238 ^ 1'b0 ;
  assign n8464 = ( n8238 & n8462 ) | ( n8238 & ~n8463 ) | ( n8462 & ~n8463 ) ;
  assign n8465 = n8376 ^ n8298 ^ x95 ;
  assign n8466 = n8410 ^ n8298 ^ 1'b0 ;
  assign n8467 = ( n8298 & n8465 ) | ( n8298 & ~n8466 ) | ( n8465 & ~n8466 ) ;
  assign n8468 = n8375 ^ n8195 ^ x94 ;
  assign n8469 = n8410 ^ n8195 ^ 1'b0 ;
  assign n8470 = ( n8195 & n8468 ) | ( n8195 & ~n8469 ) | ( n8468 & ~n8469 ) ;
  assign n8471 = n8374 ^ n8220 ^ x93 ;
  assign n8472 = n8410 ^ n8220 ^ 1'b0 ;
  assign n8473 = ( n8220 & n8471 ) | ( n8220 & ~n8472 ) | ( n8471 & ~n8472 ) ;
  assign n8474 = n8373 ^ n8265 ^ x92 ;
  assign n8475 = n8410 ^ n8265 ^ 1'b0 ;
  assign n8476 = ( n8265 & n8474 ) | ( n8265 & ~n8475 ) | ( n8474 & ~n8475 ) ;
  assign n8477 = n8372 ^ n8301 ^ x91 ;
  assign n8478 = n8410 ^ n8301 ^ 1'b0 ;
  assign n8479 = ( n8301 & n8477 ) | ( n8301 & ~n8478 ) | ( n8477 & ~n8478 ) ;
  assign n8480 = n8371 ^ n8268 ^ x90 ;
  assign n8481 = n8410 ^ n8268 ^ 1'b0 ;
  assign n8482 = ( n8268 & n8480 ) | ( n8268 & ~n8481 ) | ( n8480 & ~n8481 ) ;
  assign n8483 = n8370 ^ n8186 ^ x89 ;
  assign n8484 = n8410 ^ n8186 ^ 1'b0 ;
  assign n8485 = ( n8186 & n8483 ) | ( n8186 & ~n8484 ) | ( n8483 & ~n8484 ) ;
  assign n8486 = n8364 ^ n8219 ^ x88 ;
  assign n8487 = n8410 ^ n8219 ^ 1'b0 ;
  assign n8488 = ( n8219 & n8486 ) | ( n8219 & ~n8487 ) | ( n8486 & ~n8487 ) ;
  assign n8489 = n8358 ^ n8217 ^ x87 ;
  assign n8490 = n8410 ^ n8217 ^ 1'b0 ;
  assign n8491 = ( n8217 & n8489 ) | ( n8217 & ~n8490 ) | ( n8489 & ~n8490 ) ;
  assign n8492 = n8351 ^ n8271 ^ x80 ;
  assign n8493 = n8410 ^ n8271 ^ 1'b0 ;
  assign n8494 = ( n8271 & n8492 ) | ( n8271 & ~n8493 ) | ( n8492 & ~n8493 ) ;
  assign n8495 = n8345 ^ n8182 ^ x74 ;
  assign n8496 = n8410 ^ n8182 ^ 1'b0 ;
  assign n8497 = ( n8182 & n8495 ) | ( n8182 & ~n8496 ) | ( n8495 & ~n8496 ) ;
  assign n8498 = n8344 ^ n8313 ^ x73 ;
  assign n8499 = n8410 ^ n8313 ^ 1'b0 ;
  assign n8500 = ( n8313 & n8498 ) | ( n8313 & ~n8499 ) | ( n8498 & ~n8499 ) ;
  assign n8501 = n8343 ^ n8316 ^ x72 ;
  assign n8502 = n8410 ^ n8316 ^ 1'b0 ;
  assign n8503 = ( n8316 & n8501 ) | ( n8316 & ~n8502 ) | ( n8501 & ~n8502 ) ;
  assign n8504 = n8342 ^ n8319 ^ x71 ;
  assign n8505 = n8410 ^ n8319 ^ 1'b0 ;
  assign n8506 = ( n8319 & n8504 ) | ( n8319 & ~n8505 ) | ( n8504 & ~n8505 ) ;
  assign n8507 = n8341 ^ n8322 ^ x70 ;
  assign n8508 = n8410 ^ n8322 ^ 1'b0 ;
  assign n8509 = ( n8322 & n8507 ) | ( n8322 & ~n8508 ) | ( n8507 & ~n8508 ) ;
  assign n8510 = n8340 ^ n8198 ^ x69 ;
  assign n8511 = n8410 ^ n8198 ^ 1'b0 ;
  assign n8512 = ( n8198 & n8510 ) | ( n8198 & ~n8511 ) | ( n8510 & ~n8511 ) ;
  assign n8513 = n8339 ^ n8192 ^ x68 ;
  assign n8514 = n8410 ^ n8192 ^ 1'b0 ;
  assign n8515 = ( n8192 & n8513 ) | ( n8192 & ~n8514 ) | ( n8513 & ~n8514 ) ;
  assign n8516 = n8338 ^ n8178 ^ x67 ;
  assign n8517 = n8410 ^ n8178 ^ 1'b0 ;
  assign n8518 = ( n8178 & n8516 ) | ( n8178 & ~n8517 ) | ( n8516 & ~n8517 ) ;
  assign n8519 = n8397 ^ n8241 ^ x113 ;
  assign n8520 = n8410 ^ n8241 ^ 1'b0 ;
  assign n8521 = ( n8241 & n8519 ) | ( n8241 & ~n8520 ) | ( n8519 & ~n8520 ) ;
  assign n8522 = n8396 ^ n8244 ^ x112 ;
  assign n8523 = n8410 ^ n8244 ^ 1'b0 ;
  assign n8524 = ( n8244 & n8522 ) | ( n8244 & ~n8523 ) | ( n8522 & ~n8523 ) ;
  assign n8525 = n8395 ^ n8262 ^ x111 ;
  assign n8526 = n8410 ^ n8262 ^ 1'b0 ;
  assign n8527 = ( n8262 & n8525 ) | ( n8262 & ~n8526 ) | ( n8525 & ~n8526 ) ;
  assign n8528 = n8394 ^ n8248 ^ x110 ;
  assign n8529 = n8410 ^ n8248 ^ 1'b0 ;
  assign n8530 = ( n8248 & n8528 ) | ( n8248 & ~n8529 ) | ( n8528 & ~n8529 ) ;
  assign n8531 = n8393 ^ n8213 ^ x109 ;
  assign n8532 = n8410 ^ n8213 ^ 1'b0 ;
  assign n8533 = ( n8213 & n8531 ) | ( n8213 & ~n8532 ) | ( n8531 & ~n8532 ) ;
  assign n8534 = n8392 ^ n8218 ^ x108 ;
  assign n8535 = n8410 ^ n8218 ^ 1'b0 ;
  assign n8536 = ( n8218 & n8534 ) | ( n8218 & ~n8535 ) | ( n8534 & ~n8535 ) ;
  assign n8537 = n8391 ^ n8214 ^ x107 ;
  assign n8538 = n8410 ^ n8214 ^ 1'b0 ;
  assign n8539 = ( n8214 & n8537 ) | ( n8214 & ~n8538 ) | ( n8537 & ~n8538 ) ;
  assign n8540 = n8390 ^ n8202 ^ x106 ;
  assign n8541 = n8410 ^ n8202 ^ 1'b0 ;
  assign n8542 = ( n8202 & n8540 ) | ( n8202 & ~n8541 ) | ( n8540 & ~n8541 ) ;
  assign n8543 = n8389 ^ n8251 ^ x105 ;
  assign n8544 = n8410 ^ n8251 ^ 1'b0 ;
  assign n8545 = ( n8251 & n8543 ) | ( n8251 & ~n8544 ) | ( n8543 & ~n8544 ) ;
  assign n8546 = n8388 ^ n8286 ^ x104 ;
  assign n8547 = n8410 ^ n8286 ^ 1'b0 ;
  assign n8548 = ( n8286 & n8546 ) | ( n8286 & ~n8547 ) | ( n8546 & ~n8547 ) ;
  assign n8549 = n8387 ^ n8254 ^ x103 ;
  assign n8550 = n8410 ^ n8254 ^ 1'b0 ;
  assign n8551 = ( n8254 & n8549 ) | ( n8254 & ~n8550 ) | ( n8549 & ~n8550 ) ;
  assign n8552 = n8386 ^ n8216 ^ x102 ;
  assign n8553 = n8410 ^ n8216 ^ 1'b0 ;
  assign n8554 = ( n8216 & n8552 ) | ( n8216 & ~n8553 ) | ( n8552 & ~n8553 ) ;
  assign n8555 = n8382 ^ n8289 ^ x101 ;
  assign n8556 = n8410 ^ n8289 ^ 1'b0 ;
  assign n8557 = ( n8289 & n8555 ) | ( n8289 & ~n8556 ) | ( n8555 & ~n8556 ) ;
  assign n8558 = n8381 ^ n8257 ^ x100 ;
  assign n8559 = n8410 ^ n8257 ^ 1'b0 ;
  assign n8560 = ( n8257 & n8558 ) | ( n8257 & ~n8559 ) | ( n8558 & ~n8559 ) ;
  assign n8561 = n8380 ^ n8175 ^ x99 ;
  assign n8562 = n8410 ^ n8175 ^ 1'b0 ;
  assign n8563 = ( n8175 & n8561 ) | ( n8175 & ~n8562 ) | ( n8561 & ~n8562 ) ;
  assign n8564 = n8379 ^ n8292 ^ x98 ;
  assign n8565 = n8410 ^ n8292 ^ 1'b0 ;
  assign n8566 = ( n8292 & n8564 ) | ( n8292 & ~n8565 ) | ( n8564 & ~n8565 ) ;
  assign n8567 = n8378 ^ n8260 ^ x97 ;
  assign n8568 = n8410 ^ n8260 ^ 1'b0 ;
  assign n8569 = ( n8260 & n8567 ) | ( n8260 & ~n8568 ) | ( n8567 & ~n8568 ) ;
  assign n8570 = n8377 ^ n8295 ^ x96 ;
  assign n8571 = n8410 ^ n8295 ^ 1'b0 ;
  assign n8572 = ( n8295 & n8570 ) | ( n8295 & ~n8571 ) | ( n8570 & ~n8571 ) ;
  assign n8573 = x64 & n8410 ;
  assign n8574 = n8573 ^ x64 ^ x5 ;
  assign n8575 = ~x4 & x64 ;
  assign n8576 = n8575 ^ n8574 ^ x65 ;
  assign n8577 = ( x65 & n8575 ) | ( x65 & n8576 ) | ( n8575 & n8576 ) ;
  assign n8578 = n8577 ^ n8454 ^ x66 ;
  assign n8579 = ( x66 & n8577 ) | ( x66 & n8578 ) | ( n8577 & n8578 ) ;
  assign n8580 = ( x67 & ~n8452 ) | ( x67 & n8579 ) | ( ~n8452 & n8579 ) ;
  assign n8581 = ( x68 & ~n8518 ) | ( x68 & n8580 ) | ( ~n8518 & n8580 ) ;
  assign n8582 = ( x69 & ~n8515 ) | ( x69 & n8581 ) | ( ~n8515 & n8581 ) ;
  assign n8583 = ( x70 & ~n8512 ) | ( x70 & n8582 ) | ( ~n8512 & n8582 ) ;
  assign n8584 = ( x71 & ~n8509 ) | ( x71 & n8583 ) | ( ~n8509 & n8583 ) ;
  assign n8585 = ( x72 & ~n8506 ) | ( x72 & n8584 ) | ( ~n8506 & n8584 ) ;
  assign n8586 = ( x73 & ~n8503 ) | ( x73 & n8585 ) | ( ~n8503 & n8585 ) ;
  assign n8587 = ( x74 & ~n8500 ) | ( x74 & n8586 ) | ( ~n8500 & n8586 ) ;
  assign n8588 = ( x75 & ~n8497 ) | ( x75 & n8587 ) | ( ~n8497 & n8587 ) ;
  assign n8589 = ( x76 & ~n8450 ) | ( x76 & n8588 ) | ( ~n8450 & n8588 ) ;
  assign n8590 = ( x77 & ~n8448 ) | ( x77 & n8589 ) | ( ~n8448 & n8589 ) ;
  assign n8591 = ( x78 & ~n8446 ) | ( x78 & n8590 ) | ( ~n8446 & n8590 ) ;
  assign n8592 = ( x79 & ~n8444 ) | ( x79 & n8591 ) | ( ~n8444 & n8591 ) ;
  assign n8593 = ( x80 & ~n8442 ) | ( x80 & n8592 ) | ( ~n8442 & n8592 ) ;
  assign n8594 = ( x81 & ~n8494 ) | ( x81 & n8593 ) | ( ~n8494 & n8593 ) ;
  assign n8595 = ( x82 & ~n8440 ) | ( x82 & n8594 ) | ( ~n8440 & n8594 ) ;
  assign n8596 = ( x83 & ~n8438 ) | ( x83 & n8595 ) | ( ~n8438 & n8595 ) ;
  assign n8597 = ( x84 & ~n8436 ) | ( x84 & n8596 ) | ( ~n8436 & n8596 ) ;
  assign n8598 = ( x85 & ~n8434 ) | ( x85 & n8597 ) | ( ~n8434 & n8597 ) ;
  assign n8599 = ( x86 & ~n8432 ) | ( x86 & n8598 ) | ( ~n8432 & n8598 ) ;
  assign n8600 = ( x87 & ~n8430 ) | ( x87 & n8599 ) | ( ~n8430 & n8599 ) ;
  assign n8601 = ( x88 & ~n8491 ) | ( x88 & n8600 ) | ( ~n8491 & n8600 ) ;
  assign n8602 = ( x89 & ~n8488 ) | ( x89 & n8601 ) | ( ~n8488 & n8601 ) ;
  assign n8603 = ( x90 & ~n8485 ) | ( x90 & n8602 ) | ( ~n8485 & n8602 ) ;
  assign n8604 = ( x91 & ~n8482 ) | ( x91 & n8603 ) | ( ~n8482 & n8603 ) ;
  assign n8605 = ( x92 & ~n8479 ) | ( x92 & n8604 ) | ( ~n8479 & n8604 ) ;
  assign n8606 = ( x93 & ~n8476 ) | ( x93 & n8605 ) | ( ~n8476 & n8605 ) ;
  assign n8607 = ( x94 & ~n8473 ) | ( x94 & n8606 ) | ( ~n8473 & n8606 ) ;
  assign n8608 = ( x95 & ~n8470 ) | ( x95 & n8607 ) | ( ~n8470 & n8607 ) ;
  assign n8609 = ( x96 & ~n8467 ) | ( x96 & n8608 ) | ( ~n8467 & n8608 ) ;
  assign n8610 = ( x97 & ~n8572 ) | ( x97 & n8609 ) | ( ~n8572 & n8609 ) ;
  assign n8611 = ( x98 & ~n8569 ) | ( x98 & n8610 ) | ( ~n8569 & n8610 ) ;
  assign n8612 = ( x99 & ~n8566 ) | ( x99 & n8611 ) | ( ~n8566 & n8611 ) ;
  assign n8613 = ( x100 & ~n8563 ) | ( x100 & n8612 ) | ( ~n8563 & n8612 ) ;
  assign n8614 = ( x101 & ~n8560 ) | ( x101 & n8613 ) | ( ~n8560 & n8613 ) ;
  assign n8615 = ( x102 & ~n8557 ) | ( x102 & n8614 ) | ( ~n8557 & n8614 ) ;
  assign n8616 = ( x103 & ~n8554 ) | ( x103 & n8615 ) | ( ~n8554 & n8615 ) ;
  assign n8617 = ( x104 & ~n8551 ) | ( x104 & n8616 ) | ( ~n8551 & n8616 ) ;
  assign n8618 = ( x105 & ~n8548 ) | ( x105 & n8617 ) | ( ~n8548 & n8617 ) ;
  assign n8619 = n8607 ^ n8470 ^ x95 ;
  assign n8620 = ( x106 & ~n8545 ) | ( x106 & n8618 ) | ( ~n8545 & n8618 ) ;
  assign n8621 = n8589 ^ n8448 ^ x77 ;
  assign n8622 = n8610 ^ n8569 ^ x98 ;
  assign n8623 = n8620 ^ n8542 ^ x107 ;
  assign n8624 = n8604 ^ n8479 ^ x92 ;
  assign n8625 = n8598 ^ n8432 ^ x86 ;
  assign n8626 = n8592 ^ n8442 ^ x80 ;
  assign n8627 = n8618 ^ n8545 ^ x106 ;
  assign n8628 = n8590 ^ n8446 ^ x78 ;
  assign n8629 = ( x107 & ~n8542 ) | ( x107 & n8620 ) | ( ~n8542 & n8620 ) ;
  assign n8630 = n8330 & n8458 ;
  assign n8631 = n8587 ^ n8497 ^ x75 ;
  assign n8632 = n8579 ^ n8452 ^ x67 ;
  assign n8633 = ( x108 & ~n8539 ) | ( x108 & n8629 ) | ( ~n8539 & n8629 ) ;
  assign n8634 = ( x109 & ~n8536 ) | ( x109 & n8633 ) | ( ~n8536 & n8633 ) ;
  assign n8635 = ( x110 & ~n8533 ) | ( x110 & n8634 ) | ( ~n8533 & n8634 ) ;
  assign n8636 = ( x111 & ~n8530 ) | ( x111 & n8635 ) | ( ~n8530 & n8635 ) ;
  assign n8637 = ( x112 & ~n8527 ) | ( x112 & n8636 ) | ( ~n8527 & n8636 ) ;
  assign n8638 = ( x113 & ~n8524 ) | ( x113 & n8637 ) | ( ~n8524 & n8637 ) ;
  assign n8639 = ( x114 & ~n8521 ) | ( x114 & n8638 ) | ( ~n8521 & n8638 ) ;
  assign n8640 = ( x115 & ~n8464 ) | ( x115 & n8639 ) | ( ~n8464 & n8639 ) ;
  assign n8641 = ( x116 & ~n8428 ) | ( x116 & n8640 ) | ( ~n8428 & n8640 ) ;
  assign n8642 = ( x117 & ~n8425 ) | ( x117 & n8641 ) | ( ~n8425 & n8641 ) ;
  assign n8643 = ( x118 & ~n8424 ) | ( x118 & n8642 ) | ( ~n8424 & n8642 ) ;
  assign n8644 = n8639 ^ n8464 ^ x115 ;
  assign n8645 = ( x119 & ~n8419 ) | ( x119 & n8643 ) | ( ~n8419 & n8643 ) ;
  assign n8646 = ( x120 & ~n8416 ) | ( x120 & n8645 ) | ( ~n8416 & n8645 ) ;
  assign n8647 = ( x123 & n154 ) | ( x123 & ~n8458 ) | ( n154 & ~n8458 ) ;
  assign n8648 = ( x121 & ~n8413 ) | ( x121 & n8646 ) | ( ~n8413 & n8646 ) ;
  assign n8649 = ( x122 & ~n8461 ) | ( x122 & n8648 ) | ( ~n8461 & n8648 ) ;
  assign n8650 = ( ~x123 & n8458 ) | ( ~x123 & n8649 ) | ( n8458 & n8649 ) ;
  assign n8651 = n8647 | n8650 ;
  assign n8652 = n8630 & ~n8651 ;
  assign n8653 = ( ~n8458 & n8630 ) | ( ~n8458 & n8651 ) | ( n8630 & n8651 ) ;
  assign n8654 = n8641 ^ n8425 ^ x117 ;
  assign n8655 = n8649 ^ n8458 ^ x123 ;
  assign n8656 = n8653 ^ n8425 ^ 1'b0 ;
  assign n8657 = n8645 ^ n8416 ^ x120 ;
  assign n8658 = ( n8425 & n8654 ) | ( n8425 & ~n8656 ) | ( n8654 & ~n8656 ) ;
  assign n8659 = n8642 ^ n8424 ^ x118 ;
  assign n8660 = n8638 ^ n8521 ^ x114 ;
  assign n8661 = n8653 ^ n8470 ^ 1'b0 ;
  assign n8662 = n8653 ^ n8497 ^ 1'b0 ;
  assign n8663 = n8635 ^ n8530 ^ x111 ;
  assign n8664 = n8637 ^ n8524 ^ x113 ;
  assign n8665 = ( n8470 & n8619 ) | ( n8470 & ~n8661 ) | ( n8619 & ~n8661 ) ;
  assign n8666 = n8653 ^ n8542 ^ 1'b0 ;
  assign n8667 = n8653 ^ n8464 ^ 1'b0 ;
  assign n8668 = ( n8464 & n8644 ) | ( n8464 & ~n8667 ) | ( n8644 & ~n8667 ) ;
  assign n8669 = n8653 ^ n8424 ^ 1'b0 ;
  assign n8670 = n8643 ^ n8419 ^ x119 ;
  assign n8671 = ( n8497 & n8631 ) | ( n8497 & ~n8662 ) | ( n8631 & ~n8662 ) ;
  assign n8672 = n8653 ^ n8524 ^ 1'b0 ;
  assign n8673 = n8653 ^ n8545 ^ 1'b0 ;
  assign n8674 = n8653 ^ n8448 ^ 1'b0 ;
  assign n8675 = ( n8448 & n8621 ) | ( n8448 & ~n8674 ) | ( n8621 & ~n8674 ) ;
  assign n8676 = n8653 ^ n8416 ^ 1'b0 ;
  assign n8677 = ( n8542 & n8623 ) | ( n8542 & ~n8666 ) | ( n8623 & ~n8666 ) ;
  assign n8678 = n8653 ^ n8578 ^ 1'b0 ;
  assign n8679 = n8653 ^ n8452 ^ 1'b0 ;
  assign n8680 = n8653 ^ n8521 ^ 1'b0 ;
  assign n8681 = ( n8545 & n8627 ) | ( n8545 & ~n8673 ) | ( n8627 & ~n8673 ) ;
  assign n8682 = n8653 ^ n8530 ^ 1'b0 ;
  assign n8683 = ( n8452 & n8632 ) | ( n8452 & ~n8679 ) | ( n8632 & ~n8679 ) ;
  assign n8684 = ~n8653 & n8655 ;
  assign n8685 = n8653 ^ n8442 ^ 1'b0 ;
  assign n8686 = n8653 ^ n8432 ^ 1'b0 ;
  assign n8687 = ( n8530 & n8663 ) | ( n8530 & ~n8682 ) | ( n8663 & ~n8682 ) ;
  assign n8688 = ( n8424 & n8659 ) | ( n8424 & ~n8669 ) | ( n8659 & ~n8669 ) ;
  assign n8689 = n8653 ^ n8419 ^ 1'b0 ;
  assign n8690 = n8653 ^ n8479 ^ 1'b0 ;
  assign n8691 = n8653 ^ n8576 ^ 1'b0 ;
  assign n8692 = ( n8479 & n8624 ) | ( n8479 & ~n8690 ) | ( n8624 & ~n8690 ) ;
  assign n8693 = n8653 ^ n8446 ^ 1'b0 ;
  assign n8694 = ( n8446 & n8628 ) | ( n8446 & ~n8693 ) | ( n8628 & ~n8693 ) ;
  assign n8695 = n8653 ^ n8569 ^ 1'b0 ;
  assign n8696 = ( n8416 & n8657 ) | ( n8416 & ~n8676 ) | ( n8657 & ~n8676 ) ;
  assign n8697 = ( n8569 & n8622 ) | ( n8569 & ~n8695 ) | ( n8622 & ~n8695 ) ;
  assign n8698 = ( n8454 & n8578 ) | ( n8454 & n8678 ) | ( n8578 & n8678 ) ;
  assign n8699 = ( n8442 & n8626 ) | ( n8442 & ~n8685 ) | ( n8626 & ~n8685 ) ;
  assign n8700 = ( n8630 & ~n8652 ) | ( n8630 & n8684 ) | ( ~n8652 & n8684 ) ;
  assign n8701 = ( n8574 & n8576 ) | ( n8574 & n8691 ) | ( n8576 & n8691 ) ;
  assign n8702 = ( n8521 & n8660 ) | ( n8521 & ~n8680 ) | ( n8660 & ~n8680 ) ;
  assign n8703 = ( n8432 & n8625 ) | ( n8432 & ~n8686 ) | ( n8625 & ~n8686 ) ;
  assign n8704 = ( n8524 & n8664 ) | ( n8524 & ~n8672 ) | ( n8664 & ~n8672 ) ;
  assign n8705 = ( n8419 & n8670 ) | ( n8419 & ~n8689 ) | ( n8670 & ~n8689 ) ;
  assign n8706 = n8648 ^ n8461 ^ x122 ;
  assign n8707 = n8653 ^ n8461 ^ 1'b0 ;
  assign n8708 = ( n8461 & n8706 ) | ( n8461 & ~n8707 ) | ( n8706 & ~n8707 ) ;
  assign n8709 = n8646 ^ n8413 ^ x121 ;
  assign n8710 = n8653 ^ n8413 ^ 1'b0 ;
  assign n8711 = ( n8413 & n8709 ) | ( n8413 & ~n8710 ) | ( n8709 & ~n8710 ) ;
  assign n8712 = n8640 ^ n8428 ^ x116 ;
  assign n8713 = n8653 ^ n8428 ^ 1'b0 ;
  assign n8714 = ( n8428 & n8712 ) | ( n8428 & ~n8713 ) | ( n8712 & ~n8713 ) ;
  assign n8715 = n8601 ^ n8488 ^ x89 ;
  assign n8716 = n8653 ^ n8488 ^ 1'b0 ;
  assign n8717 = ( n8488 & n8715 ) | ( n8488 & ~n8716 ) | ( n8715 & ~n8716 ) ;
  assign n8718 = n8600 ^ n8491 ^ x88 ;
  assign n8719 = n8653 ^ n8491 ^ 1'b0 ;
  assign n8720 = ( n8491 & n8718 ) | ( n8491 & ~n8719 ) | ( n8718 & ~n8719 ) ;
  assign n8721 = n8599 ^ n8430 ^ x87 ;
  assign n8722 = n8653 ^ n8430 ^ 1'b0 ;
  assign n8723 = ( n8430 & n8721 ) | ( n8430 & ~n8722 ) | ( n8721 & ~n8722 ) ;
  assign n8724 = n8597 ^ n8434 ^ x85 ;
  assign n8725 = n8653 ^ n8434 ^ 1'b0 ;
  assign n8726 = ( n8434 & n8724 ) | ( n8434 & ~n8725 ) | ( n8724 & ~n8725 ) ;
  assign n8727 = n8596 ^ n8436 ^ x84 ;
  assign n8728 = n8653 ^ n8436 ^ 1'b0 ;
  assign n8729 = ( n8436 & n8727 ) | ( n8436 & ~n8728 ) | ( n8727 & ~n8728 ) ;
  assign n8730 = n8595 ^ n8438 ^ x83 ;
  assign n8731 = n8653 ^ n8438 ^ 1'b0 ;
  assign n8732 = ( n8438 & n8730 ) | ( n8438 & ~n8731 ) | ( n8730 & ~n8731 ) ;
  assign n8733 = n8594 ^ n8440 ^ x82 ;
  assign n8734 = n8653 ^ n8440 ^ 1'b0 ;
  assign n8735 = ( n8440 & n8733 ) | ( n8440 & ~n8734 ) | ( n8733 & ~n8734 ) ;
  assign n8736 = n8593 ^ n8494 ^ x81 ;
  assign n8737 = n8653 ^ n8494 ^ 1'b0 ;
  assign n8738 = ( n8494 & n8736 ) | ( n8494 & ~n8737 ) | ( n8736 & ~n8737 ) ;
  assign n8739 = n8591 ^ n8444 ^ x79 ;
  assign n8740 = n8653 ^ n8444 ^ 1'b0 ;
  assign n8741 = ( n8444 & n8739 ) | ( n8444 & ~n8740 ) | ( n8739 & ~n8740 ) ;
  assign n8742 = n8588 ^ n8450 ^ x76 ;
  assign n8743 = n8653 ^ n8450 ^ 1'b0 ;
  assign n8744 = ( n8450 & n8742 ) | ( n8450 & ~n8743 ) | ( n8742 & ~n8743 ) ;
  assign n8745 = n8586 ^ n8500 ^ x74 ;
  assign n8746 = n8653 ^ n8500 ^ 1'b0 ;
  assign n8747 = ( n8500 & n8745 ) | ( n8500 & ~n8746 ) | ( n8745 & ~n8746 ) ;
  assign n8748 = n8585 ^ n8503 ^ x73 ;
  assign n8749 = n8653 ^ n8503 ^ 1'b0 ;
  assign n8750 = ( n8503 & n8748 ) | ( n8503 & ~n8749 ) | ( n8748 & ~n8749 ) ;
  assign n8751 = n8584 ^ n8506 ^ x72 ;
  assign n8752 = n8653 ^ n8506 ^ 1'b0 ;
  assign n8753 = ( n8506 & n8751 ) | ( n8506 & ~n8752 ) | ( n8751 & ~n8752 ) ;
  assign n8754 = n8583 ^ n8509 ^ x71 ;
  assign n8755 = n8653 ^ n8509 ^ 1'b0 ;
  assign n8756 = ( n8509 & n8754 ) | ( n8509 & ~n8755 ) | ( n8754 & ~n8755 ) ;
  assign n8757 = n8582 ^ n8512 ^ x70 ;
  assign n8758 = n8653 ^ n8512 ^ 1'b0 ;
  assign n8759 = ( n8512 & n8757 ) | ( n8512 & ~n8758 ) | ( n8757 & ~n8758 ) ;
  assign n8760 = n8581 ^ n8515 ^ x69 ;
  assign n8761 = n8653 ^ n8515 ^ 1'b0 ;
  assign n8762 = ( n8515 & n8760 ) | ( n8515 & ~n8761 ) | ( n8760 & ~n8761 ) ;
  assign n8763 = n8580 ^ n8518 ^ x68 ;
  assign n8764 = n8653 ^ n8518 ^ 1'b0 ;
  assign n8765 = ( n8518 & n8763 ) | ( n8518 & ~n8764 ) | ( n8763 & ~n8764 ) ;
  assign n8766 = n8636 ^ n8527 ^ x112 ;
  assign n8767 = n8653 ^ n8527 ^ 1'b0 ;
  assign n8768 = ( n8527 & n8766 ) | ( n8527 & ~n8767 ) | ( n8766 & ~n8767 ) ;
  assign n8769 = n8634 ^ n8533 ^ x110 ;
  assign n8770 = n8653 ^ n8533 ^ 1'b0 ;
  assign n8771 = ( n8533 & n8769 ) | ( n8533 & ~n8770 ) | ( n8769 & ~n8770 ) ;
  assign n8772 = n8633 ^ n8536 ^ x109 ;
  assign n8773 = n8653 ^ n8536 ^ 1'b0 ;
  assign n8774 = ( n8536 & n8772 ) | ( n8536 & ~n8773 ) | ( n8772 & ~n8773 ) ;
  assign n8775 = n8629 ^ n8539 ^ x108 ;
  assign n8776 = n8653 ^ n8539 ^ 1'b0 ;
  assign n8777 = ( n8539 & n8775 ) | ( n8539 & ~n8776 ) | ( n8775 & ~n8776 ) ;
  assign n8778 = n8617 ^ n8548 ^ x105 ;
  assign n8779 = n8653 ^ n8548 ^ 1'b0 ;
  assign n8780 = ( n8548 & n8778 ) | ( n8548 & ~n8779 ) | ( n8778 & ~n8779 ) ;
  assign n8781 = n8616 ^ n8551 ^ x104 ;
  assign n8782 = n8653 ^ n8551 ^ 1'b0 ;
  assign n8783 = ( n8551 & n8781 ) | ( n8551 & ~n8782 ) | ( n8781 & ~n8782 ) ;
  assign n8784 = n8615 ^ n8554 ^ x103 ;
  assign n8785 = n8653 ^ n8554 ^ 1'b0 ;
  assign n8786 = ( n8554 & n8784 ) | ( n8554 & ~n8785 ) | ( n8784 & ~n8785 ) ;
  assign n8787 = n8614 ^ n8557 ^ x102 ;
  assign n8788 = n8653 ^ n8557 ^ 1'b0 ;
  assign n8789 = ( n8557 & n8787 ) | ( n8557 & ~n8788 ) | ( n8787 & ~n8788 ) ;
  assign n8790 = n8613 ^ n8560 ^ x101 ;
  assign n8791 = n8653 ^ n8560 ^ 1'b0 ;
  assign n8792 = ( n8560 & n8790 ) | ( n8560 & ~n8791 ) | ( n8790 & ~n8791 ) ;
  assign n8793 = n8612 ^ n8563 ^ x100 ;
  assign n8794 = n8653 ^ n8563 ^ 1'b0 ;
  assign n8795 = ( n8563 & n8793 ) | ( n8563 & ~n8794 ) | ( n8793 & ~n8794 ) ;
  assign n8796 = n8611 ^ n8566 ^ x99 ;
  assign n8797 = n8653 ^ n8566 ^ 1'b0 ;
  assign n8798 = ( n8566 & n8796 ) | ( n8566 & ~n8797 ) | ( n8796 & ~n8797 ) ;
  assign n8799 = n8609 ^ n8572 ^ x97 ;
  assign n8800 = n8653 ^ n8572 ^ 1'b0 ;
  assign n8801 = ( n8572 & n8799 ) | ( n8572 & ~n8800 ) | ( n8799 & ~n8800 ) ;
  assign n8802 = n8608 ^ n8467 ^ x96 ;
  assign n8803 = n8653 ^ n8467 ^ 1'b0 ;
  assign n8804 = ( n8467 & n8802 ) | ( n8467 & ~n8803 ) | ( n8802 & ~n8803 ) ;
  assign n8805 = n8606 ^ n8473 ^ x94 ;
  assign n8806 = n8653 ^ n8473 ^ 1'b0 ;
  assign n8807 = ( n8473 & n8805 ) | ( n8473 & ~n8806 ) | ( n8805 & ~n8806 ) ;
  assign n8808 = n8605 ^ n8476 ^ x93 ;
  assign n8809 = n8653 ^ n8476 ^ 1'b0 ;
  assign n8810 = ( n8476 & n8808 ) | ( n8476 & ~n8809 ) | ( n8808 & ~n8809 ) ;
  assign n8811 = n8603 ^ n8482 ^ x91 ;
  assign n8812 = n8653 ^ n8482 ^ 1'b0 ;
  assign n8813 = ( n8482 & n8811 ) | ( n8482 & ~n8812 ) | ( n8811 & ~n8812 ) ;
  assign n8814 = n8602 ^ n8485 ^ x90 ;
  assign n8815 = n8653 ^ n8485 ^ 1'b0 ;
  assign n8816 = ( n8485 & n8814 ) | ( n8485 & ~n8815 ) | ( n8814 & ~n8815 ) ;
  assign n8817 = ~x3 & x64 ;
  assign n8818 = x64 & n8653 ;
  assign n8819 = n8818 ^ x64 ^ x4 ;
  assign n8820 = n8819 ^ n8817 ^ x65 ;
  assign n8821 = ( x65 & n8817 ) | ( x65 & n8820 ) | ( n8817 & n8820 ) ;
  assign n8822 = n8821 ^ n8701 ^ x66 ;
  assign n8823 = ( x66 & n8821 ) | ( x66 & n8822 ) | ( n8821 & n8822 ) ;
  assign n8824 = ( x67 & ~n8698 ) | ( x67 & n8823 ) | ( ~n8698 & n8823 ) ;
  assign n8825 = ( x68 & ~n8683 ) | ( x68 & n8824 ) | ( ~n8683 & n8824 ) ;
  assign n8826 = ( x69 & ~n8765 ) | ( x69 & n8825 ) | ( ~n8765 & n8825 ) ;
  assign n8827 = ( x70 & ~n8762 ) | ( x70 & n8826 ) | ( ~n8762 & n8826 ) ;
  assign n8828 = ( x71 & ~n8759 ) | ( x71 & n8827 ) | ( ~n8759 & n8827 ) ;
  assign n8829 = ( x72 & ~n8756 ) | ( x72 & n8828 ) | ( ~n8756 & n8828 ) ;
  assign n8830 = ( x73 & ~n8753 ) | ( x73 & n8829 ) | ( ~n8753 & n8829 ) ;
  assign n8831 = ( x74 & ~n8750 ) | ( x74 & n8830 ) | ( ~n8750 & n8830 ) ;
  assign n8832 = ( x75 & ~n8747 ) | ( x75 & n8831 ) | ( ~n8747 & n8831 ) ;
  assign n8833 = n154 & n8700 ;
  assign n8834 = ( x76 & ~n8671 ) | ( x76 & n8832 ) | ( ~n8671 & n8832 ) ;
  assign n8835 = ( x77 & ~n8744 ) | ( x77 & n8834 ) | ( ~n8744 & n8834 ) ;
  assign n8836 = ( x78 & ~n8675 ) | ( x78 & n8835 ) | ( ~n8675 & n8835 ) ;
  assign n8837 = ( x79 & ~n8694 ) | ( x79 & n8836 ) | ( ~n8694 & n8836 ) ;
  assign n8838 = ( x80 & ~n8741 ) | ( x80 & n8837 ) | ( ~n8741 & n8837 ) ;
  assign n8839 = ( x81 & ~n8699 ) | ( x81 & n8838 ) | ( ~n8699 & n8838 ) ;
  assign n8840 = ( x82 & ~n8738 ) | ( x82 & n8839 ) | ( ~n8738 & n8839 ) ;
  assign n8841 = ( x83 & ~n8735 ) | ( x83 & n8840 ) | ( ~n8735 & n8840 ) ;
  assign n8842 = ( x84 & ~n8732 ) | ( x84 & n8841 ) | ( ~n8732 & n8841 ) ;
  assign n8843 = ( x85 & ~n8729 ) | ( x85 & n8842 ) | ( ~n8729 & n8842 ) ;
  assign n8844 = ( x86 & ~n8726 ) | ( x86 & n8843 ) | ( ~n8726 & n8843 ) ;
  assign n8845 = n8832 ^ n8671 ^ x76 ;
  assign n8846 = n8828 ^ n8756 ^ x72 ;
  assign n8847 = ( x87 & ~n8703 ) | ( x87 & n8844 ) | ( ~n8703 & n8844 ) ;
  assign n8848 = ( x88 & ~n8723 ) | ( x88 & n8847 ) | ( ~n8723 & n8847 ) ;
  assign n8849 = ( x89 & ~n8720 ) | ( x89 & n8848 ) | ( ~n8720 & n8848 ) ;
  assign n8850 = ( x90 & ~n8717 ) | ( x90 & n8849 ) | ( ~n8717 & n8849 ) ;
  assign n8851 = ( x91 & ~n8816 ) | ( x91 & n8850 ) | ( ~n8816 & n8850 ) ;
  assign n8852 = ( x92 & ~n8813 ) | ( x92 & n8851 ) | ( ~n8813 & n8851 ) ;
  assign n8853 = ( x93 & ~n8692 ) | ( x93 & n8852 ) | ( ~n8692 & n8852 ) ;
  assign n8854 = ( x94 & ~n8810 ) | ( x94 & n8853 ) | ( ~n8810 & n8853 ) ;
  assign n8855 = n8840 ^ n8735 ^ x83 ;
  assign n8856 = ( x95 & ~n8807 ) | ( x95 & n8854 ) | ( ~n8807 & n8854 ) ;
  assign n8857 = n8842 ^ n8729 ^ x85 ;
  assign n8858 = ( x96 & ~n8665 ) | ( x96 & n8856 ) | ( ~n8665 & n8856 ) ;
  assign n8859 = ( x97 & ~n8804 ) | ( x97 & n8858 ) | ( ~n8804 & n8858 ) ;
  assign n8860 = ( x98 & ~n8801 ) | ( x98 & n8859 ) | ( ~n8801 & n8859 ) ;
  assign n8861 = n8848 ^ n8720 ^ x89 ;
  assign n8862 = n8849 ^ n8717 ^ x90 ;
  assign n8863 = n8837 ^ n8741 ^ x80 ;
  assign n8864 = ( x99 & ~n8697 ) | ( x99 & n8860 ) | ( ~n8697 & n8860 ) ;
  assign n8865 = ( x100 & ~n8798 ) | ( x100 & n8864 ) | ( ~n8798 & n8864 ) ;
  assign n8866 = ( x101 & ~n8795 ) | ( x101 & n8865 ) | ( ~n8795 & n8865 ) ;
  assign n8867 = ( x102 & ~n8792 ) | ( x102 & n8866 ) | ( ~n8792 & n8866 ) ;
  assign n8868 = n8859 ^ n8801 ^ x98 ;
  assign n8869 = n8858 ^ n8804 ^ x97 ;
  assign n8870 = n8856 ^ n8665 ^ x96 ;
  assign n8871 = n8867 ^ n8789 ^ x103 ;
  assign n8872 = ( x103 & ~n8789 ) | ( x103 & n8867 ) | ( ~n8789 & n8867 ) ;
  assign n8873 = n8864 ^ n8798 ^ x100 ;
  assign n8874 = n8854 ^ n8807 ^ x95 ;
  assign n8875 = n8866 ^ n8792 ^ x102 ;
  assign n8876 = n8823 ^ n8698 ^ x67 ;
  assign n8877 = ( x104 & ~n8786 ) | ( x104 & n8872 ) | ( ~n8786 & n8872 ) ;
  assign n8878 = ( x105 & ~n8783 ) | ( x105 & n8877 ) | ( ~n8783 & n8877 ) ;
  assign n8879 = ( x106 & ~n8780 ) | ( x106 & n8878 ) | ( ~n8780 & n8878 ) ;
  assign n8880 = ( x107 & ~n8681 ) | ( x107 & n8879 ) | ( ~n8681 & n8879 ) ;
  assign n8881 = ( x108 & ~n8677 ) | ( x108 & n8880 ) | ( ~n8677 & n8880 ) ;
  assign n8882 = ( x109 & ~n8777 ) | ( x109 & n8881 ) | ( ~n8777 & n8881 ) ;
  assign n8883 = ( x110 & ~n8774 ) | ( x110 & n8882 ) | ( ~n8774 & n8882 ) ;
  assign n8884 = ( x111 & ~n8771 ) | ( x111 & n8883 ) | ( ~n8771 & n8883 ) ;
  assign n8885 = ( x112 & ~n8687 ) | ( x112 & n8884 ) | ( ~n8687 & n8884 ) ;
  assign n8886 = ( x113 & ~n8768 ) | ( x113 & n8885 ) | ( ~n8768 & n8885 ) ;
  assign n8887 = ( x124 & n153 ) | ( x124 & ~n8700 ) | ( n153 & ~n8700 ) ;
  assign n8888 = ( x114 & ~n8704 ) | ( x114 & n8886 ) | ( ~n8704 & n8886 ) ;
  assign n8889 = ( x115 & ~n8702 ) | ( x115 & n8888 ) | ( ~n8702 & n8888 ) ;
  assign n8890 = ( x116 & ~n8668 ) | ( x116 & n8889 ) | ( ~n8668 & n8889 ) ;
  assign n8891 = ( x117 & ~n8714 ) | ( x117 & n8890 ) | ( ~n8714 & n8890 ) ;
  assign n8892 = ( x118 & ~n8658 ) | ( x118 & n8891 ) | ( ~n8658 & n8891 ) ;
  assign n8893 = ( x119 & ~n8688 ) | ( x119 & n8892 ) | ( ~n8688 & n8892 ) ;
  assign n8894 = ( x120 & ~n8705 ) | ( x120 & n8893 ) | ( ~n8705 & n8893 ) ;
  assign n8895 = ( x121 & ~n8696 ) | ( x121 & n8894 ) | ( ~n8696 & n8894 ) ;
  assign n8896 = ( x122 & ~n8711 ) | ( x122 & n8895 ) | ( ~n8711 & n8895 ) ;
  assign n8897 = ( x123 & ~n8708 ) | ( x123 & n8896 ) | ( ~n8708 & n8896 ) ;
  assign n8898 = ( ~x124 & n8700 ) | ( ~x124 & n8897 ) | ( n8700 & n8897 ) ;
  assign n8899 = n8887 | n8898 ;
  assign n8900 = ( ~n8700 & n8833 ) | ( ~n8700 & n8899 ) | ( n8833 & n8899 ) ;
  assign n8901 = n8833 & ~n8899 ;
  assign n8902 = n8897 ^ n8700 ^ x124 ;
  assign n8903 = n8900 ^ n8756 ^ 1'b0 ;
  assign n8904 = ( n8756 & n8846 ) | ( n8756 & ~n8903 ) | ( n8846 & ~n8903 ) ;
  assign n8905 = n8900 ^ n8804 ^ 1'b0 ;
  assign n8906 = ( n8804 & n8869 ) | ( n8804 & ~n8905 ) | ( n8869 & ~n8905 ) ;
  assign n8907 = n8900 ^ n8789 ^ 1'b0 ;
  assign n8908 = n8900 ^ n8687 ^ 1'b0 ;
  assign n8909 = ( n8789 & n8871 ) | ( n8789 & ~n8907 ) | ( n8871 & ~n8907 ) ;
  assign n8910 = n8900 ^ n8698 ^ 1'b0 ;
  assign n8911 = n8900 ^ n8807 ^ 1'b0 ;
  assign n8912 = n8900 ^ n8820 ^ 1'b0 ;
  assign n8913 = ( n8819 & n8820 ) | ( n8819 & n8912 ) | ( n8820 & n8912 ) ;
  assign n8914 = n8900 ^ n8735 ^ 1'b0 ;
  assign n8915 = ( n8735 & n8855 ) | ( n8735 & ~n8914 ) | ( n8855 & ~n8914 ) ;
  assign n8916 = n8900 ^ n8786 ^ 1'b0 ;
  assign n8917 = n8900 ^ n8720 ^ 1'b0 ;
  assign n8918 = n8886 ^ n8704 ^ x114 ;
  assign n8919 = n8879 ^ n8681 ^ x107 ;
  assign n8920 = ( n8807 & n8874 ) | ( n8807 & ~n8911 ) | ( n8874 & ~n8911 ) ;
  assign n8921 = n8900 ^ n8681 ^ 1'b0 ;
  assign n8922 = n8900 ^ n8671 ^ 1'b0 ;
  assign n8923 = n8900 ^ n8665 ^ 1'b0 ;
  assign n8924 = ( n8671 & n8845 ) | ( n8671 & ~n8922 ) | ( n8845 & ~n8922 ) ;
  assign n8925 = n8900 ^ n8801 ^ 1'b0 ;
  assign n8926 = ~n8900 & n8902 ;
  assign n8927 = n8900 ^ n8729 ^ 1'b0 ;
  assign n8928 = n8872 ^ n8786 ^ x104 ;
  assign n8929 = ( n8698 & n8876 ) | ( n8698 & ~n8910 ) | ( n8876 & ~n8910 ) ;
  assign n8930 = ( n8833 & ~n8901 ) | ( n8833 & n8926 ) | ( ~n8901 & n8926 ) ;
  assign n8931 = n8900 ^ n8792 ^ 1'b0 ;
  assign n8932 = n8900 ^ n8704 ^ 1'b0 ;
  assign n8933 = n8900 ^ n8741 ^ 1'b0 ;
  assign n8934 = ( n8786 & ~n8916 ) | ( n8786 & n8928 ) | ( ~n8916 & n8928 ) ;
  assign n8935 = ( n8741 & n8863 ) | ( n8741 & ~n8933 ) | ( n8863 & ~n8933 ) ;
  assign n8936 = n8900 ^ n8717 ^ 1'b0 ;
  assign n8937 = ( n8729 & n8857 ) | ( n8729 & ~n8927 ) | ( n8857 & ~n8927 ) ;
  assign n8938 = ( n8717 & n8862 ) | ( n8717 & ~n8936 ) | ( n8862 & ~n8936 ) ;
  assign n8939 = n8900 ^ n8798 ^ 1'b0 ;
  assign n8940 = n8884 ^ n8687 ^ x112 ;
  assign n8941 = ( n8798 & n8873 ) | ( n8798 & ~n8939 ) | ( n8873 & ~n8939 ) ;
  assign n8942 = ( n8704 & n8918 ) | ( n8704 & ~n8932 ) | ( n8918 & ~n8932 ) ;
  assign n8943 = ( n8792 & n8875 ) | ( n8792 & ~n8931 ) | ( n8875 & ~n8931 ) ;
  assign n8944 = ( n8720 & n8861 ) | ( n8720 & ~n8917 ) | ( n8861 & ~n8917 ) ;
  assign n8945 = ( n8801 & n8868 ) | ( n8801 & ~n8925 ) | ( n8868 & ~n8925 ) ;
  assign n8946 = ( n8681 & n8919 ) | ( n8681 & ~n8921 ) | ( n8919 & ~n8921 ) ;
  assign n8947 = ( n8687 & ~n8908 ) | ( n8687 & n8940 ) | ( ~n8908 & n8940 ) ;
  assign n8948 = ( n8665 & n8870 ) | ( n8665 & ~n8923 ) | ( n8870 & ~n8923 ) ;
  assign n8949 = n8896 ^ n8708 ^ x123 ;
  assign n8950 = n8900 ^ n8708 ^ 1'b0 ;
  assign n8951 = ( n8708 & n8949 ) | ( n8708 & ~n8950 ) | ( n8949 & ~n8950 ) ;
  assign n8952 = n8895 ^ n8711 ^ x122 ;
  assign n8953 = n8900 ^ n8711 ^ 1'b0 ;
  assign n8954 = ( n8711 & n8952 ) | ( n8711 & ~n8953 ) | ( n8952 & ~n8953 ) ;
  assign n8955 = n8894 ^ n8696 ^ x121 ;
  assign n8956 = n8900 ^ n8696 ^ 1'b0 ;
  assign n8957 = ( n8696 & n8955 ) | ( n8696 & ~n8956 ) | ( n8955 & ~n8956 ) ;
  assign n8958 = n8850 ^ n8816 ^ x91 ;
  assign n8959 = n8900 ^ n8816 ^ 1'b0 ;
  assign n8960 = ( n8816 & n8958 ) | ( n8816 & ~n8959 ) | ( n8958 & ~n8959 ) ;
  assign n8961 = n8847 ^ n8723 ^ x88 ;
  assign n8962 = n8900 ^ n8723 ^ 1'b0 ;
  assign n8963 = ( n8723 & n8961 ) | ( n8723 & ~n8962 ) | ( n8961 & ~n8962 ) ;
  assign n8964 = n8844 ^ n8703 ^ x87 ;
  assign n8965 = n8900 ^ n8703 ^ 1'b0 ;
  assign n8966 = ( n8703 & n8964 ) | ( n8703 & ~n8965 ) | ( n8964 & ~n8965 ) ;
  assign n8967 = n8843 ^ n8726 ^ x86 ;
  assign n8968 = n8900 ^ n8726 ^ 1'b0 ;
  assign n8969 = ( n8726 & n8967 ) | ( n8726 & ~n8968 ) | ( n8967 & ~n8968 ) ;
  assign n8970 = n8841 ^ n8732 ^ x84 ;
  assign n8971 = n8900 ^ n8732 ^ 1'b0 ;
  assign n8972 = ( n8732 & n8970 ) | ( n8732 & ~n8971 ) | ( n8970 & ~n8971 ) ;
  assign n8973 = n8839 ^ n8738 ^ x82 ;
  assign n8974 = n8900 ^ n8738 ^ 1'b0 ;
  assign n8975 = ( n8738 & n8973 ) | ( n8738 & ~n8974 ) | ( n8973 & ~n8974 ) ;
  assign n8976 = n8838 ^ n8699 ^ x81 ;
  assign n8977 = n8900 ^ n8699 ^ 1'b0 ;
  assign n8978 = ( n8699 & n8976 ) | ( n8699 & ~n8977 ) | ( n8976 & ~n8977 ) ;
  assign n8979 = n8836 ^ n8694 ^ x79 ;
  assign n8980 = n8900 ^ n8694 ^ 1'b0 ;
  assign n8981 = ( n8694 & n8979 ) | ( n8694 & ~n8980 ) | ( n8979 & ~n8980 ) ;
  assign n8982 = n8835 ^ n8675 ^ x78 ;
  assign n8983 = n8900 ^ n8675 ^ 1'b0 ;
  assign n8984 = ( n8675 & n8982 ) | ( n8675 & ~n8983 ) | ( n8982 & ~n8983 ) ;
  assign n8985 = n8834 ^ n8744 ^ x77 ;
  assign n8986 = n8900 ^ n8744 ^ 1'b0 ;
  assign n8987 = ( n8744 & n8985 ) | ( n8744 & ~n8986 ) | ( n8985 & ~n8986 ) ;
  assign n8988 = n8831 ^ n8747 ^ x75 ;
  assign n8989 = n8900 ^ n8747 ^ 1'b0 ;
  assign n8990 = ( n8747 & n8988 ) | ( n8747 & ~n8989 ) | ( n8988 & ~n8989 ) ;
  assign n8991 = n8830 ^ n8750 ^ x74 ;
  assign n8992 = n8900 ^ n8750 ^ 1'b0 ;
  assign n8993 = ( n8750 & n8991 ) | ( n8750 & ~n8992 ) | ( n8991 & ~n8992 ) ;
  assign n8994 = n8829 ^ n8753 ^ x73 ;
  assign n8995 = n8900 ^ n8753 ^ 1'b0 ;
  assign n8996 = ( n8753 & n8994 ) | ( n8753 & ~n8995 ) | ( n8994 & ~n8995 ) ;
  assign n8997 = n8827 ^ n8759 ^ x71 ;
  assign n8998 = n8900 ^ n8759 ^ 1'b0 ;
  assign n8999 = ( n8759 & n8997 ) | ( n8759 & ~n8998 ) | ( n8997 & ~n8998 ) ;
  assign n9000 = n8826 ^ n8762 ^ x70 ;
  assign n9001 = n8900 ^ n8762 ^ 1'b0 ;
  assign n9002 = ( n8762 & n9000 ) | ( n8762 & ~n9001 ) | ( n9000 & ~n9001 ) ;
  assign n9003 = n8825 ^ n8765 ^ x69 ;
  assign n9004 = n8900 ^ n8765 ^ 1'b0 ;
  assign n9005 = ( n8765 & n9003 ) | ( n8765 & ~n9004 ) | ( n9003 & ~n9004 ) ;
  assign n9006 = n8824 ^ n8683 ^ x68 ;
  assign n9007 = n8900 ^ n8683 ^ 1'b0 ;
  assign n9008 = ( n8683 & n9006 ) | ( n8683 & ~n9007 ) | ( n9006 & ~n9007 ) ;
  assign n9009 = n8893 ^ n8705 ^ x120 ;
  assign n9010 = n8900 ^ n8705 ^ 1'b0 ;
  assign n9011 = ( n8705 & n9009 ) | ( n8705 & ~n9010 ) | ( n9009 & ~n9010 ) ;
  assign n9012 = n8892 ^ n8688 ^ x119 ;
  assign n9013 = n8900 ^ n8688 ^ 1'b0 ;
  assign n9014 = ( n8688 & n9012 ) | ( n8688 & ~n9013 ) | ( n9012 & ~n9013 ) ;
  assign n9015 = n8891 ^ n8658 ^ x118 ;
  assign n9016 = n8900 ^ n8658 ^ 1'b0 ;
  assign n9017 = ( n8658 & n9015 ) | ( n8658 & ~n9016 ) | ( n9015 & ~n9016 ) ;
  assign n9018 = n8890 ^ n8714 ^ x117 ;
  assign n9019 = n8900 ^ n8714 ^ 1'b0 ;
  assign n9020 = ( n8714 & n9018 ) | ( n8714 & ~n9019 ) | ( n9018 & ~n9019 ) ;
  assign n9021 = n8889 ^ n8668 ^ x116 ;
  assign n9022 = n8900 ^ n8668 ^ 1'b0 ;
  assign n9023 = ( n8668 & n9021 ) | ( n8668 & ~n9022 ) | ( n9021 & ~n9022 ) ;
  assign n9024 = n8888 ^ n8702 ^ x115 ;
  assign n9025 = n8900 ^ n8702 ^ 1'b0 ;
  assign n9026 = ( n8702 & n9024 ) | ( n8702 & ~n9025 ) | ( n9024 & ~n9025 ) ;
  assign n9027 = n8885 ^ n8768 ^ x113 ;
  assign n9028 = n8900 ^ n8768 ^ 1'b0 ;
  assign n9029 = ( n8768 & n9027 ) | ( n8768 & ~n9028 ) | ( n9027 & ~n9028 ) ;
  assign n9030 = n8883 ^ n8771 ^ x111 ;
  assign n9031 = n8900 ^ n8771 ^ 1'b0 ;
  assign n9032 = ( n8771 & n9030 ) | ( n8771 & ~n9031 ) | ( n9030 & ~n9031 ) ;
  assign n9033 = n8881 ^ n8777 ^ x109 ;
  assign n9034 = n8900 ^ n8777 ^ 1'b0 ;
  assign n9035 = ( n8777 & n9033 ) | ( n8777 & ~n9034 ) | ( n9033 & ~n9034 ) ;
  assign n9036 = n8880 ^ n8677 ^ x108 ;
  assign n9037 = n8900 ^ n8677 ^ 1'b0 ;
  assign n9038 = ( n8677 & n9036 ) | ( n8677 & ~n9037 ) | ( n9036 & ~n9037 ) ;
  assign n9039 = n8878 ^ n8780 ^ x106 ;
  assign n9040 = n8900 ^ n8780 ^ 1'b0 ;
  assign n9041 = ( n8780 & n9039 ) | ( n8780 & ~n9040 ) | ( n9039 & ~n9040 ) ;
  assign n9042 = n8877 ^ n8783 ^ x105 ;
  assign n9043 = n8900 ^ n8783 ^ 1'b0 ;
  assign n9044 = ( n8783 & n9042 ) | ( n8783 & ~n9043 ) | ( n9042 & ~n9043 ) ;
  assign n9045 = n8865 ^ n8795 ^ x101 ;
  assign n9046 = n8900 ^ n8795 ^ 1'b0 ;
  assign n9047 = ( n8795 & n9045 ) | ( n8795 & ~n9046 ) | ( n9045 & ~n9046 ) ;
  assign n9048 = n8860 ^ n8697 ^ x99 ;
  assign n9049 = n8900 ^ n8697 ^ 1'b0 ;
  assign n9050 = ( n8697 & n9048 ) | ( n8697 & ~n9049 ) | ( n9048 & ~n9049 ) ;
  assign n9051 = n8853 ^ n8810 ^ x94 ;
  assign n9052 = n8900 ^ n8810 ^ 1'b0 ;
  assign n9053 = ( n8810 & n9051 ) | ( n8810 & ~n9052 ) | ( n9051 & ~n9052 ) ;
  assign n9054 = n8852 ^ n8692 ^ x93 ;
  assign n9055 = n8900 ^ n8692 ^ 1'b0 ;
  assign n9056 = ( n8692 & n9054 ) | ( n8692 & ~n9055 ) | ( n9054 & ~n9055 ) ;
  assign n9057 = n8851 ^ n8813 ^ x92 ;
  assign n9058 = n8900 ^ n8813 ^ 1'b0 ;
  assign n9059 = ( n8813 & n9057 ) | ( n8813 & ~n9058 ) | ( n9057 & ~n9058 ) ;
  assign n9060 = n8882 ^ n8774 ^ x110 ;
  assign n9061 = n8900 ^ n8774 ^ 1'b0 ;
  assign n9062 = n8900 ^ n8822 ^ 1'b0 ;
  assign n9063 = ( n8701 & n8822 ) | ( n8701 & n9062 ) | ( n8822 & n9062 ) ;
  assign n9064 = ~x2 & x64 ;
  assign n9065 = x64 & n8900 ;
  assign n9066 = n9065 ^ x64 ^ x3 ;
  assign n9067 = n9066 ^ n9064 ^ x65 ;
  assign n9068 = ( x65 & n9064 ) | ( x65 & n9067 ) | ( n9064 & n9067 ) ;
  assign n9069 = n9068 ^ n8913 ^ x66 ;
  assign n9070 = ( x66 & n9068 ) | ( x66 & n9069 ) | ( n9068 & n9069 ) ;
  assign n9071 = ( x67 & ~n9063 ) | ( x67 & n9070 ) | ( ~n9063 & n9070 ) ;
  assign n9072 = ( x68 & ~n8929 ) | ( x68 & n9071 ) | ( ~n8929 & n9071 ) ;
  assign n9073 = ( x69 & ~n9008 ) | ( x69 & n9072 ) | ( ~n9008 & n9072 ) ;
  assign n9074 = ( x70 & ~n9005 ) | ( x70 & n9073 ) | ( ~n9005 & n9073 ) ;
  assign n9075 = ( x71 & ~n9002 ) | ( x71 & n9074 ) | ( ~n9002 & n9074 ) ;
  assign n9076 = ( x72 & ~n8999 ) | ( x72 & n9075 ) | ( ~n8999 & n9075 ) ;
  assign n9077 = ( x73 & ~n8904 ) | ( x73 & n9076 ) | ( ~n8904 & n9076 ) ;
  assign n9078 = ( x74 & ~n8996 ) | ( x74 & n9077 ) | ( ~n8996 & n9077 ) ;
  assign n9079 = ( x75 & ~n8993 ) | ( x75 & n9078 ) | ( ~n8993 & n9078 ) ;
  assign n9080 = ( x76 & ~n8990 ) | ( x76 & n9079 ) | ( ~n8990 & n9079 ) ;
  assign n9081 = ( x77 & ~n8924 ) | ( x77 & n9080 ) | ( ~n8924 & n9080 ) ;
  assign n9082 = ( x78 & ~n8987 ) | ( x78 & n9081 ) | ( ~n8987 & n9081 ) ;
  assign n9083 = ( x79 & ~n8984 ) | ( x79 & n9082 ) | ( ~n8984 & n9082 ) ;
  assign n9084 = ( x80 & ~n8981 ) | ( x80 & n9083 ) | ( ~n8981 & n9083 ) ;
  assign n9085 = ( x81 & ~n8935 ) | ( x81 & n9084 ) | ( ~n8935 & n9084 ) ;
  assign n9086 = ( x82 & ~n8978 ) | ( x82 & n9085 ) | ( ~n8978 & n9085 ) ;
  assign n9087 = ( x83 & ~n8975 ) | ( x83 & n9086 ) | ( ~n8975 & n9086 ) ;
  assign n9088 = ( x84 & ~n8915 ) | ( x84 & n9087 ) | ( ~n8915 & n9087 ) ;
  assign n9089 = ( x85 & ~n8972 ) | ( x85 & n9088 ) | ( ~n8972 & n9088 ) ;
  assign n9090 = ( x86 & ~n8937 ) | ( x86 & n9089 ) | ( ~n8937 & n9089 ) ;
  assign n9091 = ( x87 & ~n8969 ) | ( x87 & n9090 ) | ( ~n8969 & n9090 ) ;
  assign n9092 = ( x88 & ~n8966 ) | ( x88 & n9091 ) | ( ~n8966 & n9091 ) ;
  assign n9093 = ( x89 & ~n8963 ) | ( x89 & n9092 ) | ( ~n8963 & n9092 ) ;
  assign n9094 = ( x90 & ~n8944 ) | ( x90 & n9093 ) | ( ~n8944 & n9093 ) ;
  assign n9095 = ( x91 & ~n8938 ) | ( x91 & n9094 ) | ( ~n8938 & n9094 ) ;
  assign n9096 = ( x92 & ~n8960 ) | ( x92 & n9095 ) | ( ~n8960 & n9095 ) ;
  assign n9097 = ( x93 & ~n9059 ) | ( x93 & n9096 ) | ( ~n9059 & n9096 ) ;
  assign n9098 = ( x94 & ~n9056 ) | ( x94 & n9097 ) | ( ~n9056 & n9097 ) ;
  assign n9099 = ( x95 & ~n9053 ) | ( x95 & n9098 ) | ( ~n9053 & n9098 ) ;
  assign n9100 = ( x96 & ~n8920 ) | ( x96 & n9099 ) | ( ~n8920 & n9099 ) ;
  assign n9101 = ( x97 & ~n8948 ) | ( x97 & n9100 ) | ( ~n8948 & n9100 ) ;
  assign n9102 = ( x98 & ~n8906 ) | ( x98 & n9101 ) | ( ~n8906 & n9101 ) ;
  assign n9103 = n9077 ^ n8996 ^ x74 ;
  assign n9104 = n9071 ^ n8929 ^ x68 ;
  assign n9105 = n9070 ^ n9063 ^ x67 ;
  assign n9106 = ( n8774 & n9060 ) | ( n8774 & ~n9061 ) | ( n9060 & ~n9061 ) ;
  assign n9107 = ( x99 & ~n8945 ) | ( x99 & n9102 ) | ( ~n8945 & n9102 ) ;
  assign n9108 = ( x100 & ~n9050 ) | ( x100 & n9107 ) | ( ~n9050 & n9107 ) ;
  assign n9109 = ( x101 & ~n8941 ) | ( x101 & n9108 ) | ( ~n8941 & n9108 ) ;
  assign n9110 = ( x102 & ~n9047 ) | ( x102 & n9109 ) | ( ~n9047 & n9109 ) ;
  assign n9111 = ( x103 & ~n8943 ) | ( x103 & n9110 ) | ( ~n8943 & n9110 ) ;
  assign n9112 = ( x104 & ~n8909 ) | ( x104 & n9111 ) | ( ~n8909 & n9111 ) ;
  assign n9113 = ( x105 & ~n8934 ) | ( x105 & n9112 ) | ( ~n8934 & n9112 ) ;
  assign n9114 = ( x106 & ~n9044 ) | ( x106 & n9113 ) | ( ~n9044 & n9113 ) ;
  assign n9115 = ( x107 & ~n9041 ) | ( x107 & n9114 ) | ( ~n9041 & n9114 ) ;
  assign n9116 = ( x108 & ~n8946 ) | ( x108 & n9115 ) | ( ~n8946 & n9115 ) ;
  assign n9117 = ( x109 & ~n9038 ) | ( x109 & n9116 ) | ( ~n9038 & n9116 ) ;
  assign n9118 = ( x110 & ~n9035 ) | ( x110 & n9117 ) | ( ~n9035 & n9117 ) ;
  assign n9119 = ( x111 & ~n9106 ) | ( x111 & n9118 ) | ( ~n9106 & n9118 ) ;
  assign n9120 = ( x112 & ~n9032 ) | ( x112 & n9119 ) | ( ~n9032 & n9119 ) ;
  assign n9121 = ( x113 & ~n8947 ) | ( x113 & n9120 ) | ( ~n8947 & n9120 ) ;
  assign n9122 = ( x114 & ~n9029 ) | ( x114 & n9121 ) | ( ~n9029 & n9121 ) ;
  assign n9123 = ( x115 & ~n8942 ) | ( x115 & n9122 ) | ( ~n8942 & n9122 ) ;
  assign n9124 = ( x116 & ~n9026 ) | ( x116 & n9123 ) | ( ~n9026 & n9123 ) ;
  assign n9125 = ( x117 & ~n9023 ) | ( x117 & n9124 ) | ( ~n9023 & n9124 ) ;
  assign n9126 = ( x118 & ~n9020 ) | ( x118 & n9125 ) | ( ~n9020 & n9125 ) ;
  assign n9127 = ( x119 & ~n9017 ) | ( x119 & n9126 ) | ( ~n9017 & n9126 ) ;
  assign n9128 = ( x120 & ~n9014 ) | ( x120 & n9127 ) | ( ~n9014 & n9127 ) ;
  assign n9129 = ( x121 & ~n9011 ) | ( x121 & n9128 ) | ( ~n9011 & n9128 ) ;
  assign n9130 = ( x122 & ~n8957 ) | ( x122 & n9129 ) | ( ~n8957 & n9129 ) ;
  assign n9131 = ( x123 & ~n8954 ) | ( x123 & n9130 ) | ( ~n8954 & n9130 ) ;
  assign n9132 = n9131 ^ n8951 ^ x124 ;
  assign n9133 = ( x124 & ~n8951 ) | ( x124 & n9131 ) | ( ~n8951 & n9131 ) ;
  assign n9134 = ( x125 & ~n8930 ) | ( x125 & n9133 ) | ( ~n8930 & n9133 ) ;
  assign n9135 = n147 | n9134 ;
  assign n9136 = n9135 ^ n8951 ^ 1'b0 ;
  assign n9137 = ( n8951 & n9132 ) | ( n8951 & ~n9136 ) | ( n9132 & ~n9136 ) ;
  assign n9138 = n9130 ^ n8954 ^ x123 ;
  assign n9139 = n9135 ^ n8954 ^ 1'b0 ;
  assign n9140 = ( n8954 & n9138 ) | ( n8954 & ~n9139 ) | ( n9138 & ~n9139 ) ;
  assign n9141 = n9129 ^ n8957 ^ x122 ;
  assign n9142 = n9135 ^ n8957 ^ 1'b0 ;
  assign n9143 = ( n8957 & n9141 ) | ( n8957 & ~n9142 ) | ( n9141 & ~n9142 ) ;
  assign n9144 = n9128 ^ n9011 ^ x121 ;
  assign n9145 = n9135 ^ n9011 ^ 1'b0 ;
  assign n9146 = ( n9011 & n9144 ) | ( n9011 & ~n9145 ) | ( n9144 & ~n9145 ) ;
  assign n9147 = n9127 ^ n9014 ^ x120 ;
  assign n9148 = n9135 ^ n9014 ^ 1'b0 ;
  assign n9149 = ( n9014 & n9147 ) | ( n9014 & ~n9148 ) | ( n9147 & ~n9148 ) ;
  assign n9150 = n9126 ^ n9017 ^ x119 ;
  assign n9151 = n9135 ^ n9017 ^ 1'b0 ;
  assign n9152 = ( n9017 & n9150 ) | ( n9017 & ~n9151 ) | ( n9150 & ~n9151 ) ;
  assign n9153 = n9125 ^ n9020 ^ x118 ;
  assign n9154 = n9135 ^ n9020 ^ 1'b0 ;
  assign n9155 = ( n9020 & n9153 ) | ( n9020 & ~n9154 ) | ( n9153 & ~n9154 ) ;
  assign n9156 = n9124 ^ n9023 ^ x117 ;
  assign n9157 = n9135 ^ n9023 ^ 1'b0 ;
  assign n9158 = ( n9023 & n9156 ) | ( n9023 & ~n9157 ) | ( n9156 & ~n9157 ) ;
  assign n9159 = n9123 ^ n9026 ^ x116 ;
  assign n9160 = n9135 ^ n9026 ^ 1'b0 ;
  assign n9161 = ( n9026 & n9159 ) | ( n9026 & ~n9160 ) | ( n9159 & ~n9160 ) ;
  assign n9162 = n9122 ^ n8942 ^ x115 ;
  assign n9163 = n9135 ^ n8942 ^ 1'b0 ;
  assign n9164 = ( n8942 & n9162 ) | ( n8942 & ~n9163 ) | ( n9162 & ~n9163 ) ;
  assign n9165 = n9135 ^ n8996 ^ 1'b0 ;
  assign n9166 = ( n8996 & n9103 ) | ( n8996 & ~n9165 ) | ( n9103 & ~n9165 ) ;
  assign n9167 = n9135 ^ n8929 ^ 1'b0 ;
  assign n9168 = ( n8929 & n9104 ) | ( n8929 & ~n9167 ) | ( n9104 & ~n9167 ) ;
  assign n9169 = n9135 ^ n9063 ^ 1'b0 ;
  assign n9170 = ( n9063 & n9105 ) | ( n9063 & ~n9169 ) | ( n9105 & ~n9169 ) ;
  assign n9171 = n9108 ^ n8941 ^ x101 ;
  assign n9172 = n153 | n9133 ;
  assign n9173 = n9111 ^ n8909 ^ x104 ;
  assign n9174 = ( n8930 & n9135 ) | ( n8930 & ~n9172 ) | ( n9135 & ~n9172 ) ;
  assign n9175 = n9135 ^ n8909 ^ 1'b0 ;
  assign n9176 = ( n8909 & n9173 ) | ( n8909 & ~n9175 ) | ( n9173 & ~n9175 ) ;
  assign n9177 = n9109 ^ n9047 ^ x102 ;
  assign n9178 = n9121 ^ n9029 ^ x114 ;
  assign n9179 = n9135 ^ n8941 ^ 1'b0 ;
  assign n9180 = n9135 ^ n9067 ^ 1'b0 ;
  assign n9181 = n9116 ^ n9038 ^ x109 ;
  assign n9182 = ( n8941 & n9171 ) | ( n8941 & ~n9179 ) | ( n9171 & ~n9179 ) ;
  assign n9183 = n9115 ^ n8946 ^ x108 ;
  assign n9184 = n9113 ^ n9044 ^ x106 ;
  assign n9185 = n9135 ^ n8934 ^ 1'b0 ;
  assign n9186 = n9072 ^ n9008 ^ x69 ;
  assign n9187 = n9120 ^ n8947 ^ x113 ;
  assign n9188 = n9135 ^ n9035 ^ 1'b0 ;
  assign n9189 = n9110 ^ n8943 ^ x103 ;
  assign n9190 = ( n9066 & n9067 ) | ( n9066 & n9180 ) | ( n9067 & n9180 ) ;
  assign n9191 = n9135 ^ n9029 ^ 1'b0 ;
  assign n9192 = n9119 ^ n9032 ^ x112 ;
  assign n9193 = n9135 ^ n9032 ^ 1'b0 ;
  assign n9194 = ( n9032 & n9192 ) | ( n9032 & ~n9193 ) | ( n9192 & ~n9193 ) ;
  assign n9195 = n9135 ^ n9106 ^ 1'b0 ;
  assign n9196 = n9118 ^ n9106 ^ x111 ;
  assign n9197 = n9135 ^ n9041 ^ 1'b0 ;
  assign n9198 = ( n9106 & ~n9195 ) | ( n9106 & n9196 ) | ( ~n9195 & n9196 ) ;
  assign n9199 = n9135 ^ n8946 ^ 1'b0 ;
  assign n9200 = n9135 ^ n9047 ^ 1'b0 ;
  assign n9201 = n9112 ^ n8934 ^ x105 ;
  assign n9202 = ( n9047 & n9177 ) | ( n9047 & ~n9200 ) | ( n9177 & ~n9200 ) ;
  assign n9203 = n9114 ^ n9041 ^ x107 ;
  assign n9204 = ( n9029 & n9178 ) | ( n9029 & ~n9191 ) | ( n9178 & ~n9191 ) ;
  assign n9205 = n9135 ^ n8943 ^ 1'b0 ;
  assign n9206 = ( n9041 & ~n9197 ) | ( n9041 & n9203 ) | ( ~n9197 & n9203 ) ;
  assign n9207 = ( n8943 & n9189 ) | ( n8943 & ~n9205 ) | ( n9189 & ~n9205 ) ;
  assign n9208 = n9135 ^ n9038 ^ 1'b0 ;
  assign n9209 = n9117 ^ n9035 ^ x110 ;
  assign n9210 = n9135 ^ n9044 ^ 1'b0 ;
  assign n9211 = ( n8934 & ~n9185 ) | ( n8934 & n9201 ) | ( ~n9185 & n9201 ) ;
  assign n9212 = n9135 ^ n8947 ^ 1'b0 ;
  assign n9213 = ( n9038 & n9181 ) | ( n9038 & ~n9208 ) | ( n9181 & ~n9208 ) ;
  assign n9214 = ( n8947 & n9187 ) | ( n8947 & ~n9212 ) | ( n9187 & ~n9212 ) ;
  assign n9215 = ( n9044 & n9184 ) | ( n9044 & ~n9210 ) | ( n9184 & ~n9210 ) ;
  assign n9216 = n9135 ^ n9008 ^ 1'b0 ;
  assign n9217 = ( n8946 & n9183 ) | ( n8946 & ~n9199 ) | ( n9183 & ~n9199 ) ;
  assign n9218 = ( n9035 & ~n9188 ) | ( n9035 & n9209 ) | ( ~n9188 & n9209 ) ;
  assign n9219 = ( n9008 & n9186 ) | ( n9008 & ~n9216 ) | ( n9186 & ~n9216 ) ;
  assign n9220 = n9107 ^ n9050 ^ x100 ;
  assign n9221 = n9135 ^ n9050 ^ 1'b0 ;
  assign n9222 = ( n9050 & n9220 ) | ( n9050 & ~n9221 ) | ( n9220 & ~n9221 ) ;
  assign n9223 = n9102 ^ n8945 ^ x99 ;
  assign n9224 = n9135 ^ n8945 ^ 1'b0 ;
  assign n9225 = ( n8945 & n9223 ) | ( n8945 & ~n9224 ) | ( n9223 & ~n9224 ) ;
  assign n9226 = n9101 ^ n8906 ^ x98 ;
  assign n9227 = n9135 ^ n8906 ^ 1'b0 ;
  assign n9228 = ( n8906 & n9226 ) | ( n8906 & ~n9227 ) | ( n9226 & ~n9227 ) ;
  assign n9229 = n9100 ^ n8948 ^ x97 ;
  assign n9230 = n9135 ^ n8948 ^ 1'b0 ;
  assign n9231 = ( n8948 & n9229 ) | ( n8948 & ~n9230 ) | ( n9229 & ~n9230 ) ;
  assign n9232 = n9099 ^ n8920 ^ x96 ;
  assign n9233 = n9135 ^ n8920 ^ 1'b0 ;
  assign n9234 = ( n8920 & n9232 ) | ( n8920 & ~n9233 ) | ( n9232 & ~n9233 ) ;
  assign n9235 = n9098 ^ n9053 ^ x95 ;
  assign n9236 = n9135 ^ n9053 ^ 1'b0 ;
  assign n9237 = ( n9053 & n9235 ) | ( n9053 & ~n9236 ) | ( n9235 & ~n9236 ) ;
  assign n9238 = n9097 ^ n9056 ^ x94 ;
  assign n9239 = n9135 ^ n9056 ^ 1'b0 ;
  assign n9240 = ( n9056 & n9238 ) | ( n9056 & ~n9239 ) | ( n9238 & ~n9239 ) ;
  assign n9241 = n9093 ^ n8944 ^ x90 ;
  assign n9242 = n9135 ^ n8944 ^ 1'b0 ;
  assign n9243 = ( n8944 & n9241 ) | ( n8944 & ~n9242 ) | ( n9241 & ~n9242 ) ;
  assign n9244 = n9086 ^ n8975 ^ x83 ;
  assign n9245 = n9135 ^ n8975 ^ 1'b0 ;
  assign n9246 = ( n8975 & n9244 ) | ( n8975 & ~n9245 ) | ( n9244 & ~n9245 ) ;
  assign n9247 = n9085 ^ n8978 ^ x82 ;
  assign n9248 = n9135 ^ n8978 ^ 1'b0 ;
  assign n9249 = ( n8978 & n9247 ) | ( n8978 & ~n9248 ) | ( n9247 & ~n9248 ) ;
  assign n9250 = n9083 ^ n8981 ^ x80 ;
  assign n9251 = n9135 ^ n8981 ^ 1'b0 ;
  assign n9252 = ( n8981 & n9250 ) | ( n8981 & ~n9251 ) | ( n9250 & ~n9251 ) ;
  assign n9253 = n9082 ^ n8984 ^ x79 ;
  assign n9254 = n9135 ^ n8984 ^ 1'b0 ;
  assign n9255 = ( n8984 & n9253 ) | ( n8984 & ~n9254 ) | ( n9253 & ~n9254 ) ;
  assign n9256 = n9079 ^ n8990 ^ x76 ;
  assign n9257 = n9135 ^ n8990 ^ 1'b0 ;
  assign n9258 = ( n8990 & n9256 ) | ( n8990 & ~n9257 ) | ( n9256 & ~n9257 ) ;
  assign n9259 = n9078 ^ n8993 ^ x75 ;
  assign n9260 = n9135 ^ n8993 ^ 1'b0 ;
  assign n9261 = ( n8993 & n9259 ) | ( n8993 & ~n9260 ) | ( n9259 & ~n9260 ) ;
  assign n9262 = n9096 ^ n9059 ^ x93 ;
  assign n9263 = n9135 ^ n9059 ^ 1'b0 ;
  assign n9264 = ( n9059 & n9262 ) | ( n9059 & ~n9263 ) | ( n9262 & ~n9263 ) ;
  assign n9265 = n9095 ^ n8960 ^ x92 ;
  assign n9266 = n9135 ^ n8960 ^ 1'b0 ;
  assign n9267 = ( n8960 & n9265 ) | ( n8960 & ~n9266 ) | ( n9265 & ~n9266 ) ;
  assign n9268 = n9094 ^ n8938 ^ x91 ;
  assign n9269 = n9135 ^ n8938 ^ 1'b0 ;
  assign n9270 = ( n8938 & n9268 ) | ( n8938 & ~n9269 ) | ( n9268 & ~n9269 ) ;
  assign n9271 = n9092 ^ n8963 ^ x89 ;
  assign n9272 = n9135 ^ n8963 ^ 1'b0 ;
  assign n9273 = ( n8963 & n9271 ) | ( n8963 & ~n9272 ) | ( n9271 & ~n9272 ) ;
  assign n9274 = n9091 ^ n8966 ^ x88 ;
  assign n9275 = n9135 ^ n8966 ^ 1'b0 ;
  assign n9276 = ( n8966 & n9274 ) | ( n8966 & ~n9275 ) | ( n9274 & ~n9275 ) ;
  assign n9277 = n9090 ^ n8969 ^ x87 ;
  assign n9278 = n9135 ^ n8969 ^ 1'b0 ;
  assign n9279 = ( n8969 & n9277 ) | ( n8969 & ~n9278 ) | ( n9277 & ~n9278 ) ;
  assign n9280 = n9089 ^ n8937 ^ x86 ;
  assign n9281 = n9135 ^ n8937 ^ 1'b0 ;
  assign n9282 = ( n8937 & n9280 ) | ( n8937 & ~n9281 ) | ( n9280 & ~n9281 ) ;
  assign n9283 = n9088 ^ n8972 ^ x85 ;
  assign n9284 = n9135 ^ n8972 ^ 1'b0 ;
  assign n9285 = ( n8972 & n9283 ) | ( n8972 & ~n9284 ) | ( n9283 & ~n9284 ) ;
  assign n9286 = n9087 ^ n8915 ^ x84 ;
  assign n9287 = n9135 ^ n8915 ^ 1'b0 ;
  assign n9288 = ( n8915 & n9286 ) | ( n8915 & ~n9287 ) | ( n9286 & ~n9287 ) ;
  assign n9289 = n9135 ^ n8935 ^ 1'b0 ;
  assign n9290 = n9081 ^ n8987 ^ x78 ;
  assign n9291 = n9135 ^ n8987 ^ 1'b0 ;
  assign n9292 = ( n8987 & n9290 ) | ( n8987 & ~n9291 ) | ( n9290 & ~n9291 ) ;
  assign n9293 = n9080 ^ n8924 ^ x77 ;
  assign n9294 = n9135 ^ n8924 ^ 1'b0 ;
  assign n9295 = ( n8924 & n9293 ) | ( n8924 & ~n9294 ) | ( n9293 & ~n9294 ) ;
  assign n9296 = n9076 ^ n8904 ^ x73 ;
  assign n9297 = n9135 ^ n8904 ^ 1'b0 ;
  assign n9298 = ( n8904 & n9296 ) | ( n8904 & ~n9297 ) | ( n9296 & ~n9297 ) ;
  assign n9299 = n9084 ^ n8935 ^ x81 ;
  assign n9300 = ( n8935 & ~n9289 ) | ( n8935 & n9299 ) | ( ~n9289 & n9299 ) ;
  assign n9301 = n9075 ^ n8999 ^ x72 ;
  assign n9302 = n9135 ^ n8999 ^ 1'b0 ;
  assign n9303 = ( n8999 & n9301 ) | ( n8999 & ~n9302 ) | ( n9301 & ~n9302 ) ;
  assign n9304 = n9074 ^ n9002 ^ x71 ;
  assign n9305 = n9135 ^ n9002 ^ 1'b0 ;
  assign n9306 = ( n9002 & n9304 ) | ( n9002 & ~n9305 ) | ( n9304 & ~n9305 ) ;
  assign n9307 = n9073 ^ n9005 ^ x70 ;
  assign n9308 = n9135 ^ n9005 ^ 1'b0 ;
  assign n9309 = ( n9005 & n9307 ) | ( n9005 & ~n9308 ) | ( n9307 & ~n9308 ) ;
  assign n9310 = n9135 ^ n9069 ^ 1'b0 ;
  assign n9311 = ( n8913 & n9069 ) | ( n8913 & n9310 ) | ( n9069 & n9310 ) ;
  assign n9312 = x64 & n9135 ;
  assign n9313 = ~x1 & x64 ;
  assign n9314 = n9312 ^ x64 ^ x2 ;
  assign n9315 = n9314 ^ n9313 ^ x65 ;
  assign n9316 = ( x65 & n9313 ) | ( x65 & n9315 ) | ( n9313 & n9315 ) ;
  assign n9317 = n9316 ^ n9190 ^ x66 ;
  assign n9318 = ( x66 & n9316 ) | ( x66 & n9317 ) | ( n9316 & n9317 ) ;
  assign n9319 = ( x67 & ~n9311 ) | ( x67 & n9318 ) | ( ~n9311 & n9318 ) ;
  assign n9320 = ( x68 & ~n9170 ) | ( x68 & n9319 ) | ( ~n9170 & n9319 ) ;
  assign n9321 = ( x69 & ~n9168 ) | ( x69 & n9320 ) | ( ~n9168 & n9320 ) ;
  assign n9322 = ( x70 & ~n9219 ) | ( x70 & n9321 ) | ( ~n9219 & n9321 ) ;
  assign n9323 = ( x71 & ~n9309 ) | ( x71 & n9322 ) | ( ~n9309 & n9322 ) ;
  assign n9324 = ( x72 & ~n9306 ) | ( x72 & n9323 ) | ( ~n9306 & n9323 ) ;
  assign n9325 = ( x73 & ~n9303 ) | ( x73 & n9324 ) | ( ~n9303 & n9324 ) ;
  assign n9326 = ( x74 & ~n9298 ) | ( x74 & n9325 ) | ( ~n9298 & n9325 ) ;
  assign n9327 = ( x75 & ~n9166 ) | ( x75 & n9326 ) | ( ~n9166 & n9326 ) ;
  assign n9328 = ( x76 & ~n9261 ) | ( x76 & n9327 ) | ( ~n9261 & n9327 ) ;
  assign n9329 = ( x77 & ~n9258 ) | ( x77 & n9328 ) | ( ~n9258 & n9328 ) ;
  assign n9330 = ( x78 & ~n9295 ) | ( x78 & n9329 ) | ( ~n9295 & n9329 ) ;
  assign n9331 = ( x79 & ~n9292 ) | ( x79 & n9330 ) | ( ~n9292 & n9330 ) ;
  assign n9332 = ( x80 & ~n9255 ) | ( x80 & n9331 ) | ( ~n9255 & n9331 ) ;
  assign n9333 = ( x81 & ~n9252 ) | ( x81 & n9332 ) | ( ~n9252 & n9332 ) ;
  assign n9334 = ( x82 & ~n9300 ) | ( x82 & n9333 ) | ( ~n9300 & n9333 ) ;
  assign n9335 = n9318 ^ n9311 ^ x67 ;
  assign n9336 = n9319 ^ n9170 ^ x68 ;
  assign n9337 = n9320 ^ n9168 ^ x69 ;
  assign n9338 = n9321 ^ n9219 ^ x70 ;
  assign n9339 = n9322 ^ n9309 ^ x71 ;
  assign n9340 = n9323 ^ n9306 ^ x72 ;
  assign n9341 = n9325 ^ n9298 ^ x74 ;
  assign n9342 = n9326 ^ n9166 ^ x75 ;
  assign n9343 = n9327 ^ n9261 ^ x76 ;
  assign n9344 = n9328 ^ n9258 ^ x77 ;
  assign n9345 = n9324 ^ n9303 ^ x73 ;
  assign n9346 = n9329 ^ n9295 ^ x78 ;
  assign n9347 = n9330 ^ n9292 ^ x79 ;
  assign n9348 = n9331 ^ n9255 ^ x80 ;
  assign n9349 = n9332 ^ n9252 ^ x81 ;
  assign n9350 = n9333 ^ n9300 ^ x82 ;
  assign n9351 = ( x83 & ~n9249 ) | ( x83 & n9334 ) | ( ~n9249 & n9334 ) ;
  assign n9352 = n9334 ^ n9249 ^ x83 ;
  assign n9353 = ( x84 & ~n9246 ) | ( x84 & n9351 ) | ( ~n9246 & n9351 ) ;
  assign n9354 = ( x85 & ~n9288 ) | ( x85 & n9353 ) | ( ~n9288 & n9353 ) ;
  assign n9355 = ( x86 & ~n9285 ) | ( x86 & n9354 ) | ( ~n9285 & n9354 ) ;
  assign n9356 = ( x87 & ~n9282 ) | ( x87 & n9355 ) | ( ~n9282 & n9355 ) ;
  assign n9357 = ( x88 & ~n9279 ) | ( x88 & n9356 ) | ( ~n9279 & n9356 ) ;
  assign n9358 = ( x89 & ~n9276 ) | ( x89 & n9357 ) | ( ~n9276 & n9357 ) ;
  assign n9359 = ( x90 & ~n9273 ) | ( x90 & n9358 ) | ( ~n9273 & n9358 ) ;
  assign n9360 = ( x91 & ~n9243 ) | ( x91 & n9359 ) | ( ~n9243 & n9359 ) ;
  assign n9361 = ( x92 & ~n9270 ) | ( x92 & n9360 ) | ( ~n9270 & n9360 ) ;
  assign n9362 = ( x93 & ~n9267 ) | ( x93 & n9361 ) | ( ~n9267 & n9361 ) ;
  assign n9363 = ( x94 & ~n9264 ) | ( x94 & n9362 ) | ( ~n9264 & n9362 ) ;
  assign n9364 = ( x95 & ~n9240 ) | ( x95 & n9363 ) | ( ~n9240 & n9363 ) ;
  assign n9365 = ( x96 & ~n9237 ) | ( x96 & n9364 ) | ( ~n9237 & n9364 ) ;
  assign n9366 = ( x97 & ~n9234 ) | ( x97 & n9365 ) | ( ~n9234 & n9365 ) ;
  assign n9367 = ( x98 & ~n9231 ) | ( x98 & n9366 ) | ( ~n9231 & n9366 ) ;
  assign n9368 = ( x99 & ~n9228 ) | ( x99 & n9367 ) | ( ~n9228 & n9367 ) ;
  assign n9369 = ( x100 & ~n9225 ) | ( x100 & n9368 ) | ( ~n9225 & n9368 ) ;
  assign n9370 = ( x101 & ~n9222 ) | ( x101 & n9369 ) | ( ~n9222 & n9369 ) ;
  assign n9371 = ( x102 & ~n9182 ) | ( x102 & n9370 ) | ( ~n9182 & n9370 ) ;
  assign n9372 = ( x103 & ~n9202 ) | ( x103 & n9371 ) | ( ~n9202 & n9371 ) ;
  assign n9373 = ( x104 & ~n9207 ) | ( x104 & n9372 ) | ( ~n9207 & n9372 ) ;
  assign n9374 = ( x105 & ~n9176 ) | ( x105 & n9373 ) | ( ~n9176 & n9373 ) ;
  assign n9375 = ( x106 & ~n9211 ) | ( x106 & n9374 ) | ( ~n9211 & n9374 ) ;
  assign n9376 = ( x107 & ~n9215 ) | ( x107 & n9375 ) | ( ~n9215 & n9375 ) ;
  assign n9377 = ( x108 & ~n9206 ) | ( x108 & n9376 ) | ( ~n9206 & n9376 ) ;
  assign n9378 = ( x109 & ~n9217 ) | ( x109 & n9377 ) | ( ~n9217 & n9377 ) ;
  assign n9379 = ( x110 & ~n9213 ) | ( x110 & n9378 ) | ( ~n9213 & n9378 ) ;
  assign n9380 = ( x111 & ~n9218 ) | ( x111 & n9379 ) | ( ~n9218 & n9379 ) ;
  assign n9381 = ( x112 & ~n9198 ) | ( x112 & n9380 ) | ( ~n9198 & n9380 ) ;
  assign n9382 = ( x113 & ~n9194 ) | ( x113 & n9381 ) | ( ~n9194 & n9381 ) ;
  assign n9383 = ( x114 & ~n9214 ) | ( x114 & n9382 ) | ( ~n9214 & n9382 ) ;
  assign n9384 = ( x115 & ~n9204 ) | ( x115 & n9383 ) | ( ~n9204 & n9383 ) ;
  assign n9385 = ( x116 & ~n9164 ) | ( x116 & n9384 ) | ( ~n9164 & n9384 ) ;
  assign n9386 = ( x117 & ~n9161 ) | ( x117 & n9385 ) | ( ~n9161 & n9385 ) ;
  assign n9387 = ( x118 & ~n9158 ) | ( x118 & n9386 ) | ( ~n9158 & n9386 ) ;
  assign n9388 = ( x119 & ~n9155 ) | ( x119 & n9387 ) | ( ~n9155 & n9387 ) ;
  assign n9389 = ( x120 & ~n9152 ) | ( x120 & n9388 ) | ( ~n9152 & n9388 ) ;
  assign n9390 = ( x121 & ~n9149 ) | ( x121 & n9389 ) | ( ~n9149 & n9389 ) ;
  assign n9391 = ( x122 & ~n9146 ) | ( x122 & n9390 ) | ( ~n9146 & n9390 ) ;
  assign n9392 = ( x123 & ~n9143 ) | ( x123 & n9391 ) | ( ~n9143 & n9391 ) ;
  assign n9393 = ( x124 & ~n9140 ) | ( x124 & n9392 ) | ( ~n9140 & n9392 ) ;
  assign n9394 = ( x125 & ~n9137 ) | ( x125 & n9393 ) | ( ~n9137 & n9393 ) ;
  assign n9395 = ( x126 & ~n9174 ) | ( x126 & n9394 ) | ( ~n9174 & n9394 ) ;
  assign n9396 = x127 | n9395 ;
  assign n9397 = n147 | n9394 ;
  assign n9398 = ( n9174 & n9396 ) | ( n9174 & ~n9397 ) | ( n9396 & ~n9397 ) ;
  assign n9399 = n9396 ^ n9336 ^ 1'b0 ;
  assign n9400 = ( n9170 & n9336 ) | ( n9170 & n9399 ) | ( n9336 & n9399 ) ;
  assign n9401 = n9396 ^ n9350 ^ 1'b0 ;
  assign n9402 = n9396 ^ n9335 ^ 1'b0 ;
  assign n9403 = ( n9300 & n9350 ) | ( n9300 & n9401 ) | ( n9350 & n9401 ) ;
  assign n9404 = n9396 ^ n9352 ^ 1'b0 ;
  assign n9405 = ( n9249 & n9352 ) | ( n9249 & n9404 ) | ( n9352 & n9404 ) ;
  assign n9406 = n9396 ^ n9348 ^ 1'b0 ;
  assign n9407 = n9396 ^ n9315 ^ 1'b0 ;
  assign n9408 = ( n9255 & n9348 ) | ( n9255 & n9406 ) | ( n9348 & n9406 ) ;
  assign n9409 = ( n9314 & n9315 ) | ( n9314 & n9407 ) | ( n9315 & n9407 ) ;
  assign n9410 = n9396 ^ n9317 ^ 1'b0 ;
  assign n9411 = ( n9190 & n9317 ) | ( n9190 & n9410 ) | ( n9317 & n9410 ) ;
  assign n9412 = ( n9311 & n9335 ) | ( n9311 & n9402 ) | ( n9335 & n9402 ) ;
  assign n9413 = n9351 ^ n9246 ^ x84 ;
  assign n9414 = n9413 ^ n9396 ^ 1'b0 ;
  assign n9415 = ( n9246 & n9413 ) | ( n9246 & n9414 ) | ( n9413 & n9414 ) ;
  assign n9416 = n9396 ^ n9349 ^ 1'b0 ;
  assign n9417 = ( n9252 & n9349 ) | ( n9252 & n9416 ) | ( n9349 & n9416 ) ;
  assign n9418 = n9396 ^ n9347 ^ 1'b0 ;
  assign n9419 = ( n9292 & n9347 ) | ( n9292 & n9418 ) | ( n9347 & n9418 ) ;
  assign n9420 = n9396 ^ n9346 ^ 1'b0 ;
  assign n9421 = ( n9295 & n9346 ) | ( n9295 & n9420 ) | ( n9346 & n9420 ) ;
  assign n9422 = n9396 ^ n9344 ^ 1'b0 ;
  assign n9423 = ( n9258 & n9344 ) | ( n9258 & n9422 ) | ( n9344 & n9422 ) ;
  assign n9424 = n9396 ^ n9343 ^ 1'b0 ;
  assign n9425 = ( n9261 & n9343 ) | ( n9261 & n9424 ) | ( n9343 & n9424 ) ;
  assign n9426 = n9396 ^ n9342 ^ 1'b0 ;
  assign n9427 = ( n9166 & n9342 ) | ( n9166 & n9426 ) | ( n9342 & n9426 ) ;
  assign n9428 = n9396 ^ n9341 ^ 1'b0 ;
  assign n9429 = ( n9298 & n9341 ) | ( n9298 & n9428 ) | ( n9341 & n9428 ) ;
  assign n9430 = n9396 ^ n9345 ^ 1'b0 ;
  assign n9431 = ( n9303 & n9345 ) | ( n9303 & n9430 ) | ( n9345 & n9430 ) ;
  assign n9432 = n9396 ^ n9340 ^ 1'b0 ;
  assign n9433 = ( n9306 & n9340 ) | ( n9306 & n9432 ) | ( n9340 & n9432 ) ;
  assign n9434 = n9396 ^ n9339 ^ 1'b0 ;
  assign n9435 = ( n9309 & n9339 ) | ( n9309 & n9434 ) | ( n9339 & n9434 ) ;
  assign n9436 = n9396 ^ n9338 ^ 1'b0 ;
  assign n9437 = ( n9219 & n9338 ) | ( n9219 & n9436 ) | ( n9338 & n9436 ) ;
  assign n9438 = n9396 ^ n9337 ^ 1'b0 ;
  assign n9439 = ( n9168 & n9337 ) | ( n9168 & n9438 ) | ( n9337 & n9438 ) ;
  assign n9440 = ~x0 & x64 ;
  assign n9441 = x64 & n9396 ;
  assign n9442 = n9441 ^ x64 ^ x1 ;
  assign n9443 = ( x65 & n9440 ) | ( x65 & ~n9442 ) | ( n9440 & ~n9442 ) ;
  assign n9444 = ( x66 & ~n9409 ) | ( x66 & n9443 ) | ( ~n9409 & n9443 ) ;
  assign n9445 = ( x67 & ~n9411 ) | ( x67 & n9444 ) | ( ~n9411 & n9444 ) ;
  assign n9446 = ( x68 & ~n9412 ) | ( x68 & n9445 ) | ( ~n9412 & n9445 ) ;
  assign n9447 = ( x69 & ~n9400 ) | ( x69 & n9446 ) | ( ~n9400 & n9446 ) ;
  assign n9448 = ( x70 & ~n9439 ) | ( x70 & n9447 ) | ( ~n9439 & n9447 ) ;
  assign n9449 = ( x71 & ~n9437 ) | ( x71 & n9448 ) | ( ~n9437 & n9448 ) ;
  assign n9450 = ( x72 & ~n9435 ) | ( x72 & n9449 ) | ( ~n9435 & n9449 ) ;
  assign n9451 = ( x73 & ~n9433 ) | ( x73 & n9450 ) | ( ~n9433 & n9450 ) ;
  assign n9452 = ( x74 & ~n9431 ) | ( x74 & n9451 ) | ( ~n9431 & n9451 ) ;
  assign n9453 = ( x75 & ~n9429 ) | ( x75 & n9452 ) | ( ~n9429 & n9452 ) ;
  assign n9454 = ( x76 & ~n9427 ) | ( x76 & n9453 ) | ( ~n9427 & n9453 ) ;
  assign n9455 = ( x77 & ~n9425 ) | ( x77 & n9454 ) | ( ~n9425 & n9454 ) ;
  assign n9456 = ( x78 & ~n9423 ) | ( x78 & n9455 ) | ( ~n9423 & n9455 ) ;
  assign n9457 = ( x79 & ~n9421 ) | ( x79 & n9456 ) | ( ~n9421 & n9456 ) ;
  assign n9458 = ( x80 & ~n9419 ) | ( x80 & n9457 ) | ( ~n9419 & n9457 ) ;
  assign n9459 = ( x81 & ~n9408 ) | ( x81 & n9458 ) | ( ~n9408 & n9458 ) ;
  assign n9460 = ( x82 & ~n9417 ) | ( x82 & n9459 ) | ( ~n9417 & n9459 ) ;
  assign n9461 = ( x83 & ~n9403 ) | ( x83 & n9460 ) | ( ~n9403 & n9460 ) ;
  assign n9462 = ( x84 & ~n9405 ) | ( x84 & n9461 ) | ( ~n9405 & n9461 ) ;
  assign n9463 = ( x85 & ~n9415 ) | ( x85 & n9462 ) | ( ~n9415 & n9462 ) ;
  assign n9464 = n9364 ^ n9237 ^ x96 ;
  assign n9465 = n9464 ^ n9396 ^ 1'b0 ;
  assign n9466 = ( n9237 & n9464 ) | ( n9237 & n9465 ) | ( n9464 & n9465 ) ;
  assign n9467 = n9357 ^ n9276 ^ x89 ;
  assign n9468 = n9467 ^ n9396 ^ 1'b0 ;
  assign n9469 = n9353 ^ n9288 ^ x85 ;
  assign n9470 = n9360 ^ n9270 ^ x92 ;
  assign n9471 = n9469 ^ n9396 ^ 1'b0 ;
  assign n9472 = n9359 ^ n9243 ^ x91 ;
  assign n9473 = ( n9288 & n9469 ) | ( n9288 & n9471 ) | ( n9469 & n9471 ) ;
  assign n9474 = n9470 ^ n9396 ^ 1'b0 ;
  assign n9475 = n9354 ^ n9285 ^ x86 ;
  assign n9476 = n9356 ^ n9279 ^ x88 ;
  assign n9477 = n9475 ^ n9396 ^ 1'b0 ;
  assign n9478 = ( x86 & n9463 ) | ( x86 & ~n9473 ) | ( n9463 & ~n9473 ) ;
  assign n9479 = n9476 ^ n9396 ^ 1'b0 ;
  assign n9480 = ( n9276 & n9467 ) | ( n9276 & n9468 ) | ( n9467 & n9468 ) ;
  assign n9481 = n9358 ^ n9273 ^ x90 ;
  assign n9482 = n9362 ^ n9264 ^ x94 ;
  assign n9483 = n9361 ^ n9267 ^ x93 ;
  assign n9484 = ( n9279 & n9476 ) | ( n9279 & n9479 ) | ( n9476 & n9479 ) ;
  assign n9485 = ( n9270 & n9470 ) | ( n9270 & n9474 ) | ( n9470 & n9474 ) ;
  assign n9486 = ( n9285 & n9475 ) | ( n9285 & n9477 ) | ( n9475 & n9477 ) ;
  assign n9487 = n9482 ^ n9396 ^ 1'b0 ;
  assign n9488 = ( n9264 & n9482 ) | ( n9264 & n9487 ) | ( n9482 & n9487 ) ;
  assign n9489 = n9363 ^ n9240 ^ x95 ;
  assign n9490 = n9355 ^ n9282 ^ x87 ;
  assign n9491 = n9489 ^ n9396 ^ 1'b0 ;
  assign n9492 = ( n9240 & n9489 ) | ( n9240 & n9491 ) | ( n9489 & n9491 ) ;
  assign n9493 = n9490 ^ n9396 ^ 1'b0 ;
  assign n9494 = ( n9282 & n9490 ) | ( n9282 & n9493 ) | ( n9490 & n9493 ) ;
  assign n9495 = ( x87 & n9478 ) | ( x87 & ~n9486 ) | ( n9478 & ~n9486 ) ;
  assign n9496 = n9483 ^ n9396 ^ 1'b0 ;
  assign n9497 = ( n9267 & n9483 ) | ( n9267 & n9496 ) | ( n9483 & n9496 ) ;
  assign n9498 = ( x88 & ~n9494 ) | ( x88 & n9495 ) | ( ~n9494 & n9495 ) ;
  assign n9499 = ( x89 & ~n9484 ) | ( x89 & n9498 ) | ( ~n9484 & n9498 ) ;
  assign n9500 = n9472 ^ n9396 ^ 1'b0 ;
  assign n9501 = ( n9243 & n9472 ) | ( n9243 & n9500 ) | ( n9472 & n9500 ) ;
  assign n9502 = n9481 ^ n9396 ^ 1'b0 ;
  assign n9503 = ( x90 & ~n9480 ) | ( x90 & n9499 ) | ( ~n9480 & n9499 ) ;
  assign n9504 = ( n9273 & n9481 ) | ( n9273 & n9502 ) | ( n9481 & n9502 ) ;
  assign n9505 = ( x91 & n9503 ) | ( x91 & ~n9504 ) | ( n9503 & ~n9504 ) ;
  assign n9506 = ( x92 & ~n9501 ) | ( x92 & n9505 ) | ( ~n9501 & n9505 ) ;
  assign n9507 = ( x93 & ~n9485 ) | ( x93 & n9506 ) | ( ~n9485 & n9506 ) ;
  assign n9508 = ( x94 & ~n9497 ) | ( x94 & n9507 ) | ( ~n9497 & n9507 ) ;
  assign n9509 = ( x95 & ~n9488 ) | ( x95 & n9508 ) | ( ~n9488 & n9508 ) ;
  assign n9510 = ( x96 & ~n9492 ) | ( x96 & n9509 ) | ( ~n9492 & n9509 ) ;
  assign n9511 = ( x97 & ~n9466 ) | ( x97 & n9510 ) | ( ~n9466 & n9510 ) ;
  assign n9512 = n9375 ^ n9215 ^ x107 ;
  assign n9513 = n9512 ^ n9396 ^ 1'b0 ;
  assign n9514 = ( n9215 & n9512 ) | ( n9215 & n9513 ) | ( n9512 & n9513 ) ;
  assign n9515 = n9374 ^ n9211 ^ x106 ;
  assign n9516 = n9373 ^ n9176 ^ x105 ;
  assign n9517 = n9516 ^ n9396 ^ 1'b0 ;
  assign n9518 = ( n9176 & n9516 ) | ( n9176 & n9517 ) | ( n9516 & n9517 ) ;
  assign n9519 = n9372 ^ n9207 ^ x104 ;
  assign n9520 = n9519 ^ n9396 ^ 1'b0 ;
  assign n9521 = ( n9207 & n9519 ) | ( n9207 & n9520 ) | ( n9519 & n9520 ) ;
  assign n9522 = n9371 ^ n9202 ^ x103 ;
  assign n9523 = n9522 ^ n9396 ^ 1'b0 ;
  assign n9524 = ( n9202 & n9522 ) | ( n9202 & n9523 ) | ( n9522 & n9523 ) ;
  assign n9525 = n9370 ^ n9182 ^ x102 ;
  assign n9526 = n9525 ^ n9396 ^ 1'b0 ;
  assign n9527 = ( n9182 & n9525 ) | ( n9182 & n9526 ) | ( n9525 & n9526 ) ;
  assign n9528 = n9369 ^ n9222 ^ x101 ;
  assign n9529 = n9528 ^ n9396 ^ 1'b0 ;
  assign n9530 = ( n9222 & n9528 ) | ( n9222 & n9529 ) | ( n9528 & n9529 ) ;
  assign n9531 = n9515 ^ n9396 ^ 1'b0 ;
  assign n9532 = ( n9211 & n9515 ) | ( n9211 & n9531 ) | ( n9515 & n9531 ) ;
  assign n9533 = n9368 ^ n9225 ^ x100 ;
  assign n9534 = n9533 ^ n9396 ^ 1'b0 ;
  assign n9535 = ( n9225 & n9533 ) | ( n9225 & n9534 ) | ( n9533 & n9534 ) ;
  assign n9536 = n9367 ^ n9228 ^ x99 ;
  assign n9537 = n9536 ^ n9396 ^ 1'b0 ;
  assign n9538 = ( n9228 & n9536 ) | ( n9228 & n9537 ) | ( n9536 & n9537 ) ;
  assign n9539 = n9366 ^ n9231 ^ x98 ;
  assign n9540 = n9539 ^ n9396 ^ 1'b0 ;
  assign n9541 = ( n9231 & n9539 ) | ( n9231 & n9540 ) | ( n9539 & n9540 ) ;
  assign n9542 = n9365 ^ n9234 ^ x97 ;
  assign n9543 = n9542 ^ n9396 ^ 1'b0 ;
  assign n9544 = ( n9234 & n9542 ) | ( n9234 & n9543 ) | ( n9542 & n9543 ) ;
  assign n9545 = ( x98 & n9511 ) | ( x98 & ~n9544 ) | ( n9511 & ~n9544 ) ;
  assign n9546 = ( x99 & ~n9541 ) | ( x99 & n9545 ) | ( ~n9541 & n9545 ) ;
  assign n9547 = ( x100 & ~n9538 ) | ( x100 & n9546 ) | ( ~n9538 & n9546 ) ;
  assign n9548 = ( x101 & ~n9535 ) | ( x101 & n9547 ) | ( ~n9535 & n9547 ) ;
  assign n9549 = ( x102 & ~n9530 ) | ( x102 & n9548 ) | ( ~n9530 & n9548 ) ;
  assign n9550 = ( x103 & ~n9527 ) | ( x103 & n9549 ) | ( ~n9527 & n9549 ) ;
  assign n9551 = ( x104 & ~n9524 ) | ( x104 & n9550 ) | ( ~n9524 & n9550 ) ;
  assign n9552 = ( x105 & ~n9521 ) | ( x105 & n9551 ) | ( ~n9521 & n9551 ) ;
  assign n9553 = ( x106 & ~n9518 ) | ( x106 & n9552 ) | ( ~n9518 & n9552 ) ;
  assign n9554 = ( x107 & ~n9532 ) | ( x107 & n9553 ) | ( ~n9532 & n9553 ) ;
  assign n9555 = n9387 ^ n9155 ^ x119 ;
  assign n9556 = n9376 ^ n9206 ^ x108 ;
  assign n9557 = n9383 ^ n9204 ^ x115 ;
  assign n9558 = ( x108 & ~n9514 ) | ( x108 & n9554 ) | ( ~n9514 & n9554 ) ;
  assign n9559 = n9392 ^ n9140 ^ x124 ;
  assign n9560 = n9390 ^ n9146 ^ x122 ;
  assign n9561 = n9560 ^ n9396 ^ 1'b0 ;
  assign n9562 = n9391 ^ n9143 ^ x123 ;
  assign n9563 = n9382 ^ n9214 ^ x114 ;
  assign n9564 = n9388 ^ n9152 ^ x120 ;
  assign n9565 = ( n9146 & n9560 ) | ( n9146 & n9561 ) | ( n9560 & n9561 ) ;
  assign n9566 = n9377 ^ n9217 ^ x109 ;
  assign n9567 = n9555 ^ n9396 ^ 1'b0 ;
  assign n9568 = n9566 ^ n9396 ^ 1'b0 ;
  assign n9569 = ( n9217 & n9566 ) | ( n9217 & n9568 ) | ( n9566 & n9568 ) ;
  assign n9570 = n9556 ^ n9396 ^ 1'b0 ;
  assign n9571 = n9378 ^ n9213 ^ x110 ;
  assign n9572 = ( n9206 & n9556 ) | ( n9206 & n9570 ) | ( n9556 & n9570 ) ;
  assign n9573 = ( x109 & n9558 ) | ( x109 & ~n9572 ) | ( n9558 & ~n9572 ) ;
  assign n9574 = ( x110 & ~n9569 ) | ( x110 & n9573 ) | ( ~n9569 & n9573 ) ;
  assign n9575 = n9379 ^ n9218 ^ x111 ;
  assign n9576 = n9571 ^ n9396 ^ 1'b0 ;
  assign n9577 = n9575 ^ n9396 ^ 1'b0 ;
  assign n9578 = ( n9218 & n9575 ) | ( n9218 & n9577 ) | ( n9575 & n9577 ) ;
  assign n9579 = n9564 ^ n9396 ^ 1'b0 ;
  assign n9580 = n9380 ^ n9198 ^ x112 ;
  assign n9581 = ( n9213 & n9571 ) | ( n9213 & n9576 ) | ( n9571 & n9576 ) ;
  assign n9582 = n9563 ^ n9396 ^ 1'b0 ;
  assign n9583 = ( n9214 & n9563 ) | ( n9214 & n9582 ) | ( n9563 & n9582 ) ;
  assign n9584 = n9386 ^ n9158 ^ x118 ;
  assign n9585 = n9580 ^ n9396 ^ 1'b0 ;
  assign n9586 = ( n9198 & n9580 ) | ( n9198 & n9585 ) | ( n9580 & n9585 ) ;
  assign n9587 = n9385 ^ n9161 ^ x117 ;
  assign n9588 = n9584 ^ n9396 ^ 1'b0 ;
  assign n9589 = n9587 ^ n9396 ^ 1'b0 ;
  assign n9590 = n9393 ^ n9137 ^ x125 ;
  assign n9591 = n9381 ^ n9194 ^ x113 ;
  assign n9592 = n9590 ^ n9396 ^ 1'b0 ;
  assign n9593 = ( x111 & n9574 ) | ( x111 & ~n9581 ) | ( n9574 & ~n9581 ) ;
  assign n9594 = n9557 ^ n9396 ^ 1'b0 ;
  assign n9595 = n9389 ^ n9149 ^ x121 ;
  assign n9596 = n9384 ^ n9164 ^ x116 ;
  assign n9597 = n9591 ^ n9396 ^ 1'b0 ;
  assign n9598 = ( n9194 & n9591 ) | ( n9194 & n9597 ) | ( n9591 & n9597 ) ;
  assign n9599 = ( x112 & ~n9578 ) | ( x112 & n9593 ) | ( ~n9578 & n9593 ) ;
  assign n9600 = n9559 ^ n9396 ^ 1'b0 ;
  assign n9601 = ( n9161 & n9587 ) | ( n9161 & n9589 ) | ( n9587 & n9589 ) ;
  assign n9602 = ( x113 & ~n9586 ) | ( x113 & n9599 ) | ( ~n9586 & n9599 ) ;
  assign n9603 = n9596 ^ n9396 ^ 1'b0 ;
  assign n9604 = ( n9155 & n9555 ) | ( n9155 & n9567 ) | ( n9555 & n9567 ) ;
  assign n9605 = n9595 ^ n9396 ^ 1'b0 ;
  assign n9606 = ( x114 & ~n9598 ) | ( x114 & n9602 ) | ( ~n9598 & n9602 ) ;
  assign n9607 = ( x115 & ~n9583 ) | ( x115 & n9606 ) | ( ~n9583 & n9606 ) ;
  assign n9608 = ( n9152 & n9564 ) | ( n9152 & n9579 ) | ( n9564 & n9579 ) ;
  assign n9609 = ( n9149 & n9595 ) | ( n9149 & n9605 ) | ( n9595 & n9605 ) ;
  assign n9610 = ( n9204 & n9557 ) | ( n9204 & n9594 ) | ( n9557 & n9594 ) ;
  assign n9611 = n9562 ^ n9396 ^ 1'b0 ;
  assign n9612 = ( n9143 & n9562 ) | ( n9143 & n9611 ) | ( n9562 & n9611 ) ;
  assign n9613 = ( n9164 & n9596 ) | ( n9164 & n9603 ) | ( n9596 & n9603 ) ;
  assign n9614 = ( n9140 & n9559 ) | ( n9140 & n9600 ) | ( n9559 & n9600 ) ;
  assign n9615 = ( n9137 & n9590 ) | ( n9137 & n9592 ) | ( n9590 & n9592 ) ;
  assign n9616 = ( x116 & n9607 ) | ( x116 & ~n9610 ) | ( n9607 & ~n9610 ) ;
  assign n9617 = ( x117 & ~n9613 ) | ( x117 & n9616 ) | ( ~n9613 & n9616 ) ;
  assign n9618 = ( x118 & ~n9601 ) | ( x118 & n9617 ) | ( ~n9601 & n9617 ) ;
  assign n9619 = ( n9158 & n9584 ) | ( n9158 & n9588 ) | ( n9584 & n9588 ) ;
  assign n9620 = ( x119 & n9618 ) | ( x119 & ~n9619 ) | ( n9618 & ~n9619 ) ;
  assign n9621 = ( x120 & ~n9604 ) | ( x120 & n9620 ) | ( ~n9604 & n9620 ) ;
  assign n9622 = ( x121 & ~n9608 ) | ( x121 & n9621 ) | ( ~n9608 & n9621 ) ;
  assign n9623 = ( x122 & ~n9609 ) | ( x122 & n9622 ) | ( ~n9609 & n9622 ) ;
  assign n9624 = ( x123 & ~n9565 ) | ( x123 & n9623 ) | ( ~n9565 & n9623 ) ;
  assign n9625 = ( x124 & ~n9612 ) | ( x124 & n9624 ) | ( ~n9612 & n9624 ) ;
  assign n9626 = ( x125 & ~n9614 ) | ( x125 & n9625 ) | ( ~n9614 & n9625 ) ;
  assign n9627 = ( x126 & ~n9615 ) | ( x126 & n9626 ) | ( ~n9615 & n9626 ) ;
  assign n9628 = ( x127 & ~n9398 ) | ( x127 & n9627 ) | ( ~n9398 & n9627 ) ;
  assign n9629 = x64 & n6415 ;
  assign n9630 = n9629 ^ x64 ^ x13 ;
  assign n9631 = n9630 ^ n6757 ^ x65 ;
  assign n9632 = ( x65 & n6757 ) | ( x65 & n9631 ) | ( n6757 & n9631 ) ;
  assign n9633 = n9632 ^ n6453 ^ x66 ;
  assign n9634 = ( x66 & n9632 ) | ( x66 & n9633 ) | ( n9632 & n9633 ) ;
  assign n9635 = ( x67 & ~n6451 ) | ( x67 & n9634 ) | ( ~n6451 & n9634 ) ;
  assign n9636 = ( x68 & ~n6506 ) | ( x68 & n9635 ) | ( ~n6506 & n9635 ) ;
  assign n9637 = ( x69 & ~n6503 ) | ( x69 & n9636 ) | ( ~n6503 & n9636 ) ;
  assign n9638 = ( x70 & ~n6449 ) | ( x70 & n9637 ) | ( ~n6449 & n9637 ) ;
  assign n9639 = ( x71 & ~n6500 ) | ( x71 & n9638 ) | ( ~n6500 & n9638 ) ;
  assign n9640 = ( x72 & ~n6497 ) | ( x72 & n9639 ) | ( ~n6497 & n9639 ) ;
  assign n9641 = ( x73 & ~n6447 ) | ( x73 & n9640 ) | ( ~n6447 & n9640 ) ;
  assign n9642 = ( x74 & ~n6445 ) | ( x74 & n9641 ) | ( ~n6445 & n9641 ) ;
  assign n9643 = ( x75 & ~n6494 ) | ( x75 & n9642 ) | ( ~n6494 & n9642 ) ;
  assign n9644 = ( x76 & ~n6491 ) | ( x76 & n9643 ) | ( ~n6491 & n9643 ) ;
  assign n9645 = ( x77 & ~n6488 ) | ( x77 & n9644 ) | ( ~n6488 & n9644 ) ;
  assign n9646 = n9638 ^ n6500 ^ x71 ;
  assign n9647 = ( x78 & ~n6485 ) | ( x78 & n9645 ) | ( ~n6485 & n9645 ) ;
  assign n9648 = ( x79 & ~n6482 ) | ( x79 & n9647 ) | ( ~n6482 & n9647 ) ;
  assign n9649 = ( x80 & ~n6443 ) | ( x80 & n9648 ) | ( ~n6443 & n9648 ) ;
  assign n9650 = ( x81 & ~n6441 ) | ( x81 & n9649 ) | ( ~n6441 & n9649 ) ;
  assign n9651 = ( x82 & ~n6479 ) | ( x82 & n9650 ) | ( ~n6479 & n9650 ) ;
  assign n9652 = ( x83 & ~n6439 ) | ( x83 & n9651 ) | ( ~n6439 & n9651 ) ;
  assign n9653 = ( x84 & ~n6476 ) | ( x84 & n9652 ) | ( ~n6476 & n9652 ) ;
  assign n9654 = ( x85 & ~n6437 ) | ( x85 & n9653 ) | ( ~n6437 & n9653 ) ;
  assign n9655 = ( x86 & ~n6435 ) | ( x86 & n9654 ) | ( ~n6435 & n9654 ) ;
  assign n9656 = ( x87 & ~n6473 ) | ( x87 & n9655 ) | ( ~n6473 & n9655 ) ;
  assign n9657 = ( x88 & ~n6433 ) | ( x88 & n9656 ) | ( ~n6433 & n9656 ) ;
  assign n9658 = ( x89 & ~n6431 ) | ( x89 & n9657 ) | ( ~n6431 & n9657 ) ;
  assign n9659 = ( x90 & ~n6429 ) | ( x90 & n9658 ) | ( ~n6429 & n9658 ) ;
  assign n9660 = ( x91 & ~n6427 ) | ( x91 & n9659 ) | ( ~n6427 & n9659 ) ;
  assign n9661 = ( x92 & ~n6470 ) | ( x92 & n9660 ) | ( ~n6470 & n9660 ) ;
  assign n9662 = ( x93 & ~n6467 ) | ( x93 & n9661 ) | ( ~n6467 & n9661 ) ;
  assign n9663 = n9662 ^ n6548 ^ x94 ;
  assign n9664 = n9648 ^ n6443 ^ x80 ;
  assign n9665 = n9639 ^ n6497 ^ x72 ;
  assign n9666 = n9642 ^ n6494 ^ x75 ;
  assign n9667 = n9651 ^ n6439 ^ x83 ;
  assign n9668 = n9652 ^ n6476 ^ x84 ;
  assign n9669 = n9643 ^ n6491 ^ x76 ;
  assign n9670 = n9654 ^ n6435 ^ x86 ;
  assign n9671 = n9644 ^ n6488 ^ x77 ;
  assign n9672 = n9661 ^ n6467 ^ x93 ;
  assign n9673 = n9657 ^ n6431 ^ x89 ;
  assign n9674 = ( x94 & ~n6548 ) | ( x94 & n9662 ) | ( ~n6548 & n9662 ) ;
  assign n9675 = n9659 ^ n6427 ^ x91 ;
  assign n9676 = n9660 ^ n6470 ^ x92 ;
  assign n9677 = n9645 ^ n6485 ^ x78 ;
  assign n9678 = n9636 ^ n6503 ^ x69 ;
  assign n9679 = ( x95 & ~n6425 ) | ( x95 & n9674 ) | ( ~n6425 & n9674 ) ;
  assign n9680 = n9635 ^ n6506 ^ x68 ;
  assign n9681 = ( x96 & ~n6423 ) | ( x96 & n9679 ) | ( ~n6423 & n9679 ) ;
  assign n9682 = ( x97 & ~n6545 ) | ( x97 & n9681 ) | ( ~n6545 & n9681 ) ;
  assign n9683 = ( x98 & ~n6542 ) | ( x98 & n9682 ) | ( ~n6542 & n9682 ) ;
  assign n9684 = ( x99 & ~n6421 ) | ( x99 & n9683 ) | ( ~n6421 & n9683 ) ;
  assign n9685 = ( x100 & ~n6539 ) | ( x100 & n9684 ) | ( ~n6539 & n9684 ) ;
  assign n9686 = ( x101 & ~n6536 ) | ( x101 & n9685 ) | ( ~n6536 & n9685 ) ;
  assign n9687 = ( x102 & ~n6533 ) | ( x102 & n9686 ) | ( ~n6533 & n9686 ) ;
  assign n9688 = ( x103 & ~n6530 ) | ( x103 & n9687 ) | ( ~n6530 & n9687 ) ;
  assign n9689 = ( x104 & ~n6527 ) | ( x104 & n9688 ) | ( ~n6527 & n9688 ) ;
  assign n9690 = ( x105 & ~n6418 ) | ( x105 & n9689 ) | ( ~n6418 & n9689 ) ;
  assign n9691 = ( x106 & ~n6524 ) | ( x106 & n9690 ) | ( ~n6524 & n9690 ) ;
  assign n9692 = ( x107 & ~n6521 ) | ( x107 & n9691 ) | ( ~n6521 & n9691 ) ;
  assign n9693 = ( x108 & ~n6518 ) | ( x108 & n9692 ) | ( ~n6518 & n9692 ) ;
  assign n9694 = ( x109 & ~n6515 ) | ( x109 & n9693 ) | ( ~n6515 & n9693 ) ;
  assign n9695 = ( x110 & ~n6512 ) | ( x110 & n9694 ) | ( ~n6512 & n9694 ) ;
  assign n9696 = ( x111 & ~n6509 ) | ( x111 & n9695 ) | ( ~n6509 & n9695 ) ;
  assign n9697 = ( x112 & ~n6464 ) | ( x112 & n9696 ) | ( ~n6464 & n9696 ) ;
  assign n9698 = ( x113 & ~n6461 ) | ( x113 & n9697 ) | ( ~n6461 & n9697 ) ;
  assign n9699 = ( x114 & ~n6458 ) | ( x114 & n9698 ) | ( ~n6458 & n9698 ) ;
  assign n9700 = ( x115 & ~n6455 ) | ( x115 & n9699 ) | ( ~n6455 & n9699 ) ;
  assign n9701 = n6965 | n9700 ;
  assign n9702 = ( x12 & ~n9700 ) | ( x12 & n9701 ) | ( ~n9700 & n9701 ) ;
  assign n9703 = ~n6970 & n9702 ;
  assign n9704 = ( n9701 & n9702 ) | ( n9701 & n9703 ) | ( n9702 & n9703 ) ;
  assign n9705 = n174 | n9700 ;
  assign n9706 = n9705 ^ n6439 ^ 1'b0 ;
  assign n9707 = n9705 ^ n6485 ^ 1'b0 ;
  assign n9708 = ( n6485 & n9677 ) | ( n6485 & ~n9707 ) | ( n9677 & ~n9707 ) ;
  assign n9709 = n9705 ^ n6548 ^ 1'b0 ;
  assign n9710 = n9705 ^ n6506 ^ 1'b0 ;
  assign n9711 = ( n6506 & n9680 ) | ( n6506 & ~n9710 ) | ( n9680 & ~n9710 ) ;
  assign n9712 = n9705 ^ n6476 ^ 1'b0 ;
  assign n9713 = n9705 ^ n9631 ^ 1'b0 ;
  assign n9714 = ( n9630 & n9631 ) | ( n9630 & n9713 ) | ( n9631 & n9713 ) ;
  assign n9715 = n9705 ^ n6467 ^ 1'b0 ;
  assign n9716 = n9705 ^ n6443 ^ 1'b0 ;
  assign n9717 = ( n6467 & n9672 ) | ( n6467 & ~n9715 ) | ( n9672 & ~n9715 ) ;
  assign n9718 = ( n6439 & n9667 ) | ( n6439 & ~n9706 ) | ( n9667 & ~n9706 ) ;
  assign n9719 = ( n6443 & n9664 ) | ( n6443 & ~n9716 ) | ( n9664 & ~n9716 ) ;
  assign n9720 = ( n6548 & n9663 ) | ( n6548 & ~n9709 ) | ( n9663 & ~n9709 ) ;
  assign n9721 = ( n6476 & n9668 ) | ( n6476 & ~n9712 ) | ( n9668 & ~n9712 ) ;
  assign n9722 = n9705 ^ n6497 ^ 1'b0 ;
  assign n9723 = ( n6497 & n9665 ) | ( n6497 & ~n9722 ) | ( n9665 & ~n9722 ) ;
  assign n9724 = n9705 ^ n6494 ^ 1'b0 ;
  assign n9725 = n9705 ^ n6503 ^ 1'b0 ;
  assign n9726 = n9705 ^ n6488 ^ 1'b0 ;
  assign n9727 = n9705 ^ n6500 ^ 1'b0 ;
  assign n9728 = ( n6500 & n9646 ) | ( n6500 & ~n9727 ) | ( n9646 & ~n9727 ) ;
  assign n9729 = ( n6488 & n9671 ) | ( n6488 & ~n9726 ) | ( n9671 & ~n9726 ) ;
  assign n9730 = n9705 ^ n9633 ^ 1'b0 ;
  assign n9731 = ( n6453 & n9633 ) | ( n6453 & n9730 ) | ( n9633 & n9730 ) ;
  assign n9732 = ( n6494 & n9666 ) | ( n6494 & ~n9724 ) | ( n9666 & ~n9724 ) ;
  assign n9733 = ( n6503 & n9678 ) | ( n6503 & ~n9725 ) | ( n9678 & ~n9725 ) ;
  assign n9734 = n9705 ^ n6435 ^ 1'b0 ;
  assign n9735 = n9705 ^ n6427 ^ 1'b0 ;
  assign n9736 = n9705 ^ n6470 ^ 1'b0 ;
  assign n9737 = ( n6470 & n9676 ) | ( n6470 & ~n9736 ) | ( n9676 & ~n9736 ) ;
  assign n9738 = ( n6427 & n9675 ) | ( n6427 & ~n9735 ) | ( n9675 & ~n9735 ) ;
  assign n9739 = n9705 ^ n6431 ^ 1'b0 ;
  assign n9740 = n9705 ^ n6491 ^ 1'b0 ;
  assign n9741 = ( n6431 & n9673 ) | ( n6431 & ~n9739 ) | ( n9673 & ~n9739 ) ;
  assign n9742 = ( n6435 & n9670 ) | ( n6435 & ~n9734 ) | ( n9670 & ~n9734 ) ;
  assign n9743 = ( n6491 & n9669 ) | ( n6491 & ~n9740 ) | ( n9669 & ~n9740 ) ;
  assign n9744 = n9698 ^ n6458 ^ x114 ;
  assign n9745 = n9705 ^ n6458 ^ 1'b0 ;
  assign n9746 = ( n6458 & n9744 ) | ( n6458 & ~n9745 ) | ( n9744 & ~n9745 ) ;
  assign n9747 = n9697 ^ n6461 ^ x113 ;
  assign n9748 = n9705 ^ n6461 ^ 1'b0 ;
  assign n9749 = ( n6461 & n9747 ) | ( n6461 & ~n9748 ) | ( n9747 & ~n9748 ) ;
  assign n9750 = n9682 ^ n6542 ^ x98 ;
  assign n9751 = n9705 ^ n6542 ^ 1'b0 ;
  assign n9752 = ( n6542 & n9750 ) | ( n6542 & ~n9751 ) | ( n9750 & ~n9751 ) ;
  assign n9753 = n9681 ^ n6545 ^ x97 ;
  assign n9754 = n9705 ^ n6545 ^ 1'b0 ;
  assign n9755 = ( n6545 & n9753 ) | ( n6545 & ~n9754 ) | ( n9753 & ~n9754 ) ;
  assign n9756 = n9679 ^ n6423 ^ x96 ;
  assign n9757 = n9705 ^ n6423 ^ 1'b0 ;
  assign n9758 = ( n6423 & n9756 ) | ( n6423 & ~n9757 ) | ( n9756 & ~n9757 ) ;
  assign n9759 = n9674 ^ n6425 ^ x95 ;
  assign n9760 = n9705 ^ n6425 ^ 1'b0 ;
  assign n9761 = ( n6425 & n9759 ) | ( n6425 & ~n9760 ) | ( n9759 & ~n9760 ) ;
  assign n9762 = n9658 ^ n6429 ^ x90 ;
  assign n9763 = n9705 ^ n6429 ^ 1'b0 ;
  assign n9764 = ( n6429 & n9762 ) | ( n6429 & ~n9763 ) | ( n9762 & ~n9763 ) ;
  assign n9765 = n9656 ^ n6433 ^ x88 ;
  assign n9766 = n9705 ^ n6433 ^ 1'b0 ;
  assign n9767 = ( n6433 & n9765 ) | ( n6433 & ~n9766 ) | ( n9765 & ~n9766 ) ;
  assign n9768 = n9655 ^ n6473 ^ x87 ;
  assign n9769 = n9705 ^ n6473 ^ 1'b0 ;
  assign n9770 = ( n6473 & n9768 ) | ( n6473 & ~n9769 ) | ( n9768 & ~n9769 ) ;
  assign n9771 = n9653 ^ n6437 ^ x85 ;
  assign n9772 = n9705 ^ n6437 ^ 1'b0 ;
  assign n9773 = ( n6437 & n9771 ) | ( n6437 & ~n9772 ) | ( n9771 & ~n9772 ) ;
  assign n9774 = n9650 ^ n6479 ^ x82 ;
  assign n9775 = n9705 ^ n6479 ^ 1'b0 ;
  assign n9776 = ( n6479 & n9774 ) | ( n6479 & ~n9775 ) | ( n9774 & ~n9775 ) ;
  assign n9777 = n9649 ^ n6441 ^ x81 ;
  assign n9778 = n9705 ^ n6441 ^ 1'b0 ;
  assign n9779 = ( n6441 & n9777 ) | ( n6441 & ~n9778 ) | ( n9777 & ~n9778 ) ;
  assign n9780 = n9647 ^ n6482 ^ x79 ;
  assign n9781 = n9705 ^ n6482 ^ 1'b0 ;
  assign n9782 = ( n6482 & n9780 ) | ( n6482 & ~n9781 ) | ( n9780 & ~n9781 ) ;
  assign n9783 = n9641 ^ n6445 ^ x74 ;
  assign n9784 = n9705 ^ n6445 ^ 1'b0 ;
  assign n9785 = ( n6445 & n9783 ) | ( n6445 & ~n9784 ) | ( n9783 & ~n9784 ) ;
  assign n9786 = n9640 ^ n6447 ^ x73 ;
  assign n9787 = n9705 ^ n6447 ^ 1'b0 ;
  assign n9788 = ( n6447 & n9786 ) | ( n6447 & ~n9787 ) | ( n9786 & ~n9787 ) ;
  assign n9789 = n9637 ^ n6449 ^ x70 ;
  assign n9790 = n9705 ^ n6449 ^ 1'b0 ;
  assign n9791 = ( n6449 & n9789 ) | ( n6449 & ~n9790 ) | ( n9789 & ~n9790 ) ;
  assign n9792 = n9634 ^ n6451 ^ x67 ;
  assign n9793 = n9705 ^ n6451 ^ 1'b0 ;
  assign n9794 = ( n6451 & n9792 ) | ( n6451 & ~n9793 ) | ( n9792 & ~n9793 ) ;
  assign n9795 = n9696 ^ n6464 ^ x112 ;
  assign n9796 = n9705 ^ n6464 ^ 1'b0 ;
  assign n9797 = ( n6464 & n9795 ) | ( n6464 & ~n9796 ) | ( n9795 & ~n9796 ) ;
  assign n9798 = n9695 ^ n6509 ^ x111 ;
  assign n9799 = n9694 ^ n6512 ^ x110 ;
  assign n9800 = n9705 ^ n6512 ^ 1'b0 ;
  assign n9801 = ( n6512 & n9799 ) | ( n6512 & ~n9800 ) | ( n9799 & ~n9800 ) ;
  assign n9802 = n9693 ^ n6515 ^ x109 ;
  assign n9803 = n9705 ^ n6509 ^ 1'b0 ;
  assign n9804 = ( n6509 & n9798 ) | ( n6509 & ~n9803 ) | ( n9798 & ~n9803 ) ;
  assign n9805 = n9705 ^ n6515 ^ 1'b0 ;
  assign n9806 = ( n6515 & n9802 ) | ( n6515 & ~n9805 ) | ( n9802 & ~n9805 ) ;
  assign n9807 = n9692 ^ n6518 ^ x108 ;
  assign n9808 = n9705 ^ n6518 ^ 1'b0 ;
  assign n9809 = ( n6518 & n9807 ) | ( n6518 & ~n9808 ) | ( n9807 & ~n9808 ) ;
  assign n9810 = n9691 ^ n6521 ^ x107 ;
  assign n9811 = n9705 ^ n6521 ^ 1'b0 ;
  assign n9812 = ( n6521 & n9810 ) | ( n6521 & ~n9811 ) | ( n9810 & ~n9811 ) ;
  assign n9813 = n9690 ^ n6524 ^ x106 ;
  assign n9814 = n9705 ^ n6524 ^ 1'b0 ;
  assign n9815 = ( n6524 & n9813 ) | ( n6524 & ~n9814 ) | ( n9813 & ~n9814 ) ;
  assign n9816 = n9689 ^ n6418 ^ x105 ;
  assign n9817 = n9705 ^ n6418 ^ 1'b0 ;
  assign n9818 = ( n6418 & n9816 ) | ( n6418 & ~n9817 ) | ( n9816 & ~n9817 ) ;
  assign n9819 = n9688 ^ n6527 ^ x104 ;
  assign n9820 = n9705 ^ n6527 ^ 1'b0 ;
  assign n9821 = ( n6527 & n9819 ) | ( n6527 & ~n9820 ) | ( n9819 & ~n9820 ) ;
  assign n9822 = n9687 ^ n6530 ^ x103 ;
  assign n9823 = n9705 ^ n6530 ^ 1'b0 ;
  assign n9824 = ( n6530 & n9822 ) | ( n6530 & ~n9823 ) | ( n9822 & ~n9823 ) ;
  assign n9825 = n9686 ^ n6533 ^ x102 ;
  assign n9826 = n9705 ^ n6533 ^ 1'b0 ;
  assign n9827 = ( n6533 & n9825 ) | ( n6533 & ~n9826 ) | ( n9825 & ~n9826 ) ;
  assign n9828 = n9685 ^ n6536 ^ x101 ;
  assign n9829 = n9705 ^ n6536 ^ 1'b0 ;
  assign n9830 = ( n6536 & n9828 ) | ( n6536 & ~n9829 ) | ( n9828 & ~n9829 ) ;
  assign n9831 = n9684 ^ n6539 ^ x100 ;
  assign n9832 = n9705 ^ n6539 ^ 1'b0 ;
  assign n9833 = ( n6539 & n9831 ) | ( n6539 & ~n9832 ) | ( n9831 & ~n9832 ) ;
  assign n9834 = n9683 ^ n6421 ^ x99 ;
  assign n9835 = n9705 ^ n6421 ^ 1'b0 ;
  assign n9836 = ( n6421 & n9834 ) | ( n6421 & ~n9835 ) | ( n9834 & ~n9835 ) ;
  assign n9837 = n6455 & n9705 ;
  assign n9838 = n174 & n6455 ;
  assign n9839 = n9704 ^ n6967 ^ x65 ;
  assign n9840 = ( x65 & n6967 ) | ( x65 & n9839 ) | ( n6967 & n9839 ) ;
  assign n9841 = n9840 ^ n9714 ^ x66 ;
  assign n9842 = ( x66 & n9840 ) | ( x66 & n9841 ) | ( n9840 & n9841 ) ;
  assign n9843 = ( x67 & ~n9731 ) | ( x67 & n9842 ) | ( ~n9731 & n9842 ) ;
  assign n9844 = ( x68 & ~n9794 ) | ( x68 & n9843 ) | ( ~n9794 & n9843 ) ;
  assign n9845 = ( x69 & ~n9711 ) | ( x69 & n9844 ) | ( ~n9711 & n9844 ) ;
  assign n9846 = ( x70 & ~n9733 ) | ( x70 & n9845 ) | ( ~n9733 & n9845 ) ;
  assign n9847 = ( x71 & ~n9791 ) | ( x71 & n9846 ) | ( ~n9791 & n9846 ) ;
  assign n9848 = ( x72 & ~n9728 ) | ( x72 & n9847 ) | ( ~n9728 & n9847 ) ;
  assign n9849 = ( x73 & ~n9723 ) | ( x73 & n9848 ) | ( ~n9723 & n9848 ) ;
  assign n9850 = ( x74 & ~n9788 ) | ( x74 & n9849 ) | ( ~n9788 & n9849 ) ;
  assign n9851 = ( x75 & ~n9785 ) | ( x75 & n9850 ) | ( ~n9785 & n9850 ) ;
  assign n9852 = ( x76 & ~n9732 ) | ( x76 & n9851 ) | ( ~n9732 & n9851 ) ;
  assign n9853 = ( x77 & ~n9743 ) | ( x77 & n9852 ) | ( ~n9743 & n9852 ) ;
  assign n9854 = ( x78 & ~n9729 ) | ( x78 & n9853 ) | ( ~n9729 & n9853 ) ;
  assign n9855 = ( x79 & ~n9708 ) | ( x79 & n9854 ) | ( ~n9708 & n9854 ) ;
  assign n9856 = ( x80 & ~n9782 ) | ( x80 & n9855 ) | ( ~n9782 & n9855 ) ;
  assign n9857 = ( x81 & ~n9719 ) | ( x81 & n9856 ) | ( ~n9719 & n9856 ) ;
  assign n9858 = ( x82 & ~n9779 ) | ( x82 & n9857 ) | ( ~n9779 & n9857 ) ;
  assign n9859 = ( x83 & ~n9776 ) | ( x83 & n9858 ) | ( ~n9776 & n9858 ) ;
  assign n9860 = ( x84 & ~n9718 ) | ( x84 & n9859 ) | ( ~n9718 & n9859 ) ;
  assign n9861 = ( x85 & ~n9721 ) | ( x85 & n9860 ) | ( ~n9721 & n9860 ) ;
  assign n9862 = ( x86 & ~n9773 ) | ( x86 & n9861 ) | ( ~n9773 & n9861 ) ;
  assign n9863 = ( x87 & ~n9742 ) | ( x87 & n9862 ) | ( ~n9742 & n9862 ) ;
  assign n9864 = ( x116 & n171 ) | ( x116 & ~n9837 ) | ( n171 & ~n9837 ) ;
  assign n9865 = n322 | n9837 ;
  assign n9866 = ( x88 & ~n9770 ) | ( x88 & n9863 ) | ( ~n9770 & n9863 ) ;
  assign n9867 = ( x89 & ~n9767 ) | ( x89 & n9866 ) | ( ~n9767 & n9866 ) ;
  assign n9868 = ( x90 & ~n9741 ) | ( x90 & n9867 ) | ( ~n9741 & n9867 ) ;
  assign n9869 = ( x91 & ~n9764 ) | ( x91 & n9868 ) | ( ~n9764 & n9868 ) ;
  assign n9870 = n9863 ^ n9770 ^ x88 ;
  assign n9871 = n9862 ^ n9742 ^ x87 ;
  assign n9872 = n9861 ^ n9773 ^ x86 ;
  assign n9873 = n9860 ^ n9721 ^ x85 ;
  assign n9874 = n9858 ^ n9776 ^ x83 ;
  assign n9875 = n9857 ^ n9779 ^ x82 ;
  assign n9876 = n9856 ^ n9719 ^ x81 ;
  assign n9877 = n9842 ^ n9731 ^ x67 ;
  assign n9878 = n9843 ^ n9794 ^ x68 ;
  assign n9879 = ( x92 & ~n9738 ) | ( x92 & n9869 ) | ( ~n9738 & n9869 ) ;
  assign n9880 = n9869 ^ n9738 ^ x92 ;
  assign n9881 = n9868 ^ n9764 ^ x91 ;
  assign n9882 = n9849 ^ n9788 ^ x74 ;
  assign n9883 = n9852 ^ n9743 ^ x77 ;
  assign n9884 = n9855 ^ n9782 ^ x80 ;
  assign n9885 = n9867 ^ n9741 ^ x90 ;
  assign n9886 = n9845 ^ n9733 ^ x70 ;
  assign n9887 = n174 & n9865 ;
  assign n9888 = ( x93 & ~n9737 ) | ( x93 & n9879 ) | ( ~n9737 & n9879 ) ;
  assign n9889 = ( x94 & ~n9717 ) | ( x94 & n9888 ) | ( ~n9717 & n9888 ) ;
  assign n9890 = n9888 ^ n9717 ^ x94 ;
  assign n9891 = ( x95 & ~n9720 ) | ( x95 & n9889 ) | ( ~n9720 & n9889 ) ;
  assign n9892 = ( x96 & ~n9761 ) | ( x96 & n9891 ) | ( ~n9761 & n9891 ) ;
  assign n9893 = ( x97 & ~n9758 ) | ( x97 & n9892 ) | ( ~n9758 & n9892 ) ;
  assign n9894 = ( x98 & ~n9755 ) | ( x98 & n9893 ) | ( ~n9755 & n9893 ) ;
  assign n9895 = ( x99 & ~n9752 ) | ( x99 & n9894 ) | ( ~n9752 & n9894 ) ;
  assign n9896 = ( x100 & ~n9836 ) | ( x100 & n9895 ) | ( ~n9836 & n9895 ) ;
  assign n9897 = ( x101 & ~n9833 ) | ( x101 & n9896 ) | ( ~n9833 & n9896 ) ;
  assign n9898 = ( x102 & ~n9830 ) | ( x102 & n9897 ) | ( ~n9830 & n9897 ) ;
  assign n9899 = ( x103 & ~n9827 ) | ( x103 & n9898 ) | ( ~n9827 & n9898 ) ;
  assign n9900 = ( x104 & ~n9824 ) | ( x104 & n9899 ) | ( ~n9824 & n9899 ) ;
  assign n9901 = ( x105 & ~n9821 ) | ( x105 & n9900 ) | ( ~n9821 & n9900 ) ;
  assign n9902 = ( x106 & ~n9818 ) | ( x106 & n9901 ) | ( ~n9818 & n9901 ) ;
  assign n9903 = ( x107 & ~n9815 ) | ( x107 & n9902 ) | ( ~n9815 & n9902 ) ;
  assign n9904 = ( x108 & ~n9812 ) | ( x108 & n9903 ) | ( ~n9812 & n9903 ) ;
  assign n9905 = ( x109 & ~n9809 ) | ( x109 & n9904 ) | ( ~n9809 & n9904 ) ;
  assign n9906 = ( x110 & ~n9806 ) | ( x110 & n9905 ) | ( ~n9806 & n9905 ) ;
  assign n9907 = ( x111 & ~n9801 ) | ( x111 & n9906 ) | ( ~n9801 & n9906 ) ;
  assign n9908 = ( x112 & ~n9804 ) | ( x112 & n9907 ) | ( ~n9804 & n9907 ) ;
  assign n9909 = ( x113 & ~n9797 ) | ( x113 & n9908 ) | ( ~n9797 & n9908 ) ;
  assign n9910 = ( x114 & ~n9749 ) | ( x114 & n9909 ) | ( ~n9749 & n9909 ) ;
  assign n9911 = ( x115 & ~n9746 ) | ( x115 & n9910 ) | ( ~n9746 & n9910 ) ;
  assign n9912 = ( ~x116 & n171 ) | ( ~x116 & n9865 ) | ( n171 & n9865 ) ;
  assign n9913 = ( n9864 & ~n9911 ) | ( n9864 & n9912 ) | ( ~n9911 & n9912 ) ;
  assign n9914 = n9911 | n9913 ;
  assign n9915 = ( ~n9865 & n9887 ) | ( ~n9865 & n9914 ) | ( n9887 & n9914 ) ;
  assign n9916 = n9915 ^ n9717 ^ 1'b0 ;
  assign n9917 = ( n9717 & n9890 ) | ( n9717 & ~n9916 ) | ( n9890 & ~n9916 ) ;
  assign n9918 = n9915 ^ n9738 ^ 1'b0 ;
  assign n9919 = ( n9738 & n9880 ) | ( n9738 & ~n9918 ) | ( n9880 & ~n9918 ) ;
  assign n9920 = n9915 ^ n9764 ^ 1'b0 ;
  assign n9921 = ( n9764 & n9881 ) | ( n9764 & ~n9920 ) | ( n9881 & ~n9920 ) ;
  assign n9922 = n9915 ^ n9741 ^ 1'b0 ;
  assign n9923 = ( n9741 & n9885 ) | ( n9741 & ~n9922 ) | ( n9885 & ~n9922 ) ;
  assign n9924 = n9915 ^ n9770 ^ 1'b0 ;
  assign n9925 = ( n9770 & n9870 ) | ( n9770 & ~n9924 ) | ( n9870 & ~n9924 ) ;
  assign n9926 = n9915 ^ n9742 ^ 1'b0 ;
  assign n9927 = ( n9742 & n9871 ) | ( n9742 & ~n9926 ) | ( n9871 & ~n9926 ) ;
  assign n9928 = n9915 ^ n9773 ^ 1'b0 ;
  assign n9929 = ( n9773 & n9872 ) | ( n9773 & ~n9928 ) | ( n9872 & ~n9928 ) ;
  assign n9930 = n9915 ^ n9721 ^ 1'b0 ;
  assign n9931 = ( n9721 & n9873 ) | ( n9721 & ~n9930 ) | ( n9873 & ~n9930 ) ;
  assign n9932 = n9915 ^ n9776 ^ 1'b0 ;
  assign n9933 = ( n9776 & n9874 ) | ( n9776 & ~n9932 ) | ( n9874 & ~n9932 ) ;
  assign n9934 = n9915 ^ n9779 ^ 1'b0 ;
  assign n9935 = ( n9779 & n9875 ) | ( n9779 & ~n9934 ) | ( n9875 & ~n9934 ) ;
  assign n9936 = n9915 ^ n9719 ^ 1'b0 ;
  assign n9937 = ( n9719 & n9876 ) | ( n9719 & ~n9936 ) | ( n9876 & ~n9936 ) ;
  assign n9938 = n9915 ^ n9782 ^ 1'b0 ;
  assign n9939 = ( n9782 & n9884 ) | ( n9782 & ~n9938 ) | ( n9884 & ~n9938 ) ;
  assign n9940 = n9915 ^ n9743 ^ 1'b0 ;
  assign n9941 = ( n9743 & n9883 ) | ( n9743 & ~n9940 ) | ( n9883 & ~n9940 ) ;
  assign n9942 = n9915 ^ n9788 ^ 1'b0 ;
  assign n9943 = ( n9788 & n9882 ) | ( n9788 & ~n9942 ) | ( n9882 & ~n9942 ) ;
  assign n9944 = n9915 ^ n9733 ^ 1'b0 ;
  assign n9945 = ( n9733 & n9886 ) | ( n9733 & ~n9944 ) | ( n9886 & ~n9944 ) ;
  assign n9946 = n9915 ^ n9794 ^ 1'b0 ;
  assign n9947 = ( n9794 & n9878 ) | ( n9794 & ~n9946 ) | ( n9878 & ~n9946 ) ;
  assign n9948 = n9915 ^ n9731 ^ 1'b0 ;
  assign n9949 = ( n9731 & n9877 ) | ( n9731 & ~n9948 ) | ( n9877 & ~n9948 ) ;
  assign n9950 = n9915 ^ n9841 ^ 1'b0 ;
  assign n9951 = ( n9714 & n9841 ) | ( n9714 & n9950 ) | ( n9841 & n9950 ) ;
  assign n9952 = n9915 ^ n9839 ^ 1'b0 ;
  assign n9953 = ( n9704 & n9839 ) | ( n9704 & n9952 ) | ( n9839 & n9952 ) ;
  assign n9954 = n9838 & n9914 ;
  assign n9955 = n9910 ^ n9746 ^ x115 ;
  assign n9956 = n9915 ^ n9746 ^ 1'b0 ;
  assign n9957 = ( n9746 & n9955 ) | ( n9746 & ~n9956 ) | ( n9955 & ~n9956 ) ;
  assign n9958 = n9909 ^ n9749 ^ x114 ;
  assign n9959 = n9915 ^ n9749 ^ 1'b0 ;
  assign n9960 = ( n9749 & n9958 ) | ( n9749 & ~n9959 ) | ( n9958 & ~n9959 ) ;
  assign n9961 = n9893 ^ n9755 ^ x98 ;
  assign n9962 = n9915 ^ n9755 ^ 1'b0 ;
  assign n9963 = ( n9755 & n9961 ) | ( n9755 & ~n9962 ) | ( n9961 & ~n9962 ) ;
  assign n9964 = n9892 ^ n9758 ^ x97 ;
  assign n9965 = n9915 ^ n9758 ^ 1'b0 ;
  assign n9966 = ( n9758 & n9964 ) | ( n9758 & ~n9965 ) | ( n9964 & ~n9965 ) ;
  assign n9967 = n9891 ^ n9761 ^ x96 ;
  assign n9968 = n9915 ^ n9761 ^ 1'b0 ;
  assign n9969 = ( n9761 & n9967 ) | ( n9761 & ~n9968 ) | ( n9967 & ~n9968 ) ;
  assign n9970 = n9889 ^ n9720 ^ x95 ;
  assign n9971 = n9915 ^ n9720 ^ 1'b0 ;
  assign n9972 = ( n9720 & n9970 ) | ( n9720 & ~n9971 ) | ( n9970 & ~n9971 ) ;
  assign n9973 = n9879 ^ n9737 ^ x93 ;
  assign n9974 = n9915 ^ n9737 ^ 1'b0 ;
  assign n9975 = ( n9737 & n9973 ) | ( n9737 & ~n9974 ) | ( n9973 & ~n9974 ) ;
  assign n9976 = n9866 ^ n9767 ^ x89 ;
  assign n9977 = n9915 ^ n9767 ^ 1'b0 ;
  assign n9978 = ( n9767 & n9976 ) | ( n9767 & ~n9977 ) | ( n9976 & ~n9977 ) ;
  assign n9979 = n9859 ^ n9718 ^ x84 ;
  assign n9980 = n9915 ^ n9718 ^ 1'b0 ;
  assign n9981 = ( n9718 & n9979 ) | ( n9718 & ~n9980 ) | ( n9979 & ~n9980 ) ;
  assign n9982 = n9854 ^ n9708 ^ x79 ;
  assign n9983 = n9915 ^ n9708 ^ 1'b0 ;
  assign n9984 = ( n9708 & n9982 ) | ( n9708 & ~n9983 ) | ( n9982 & ~n9983 ) ;
  assign n9985 = n9853 ^ n9729 ^ x78 ;
  assign n9986 = n9915 ^ n9729 ^ 1'b0 ;
  assign n9987 = ( n9729 & n9985 ) | ( n9729 & ~n9986 ) | ( n9985 & ~n9986 ) ;
  assign n9988 = n9851 ^ n9732 ^ x76 ;
  assign n9989 = n9915 ^ n9732 ^ 1'b0 ;
  assign n9990 = ( n9732 & n9988 ) | ( n9732 & ~n9989 ) | ( n9988 & ~n9989 ) ;
  assign n9991 = n9850 ^ n9785 ^ x75 ;
  assign n9992 = n9915 ^ n9785 ^ 1'b0 ;
  assign n9993 = ( n9785 & n9991 ) | ( n9785 & ~n9992 ) | ( n9991 & ~n9992 ) ;
  assign n9994 = n9848 ^ n9723 ^ x73 ;
  assign n9995 = n9915 ^ n9723 ^ 1'b0 ;
  assign n9996 = ( n9723 & n9994 ) | ( n9723 & ~n9995 ) | ( n9994 & ~n9995 ) ;
  assign n9997 = n9847 ^ n9728 ^ x72 ;
  assign n9998 = n9915 ^ n9728 ^ 1'b0 ;
  assign n9999 = ( n9728 & n9997 ) | ( n9728 & ~n9998 ) | ( n9997 & ~n9998 ) ;
  assign n10000 = n9846 ^ n9791 ^ x71 ;
  assign n10001 = n9915 ^ n9791 ^ 1'b0 ;
  assign n10002 = ( n9791 & n10000 ) | ( n9791 & ~n10001 ) | ( n10000 & ~n10001 ) ;
  assign n10003 = n9844 ^ n9711 ^ x69 ;
  assign n10004 = n9915 ^ n9711 ^ 1'b0 ;
  assign n10005 = ( n9711 & n10003 ) | ( n9711 & ~n10004 ) | ( n10003 & ~n10004 ) ;
  assign n10006 = n9908 ^ n9797 ^ x113 ;
  assign n10007 = n9915 ^ n9797 ^ 1'b0 ;
  assign n10008 = ( n9797 & n10006 ) | ( n9797 & ~n10007 ) | ( n10006 & ~n10007 ) ;
  assign n10009 = n9915 ^ n9804 ^ 1'b0 ;
  assign n10010 = n9906 ^ n9801 ^ x111 ;
  assign n10011 = n9915 ^ n9801 ^ 1'b0 ;
  assign n10012 = ( n9801 & n10010 ) | ( n9801 & ~n10011 ) | ( n10010 & ~n10011 ) ;
  assign n10013 = n9905 ^ n9806 ^ x110 ;
  assign n10014 = n9915 ^ n9806 ^ 1'b0 ;
  assign n10015 = ( n9806 & n10013 ) | ( n9806 & ~n10014 ) | ( n10013 & ~n10014 ) ;
  assign n10016 = n9904 ^ n9809 ^ x109 ;
  assign n10017 = n9915 ^ n9809 ^ 1'b0 ;
  assign n10018 = ( n9809 & n10016 ) | ( n9809 & ~n10017 ) | ( n10016 & ~n10017 ) ;
  assign n10019 = n9903 ^ n9812 ^ x108 ;
  assign n10020 = n9915 ^ n9812 ^ 1'b0 ;
  assign n10021 = n9907 ^ n9804 ^ x112 ;
  assign n10022 = ( n9804 & ~n10009 ) | ( n9804 & n10021 ) | ( ~n10009 & n10021 ) ;
  assign n10023 = ( n9812 & n10019 ) | ( n9812 & ~n10020 ) | ( n10019 & ~n10020 ) ;
  assign n10024 = n9902 ^ n9815 ^ x107 ;
  assign n10025 = n9915 ^ n9815 ^ 1'b0 ;
  assign n10026 = ( n9815 & n10024 ) | ( n9815 & ~n10025 ) | ( n10024 & ~n10025 ) ;
  assign n10027 = n9901 ^ n9818 ^ x106 ;
  assign n10028 = n9915 ^ n9818 ^ 1'b0 ;
  assign n10029 = ( n9818 & n10027 ) | ( n9818 & ~n10028 ) | ( n10027 & ~n10028 ) ;
  assign n10030 = n9900 ^ n9821 ^ x105 ;
  assign n10031 = n9915 ^ n9821 ^ 1'b0 ;
  assign n10032 = ( n9821 & n10030 ) | ( n9821 & ~n10031 ) | ( n10030 & ~n10031 ) ;
  assign n10033 = n9899 ^ n9824 ^ x104 ;
  assign n10034 = n9915 ^ n9824 ^ 1'b0 ;
  assign n10035 = ( n9824 & n10033 ) | ( n9824 & ~n10034 ) | ( n10033 & ~n10034 ) ;
  assign n10036 = n9898 ^ n9827 ^ x103 ;
  assign n10037 = n9915 ^ n9827 ^ 1'b0 ;
  assign n10038 = ( n9827 & n10036 ) | ( n9827 & ~n10037 ) | ( n10036 & ~n10037 ) ;
  assign n10039 = n9897 ^ n9830 ^ x102 ;
  assign n10040 = n9915 ^ n9830 ^ 1'b0 ;
  assign n10041 = ( n9830 & n10039 ) | ( n9830 & ~n10040 ) | ( n10039 & ~n10040 ) ;
  assign n10042 = n9896 ^ n9833 ^ x101 ;
  assign n10043 = n9915 ^ n9833 ^ 1'b0 ;
  assign n10044 = ( n9833 & n10042 ) | ( n9833 & ~n10043 ) | ( n10042 & ~n10043 ) ;
  assign n10045 = n9895 ^ n9836 ^ x100 ;
  assign n10046 = n9915 ^ n9836 ^ 1'b0 ;
  assign n10047 = ( n9836 & n10045 ) | ( n9836 & ~n10046 ) | ( n10045 & ~n10046 ) ;
  assign n10048 = n9894 ^ n9752 ^ x99 ;
  assign n10049 = n9915 ^ n9752 ^ 1'b0 ;
  assign n10050 = ( n9752 & n10048 ) | ( n9752 & ~n10049 ) | ( n10048 & ~n10049 ) ;
  assign n10051 = x64 & n9915 ;
  assign n10052 = n10051 ^ x64 ^ x11 ;
  assign n10053 = n322 | n9954 ;
  assign n10054 = n10052 ^ n7180 ^ x65 ;
  assign n10055 = ( x65 & n7180 ) | ( x65 & n10054 ) | ( n7180 & n10054 ) ;
  assign n10056 = n10055 ^ n9953 ^ x66 ;
  assign n10057 = ( x66 & n10055 ) | ( x66 & n10056 ) | ( n10055 & n10056 ) ;
  assign n10058 = ( x67 & ~n9951 ) | ( x67 & n10057 ) | ( ~n9951 & n10057 ) ;
  assign n10059 = ( x68 & ~n9949 ) | ( x68 & n10058 ) | ( ~n9949 & n10058 ) ;
  assign n10060 = ( x69 & ~n9947 ) | ( x69 & n10059 ) | ( ~n9947 & n10059 ) ;
  assign n10061 = ( x70 & ~n10005 ) | ( x70 & n10060 ) | ( ~n10005 & n10060 ) ;
  assign n10062 = ( x71 & ~n9945 ) | ( x71 & n10061 ) | ( ~n9945 & n10061 ) ;
  assign n10063 = ( x72 & ~n10002 ) | ( x72 & n10062 ) | ( ~n10002 & n10062 ) ;
  assign n10064 = ( x73 & ~n9999 ) | ( x73 & n10063 ) | ( ~n9999 & n10063 ) ;
  assign n10065 = ( x74 & ~n9996 ) | ( x74 & n10064 ) | ( ~n9996 & n10064 ) ;
  assign n10066 = ( x75 & ~n9943 ) | ( x75 & n10065 ) | ( ~n9943 & n10065 ) ;
  assign n10067 = ( x76 & ~n9993 ) | ( x76 & n10066 ) | ( ~n9993 & n10066 ) ;
  assign n10068 = ( x77 & ~n9990 ) | ( x77 & n10067 ) | ( ~n9990 & n10067 ) ;
  assign n10069 = ( x78 & ~n9941 ) | ( x78 & n10068 ) | ( ~n9941 & n10068 ) ;
  assign n10070 = ( x79 & ~n9987 ) | ( x79 & n10069 ) | ( ~n9987 & n10069 ) ;
  assign n10071 = n10070 ^ n9984 ^ x80 ;
  assign n10072 = n10068 ^ n9941 ^ x78 ;
  assign n10073 = n10067 ^ n9990 ^ x77 ;
  assign n10074 = n10064 ^ n9996 ^ x74 ;
  assign n10075 = n10063 ^ n9999 ^ x73 ;
  assign n10076 = n10057 ^ n9951 ^ x67 ;
  assign n10077 = ( x80 & ~n9984 ) | ( x80 & n10070 ) | ( ~n9984 & n10070 ) ;
  assign n10078 = ( x81 & ~n9939 ) | ( x81 & n10077 ) | ( ~n9939 & n10077 ) ;
  assign n10079 = n10078 ^ n9937 ^ x82 ;
  assign n10080 = n10077 ^ n9939 ^ x81 ;
  assign n10081 = ( x82 & ~n9937 ) | ( x82 & n10078 ) | ( ~n9937 & n10078 ) ;
  assign n10082 = ( x83 & ~n9935 ) | ( x83 & n10081 ) | ( ~n9935 & n10081 ) ;
  assign n10083 = n171 & n10053 ;
  assign n10084 = n10081 ^ n9935 ^ x83 ;
  assign n10085 = ( x84 & ~n9933 ) | ( x84 & n10082 ) | ( ~n9933 & n10082 ) ;
  assign n10086 = ( x85 & ~n9981 ) | ( x85 & n10085 ) | ( ~n9981 & n10085 ) ;
  assign n10087 = n10085 ^ n9981 ^ x85 ;
  assign n10088 = ( x86 & ~n9931 ) | ( x86 & n10086 ) | ( ~n9931 & n10086 ) ;
  assign n10089 = n10088 ^ n9929 ^ x87 ;
  assign n10090 = ( x87 & ~n9929 ) | ( x87 & n10088 ) | ( ~n9929 & n10088 ) ;
  assign n10091 = ( x88 & ~n9927 ) | ( x88 & n10090 ) | ( ~n9927 & n10090 ) ;
  assign n10092 = n10091 ^ n9925 ^ x89 ;
  assign n10093 = ( x89 & ~n9925 ) | ( x89 & n10091 ) | ( ~n9925 & n10091 ) ;
  assign n10094 = ( x90 & ~n9978 ) | ( x90 & n10093 ) | ( ~n9978 & n10093 ) ;
  assign n10095 = ( x91 & ~n9923 ) | ( x91 & n10094 ) | ( ~n9923 & n10094 ) ;
  assign n10096 = ( x92 & ~n9921 ) | ( x92 & n10095 ) | ( ~n9921 & n10095 ) ;
  assign n10097 = ( x93 & ~n9919 ) | ( x93 & n10096 ) | ( ~n9919 & n10096 ) ;
  assign n10098 = ( x94 & ~n9975 ) | ( x94 & n10097 ) | ( ~n9975 & n10097 ) ;
  assign n10099 = n10098 ^ n9917 ^ x95 ;
  assign n10100 = ( x95 & ~n9917 ) | ( x95 & n10098 ) | ( ~n9917 & n10098 ) ;
  assign n10101 = ( x96 & ~n9972 ) | ( x96 & n10100 ) | ( ~n9972 & n10100 ) ;
  assign n10102 = n10100 ^ n9972 ^ x96 ;
  assign n10103 = ( x97 & ~n9969 ) | ( x97 & n10101 ) | ( ~n9969 & n10101 ) ;
  assign n10104 = n10101 ^ n9969 ^ x97 ;
  assign n10105 = n10094 ^ n9923 ^ x91 ;
  assign n10106 = n10096 ^ n9919 ^ x93 ;
  assign n10107 = ( x98 & ~n9966 ) | ( x98 & n10103 ) | ( ~n9966 & n10103 ) ;
  assign n10108 = ( x99 & ~n9963 ) | ( x99 & n10107 ) | ( ~n9963 & n10107 ) ;
  assign n10109 = ( x100 & ~n10050 ) | ( x100 & n10108 ) | ( ~n10050 & n10108 ) ;
  assign n10110 = ( x101 & ~n10047 ) | ( x101 & n10109 ) | ( ~n10047 & n10109 ) ;
  assign n10111 = ( x102 & ~n10044 ) | ( x102 & n10110 ) | ( ~n10044 & n10110 ) ;
  assign n10112 = ( x103 & ~n10041 ) | ( x103 & n10111 ) | ( ~n10041 & n10111 ) ;
  assign n10113 = ( x104 & ~n10038 ) | ( x104 & n10112 ) | ( ~n10038 & n10112 ) ;
  assign n10114 = ( x105 & ~n10035 ) | ( x105 & n10113 ) | ( ~n10035 & n10113 ) ;
  assign n10115 = ( x106 & ~n10032 ) | ( x106 & n10114 ) | ( ~n10032 & n10114 ) ;
  assign n10116 = ( x107 & ~n10029 ) | ( x107 & n10115 ) | ( ~n10029 & n10115 ) ;
  assign n10117 = ( x108 & ~n10026 ) | ( x108 & n10116 ) | ( ~n10026 & n10116 ) ;
  assign n10118 = ( x109 & ~n10023 ) | ( x109 & n10117 ) | ( ~n10023 & n10117 ) ;
  assign n10119 = ( x110 & ~n10018 ) | ( x110 & n10118 ) | ( ~n10018 & n10118 ) ;
  assign n10120 = ( x111 & ~n10015 ) | ( x111 & n10119 ) | ( ~n10015 & n10119 ) ;
  assign n10121 = ( x112 & ~n10012 ) | ( x112 & n10120 ) | ( ~n10012 & n10120 ) ;
  assign n10122 = ( x113 & ~n10022 ) | ( x113 & n10121 ) | ( ~n10022 & n10121 ) ;
  assign n10123 = ( x114 & ~n10008 ) | ( x114 & n10122 ) | ( ~n10008 & n10122 ) ;
  assign n10124 = ( x115 & ~n9960 ) | ( x115 & n10123 ) | ( ~n9960 & n10123 ) ;
  assign n10125 = ( x116 & ~n9957 ) | ( x116 & n10124 ) | ( ~n9957 & n10124 ) ;
  assign n10126 = ( x117 & n10053 ) | ( x117 & ~n10125 ) | ( n10053 & ~n10125 ) ;
  assign n10127 = ( x117 & n9954 ) | ( x117 & n10125 ) | ( n9954 & n10125 ) ;
  assign n10128 = ( n7187 & n10126 ) | ( n7187 & ~n10127 ) | ( n10126 & ~n10127 ) ;
  assign n10129 = n10125 | n10128 ;
  assign n10130 = ( ~n10053 & n10083 ) | ( ~n10053 & n10129 ) | ( n10083 & n10129 ) ;
  assign n10131 = n10108 ^ n10050 ^ x100 ;
  assign n10132 = n10130 ^ n10050 ^ 1'b0 ;
  assign n10133 = ( n10050 & n10131 ) | ( n10050 & ~n10132 ) | ( n10131 & ~n10132 ) ;
  assign n10134 = n10130 ^ n9969 ^ 1'b0 ;
  assign n10135 = ( n9969 & n10104 ) | ( n9969 & ~n10134 ) | ( n10104 & ~n10134 ) ;
  assign n10136 = n10130 ^ n9972 ^ 1'b0 ;
  assign n10137 = ( n9972 & n10102 ) | ( n9972 & ~n10136 ) | ( n10102 & ~n10136 ) ;
  assign n10138 = n10130 ^ n9917 ^ 1'b0 ;
  assign n10139 = ( n9917 & n10099 ) | ( n9917 & ~n10138 ) | ( n10099 & ~n10138 ) ;
  assign n10140 = n10130 ^ n9919 ^ 1'b0 ;
  assign n10141 = ( n9919 & n10106 ) | ( n9919 & ~n10140 ) | ( n10106 & ~n10140 ) ;
  assign n10142 = n10130 ^ n9923 ^ 1'b0 ;
  assign n10143 = ( n9923 & n10105 ) | ( n9923 & ~n10142 ) | ( n10105 & ~n10142 ) ;
  assign n10144 = n10130 ^ n9925 ^ 1'b0 ;
  assign n10145 = ( n9925 & n10092 ) | ( n9925 & ~n10144 ) | ( n10092 & ~n10144 ) ;
  assign n10146 = n10130 ^ n9929 ^ 1'b0 ;
  assign n10147 = ( n9929 & n10089 ) | ( n9929 & ~n10146 ) | ( n10089 & ~n10146 ) ;
  assign n10148 = n10130 ^ n9981 ^ 1'b0 ;
  assign n10149 = ( n9981 & n10087 ) | ( n9981 & ~n10148 ) | ( n10087 & ~n10148 ) ;
  assign n10150 = n10130 ^ n9935 ^ 1'b0 ;
  assign n10151 = ( n9935 & n10084 ) | ( n9935 & ~n10150 ) | ( n10084 & ~n10150 ) ;
  assign n10152 = n10130 ^ n9937 ^ 1'b0 ;
  assign n10153 = ( n9937 & n10079 ) | ( n9937 & ~n10152 ) | ( n10079 & ~n10152 ) ;
  assign n10154 = n10130 ^ n9939 ^ 1'b0 ;
  assign n10155 = ( n9939 & n10080 ) | ( n9939 & ~n10154 ) | ( n10080 & ~n10154 ) ;
  assign n10156 = n10130 ^ n9984 ^ 1'b0 ;
  assign n10157 = ( n9984 & n10071 ) | ( n9984 & ~n10156 ) | ( n10071 & ~n10156 ) ;
  assign n10158 = n10130 ^ n9941 ^ 1'b0 ;
  assign n10159 = ( n9941 & n10072 ) | ( n9941 & ~n10158 ) | ( n10072 & ~n10158 ) ;
  assign n10160 = n10130 ^ n9990 ^ 1'b0 ;
  assign n10161 = ( n9990 & n10073 ) | ( n9990 & ~n10160 ) | ( n10073 & ~n10160 ) ;
  assign n10162 = n10130 ^ n9996 ^ 1'b0 ;
  assign n10163 = ( n9996 & n10074 ) | ( n9996 & ~n10162 ) | ( n10074 & ~n10162 ) ;
  assign n10164 = n10130 ^ n9999 ^ 1'b0 ;
  assign n10165 = ( n9999 & n10075 ) | ( n9999 & ~n10164 ) | ( n10075 & ~n10164 ) ;
  assign n10166 = n10130 ^ n9951 ^ 1'b0 ;
  assign n10167 = ( n9951 & n10076 ) | ( n9951 & ~n10166 ) | ( n10076 & ~n10166 ) ;
  assign n10168 = n10130 ^ n10056 ^ 1'b0 ;
  assign n10169 = ( n9953 & n10056 ) | ( n9953 & n10168 ) | ( n10056 & n10168 ) ;
  assign n10170 = n10083 & ~n10129 ;
  assign n10171 = ( n322 & n10083 ) | ( n322 & ~n10170 ) | ( n10083 & ~n10170 ) ;
  assign n10172 = n10124 ^ n9957 ^ x116 ;
  assign n10173 = n10130 ^ n9957 ^ 1'b0 ;
  assign n10174 = ( n9957 & n10172 ) | ( n9957 & ~n10173 ) | ( n10172 & ~n10173 ) ;
  assign n10175 = n10123 ^ n9960 ^ x115 ;
  assign n10176 = n10130 ^ n9960 ^ 1'b0 ;
  assign n10177 = ( n9960 & n10175 ) | ( n9960 & ~n10176 ) | ( n10175 & ~n10176 ) ;
  assign n10178 = n10122 ^ n10008 ^ x114 ;
  assign n10179 = n10130 ^ n10008 ^ 1'b0 ;
  assign n10180 = ( n10008 & n10178 ) | ( n10008 & ~n10179 ) | ( n10178 & ~n10179 ) ;
  assign n10181 = n10103 ^ n9966 ^ x98 ;
  assign n10182 = n10130 ^ n9966 ^ 1'b0 ;
  assign n10183 = ( n9966 & n10181 ) | ( n9966 & ~n10182 ) | ( n10181 & ~n10182 ) ;
  assign n10184 = n10097 ^ n9975 ^ x94 ;
  assign n10185 = n10130 ^ n9975 ^ 1'b0 ;
  assign n10186 = ( n9975 & n10184 ) | ( n9975 & ~n10185 ) | ( n10184 & ~n10185 ) ;
  assign n10187 = n10095 ^ n9921 ^ x92 ;
  assign n10188 = n10130 ^ n9921 ^ 1'b0 ;
  assign n10189 = ( n9921 & n10187 ) | ( n9921 & ~n10188 ) | ( n10187 & ~n10188 ) ;
  assign n10190 = n10093 ^ n9978 ^ x90 ;
  assign n10191 = n10130 ^ n9978 ^ 1'b0 ;
  assign n10192 = ( n9978 & n10190 ) | ( n9978 & ~n10191 ) | ( n10190 & ~n10191 ) ;
  assign n10193 = n10090 ^ n9927 ^ x88 ;
  assign n10194 = n10130 ^ n9927 ^ 1'b0 ;
  assign n10195 = ( n9927 & n10193 ) | ( n9927 & ~n10194 ) | ( n10193 & ~n10194 ) ;
  assign n10196 = n10086 ^ n9931 ^ x86 ;
  assign n10197 = n10130 ^ n9931 ^ 1'b0 ;
  assign n10198 = ( n9931 & n10196 ) | ( n9931 & ~n10197 ) | ( n10196 & ~n10197 ) ;
  assign n10199 = n10082 ^ n9933 ^ x84 ;
  assign n10200 = n10130 ^ n9933 ^ 1'b0 ;
  assign n10201 = ( n9933 & n10199 ) | ( n9933 & ~n10200 ) | ( n10199 & ~n10200 ) ;
  assign n10202 = n10069 ^ n9987 ^ x79 ;
  assign n10203 = n10130 ^ n9987 ^ 1'b0 ;
  assign n10204 = ( n9987 & n10202 ) | ( n9987 & ~n10203 ) | ( n10202 & ~n10203 ) ;
  assign n10205 = n10066 ^ n9993 ^ x76 ;
  assign n10206 = n10130 ^ n9993 ^ 1'b0 ;
  assign n10207 = ( n9993 & n10205 ) | ( n9993 & ~n10206 ) | ( n10205 & ~n10206 ) ;
  assign n10208 = n10065 ^ n9943 ^ x75 ;
  assign n10209 = n10130 ^ n9943 ^ 1'b0 ;
  assign n10210 = ( n9943 & n10208 ) | ( n9943 & ~n10209 ) | ( n10208 & ~n10209 ) ;
  assign n10211 = n10062 ^ n10002 ^ x72 ;
  assign n10212 = n10130 ^ n10002 ^ 1'b0 ;
  assign n10213 = ( n10002 & n10211 ) | ( n10002 & ~n10212 ) | ( n10211 & ~n10212 ) ;
  assign n10214 = n10061 ^ n9945 ^ x71 ;
  assign n10215 = n10130 ^ n9945 ^ 1'b0 ;
  assign n10216 = ( n9945 & n10214 ) | ( n9945 & ~n10215 ) | ( n10214 & ~n10215 ) ;
  assign n10217 = n10060 ^ n10005 ^ x70 ;
  assign n10218 = n10130 ^ n10005 ^ 1'b0 ;
  assign n10219 = ( n10005 & n10217 ) | ( n10005 & ~n10218 ) | ( n10217 & ~n10218 ) ;
  assign n10220 = n10059 ^ n9947 ^ x69 ;
  assign n10221 = n10130 ^ n9947 ^ 1'b0 ;
  assign n10222 = ( n9947 & n10220 ) | ( n9947 & ~n10221 ) | ( n10220 & ~n10221 ) ;
  assign n10223 = n10058 ^ n9949 ^ x68 ;
  assign n10224 = n10130 ^ n9949 ^ 1'b0 ;
  assign n10225 = ( n9949 & n10223 ) | ( n9949 & ~n10224 ) | ( n10223 & ~n10224 ) ;
  assign n10226 = n10121 ^ n10022 ^ x113 ;
  assign n10227 = n10130 ^ n10022 ^ 1'b0 ;
  assign n10228 = ( n10022 & n10226 ) | ( n10022 & ~n10227 ) | ( n10226 & ~n10227 ) ;
  assign n10229 = n10120 ^ n10012 ^ x112 ;
  assign n10230 = n10130 ^ n10012 ^ 1'b0 ;
  assign n10231 = ( n10012 & n10229 ) | ( n10012 & ~n10230 ) | ( n10229 & ~n10230 ) ;
  assign n10232 = n10119 ^ n10015 ^ x111 ;
  assign n10233 = n10130 ^ n10015 ^ 1'b0 ;
  assign n10234 = ( n10015 & n10232 ) | ( n10015 & ~n10233 ) | ( n10232 & ~n10233 ) ;
  assign n10235 = n10118 ^ n10018 ^ x110 ;
  assign n10236 = n10130 ^ n10018 ^ 1'b0 ;
  assign n10237 = ( n10018 & n10235 ) | ( n10018 & ~n10236 ) | ( n10235 & ~n10236 ) ;
  assign n10238 = n10117 ^ n10023 ^ x109 ;
  assign n10239 = n10130 ^ n10023 ^ 1'b0 ;
  assign n10240 = ( n10023 & n10238 ) | ( n10023 & ~n10239 ) | ( n10238 & ~n10239 ) ;
  assign n10241 = n10116 ^ n10026 ^ x108 ;
  assign n10242 = n10130 ^ n10026 ^ 1'b0 ;
  assign n10243 = ( n10026 & n10241 ) | ( n10026 & ~n10242 ) | ( n10241 & ~n10242 ) ;
  assign n10244 = n10115 ^ n10029 ^ x107 ;
  assign n10245 = n10130 ^ n10029 ^ 1'b0 ;
  assign n10246 = ( n10029 & n10244 ) | ( n10029 & ~n10245 ) | ( n10244 & ~n10245 ) ;
  assign n10247 = n10114 ^ n10032 ^ x106 ;
  assign n10248 = n10130 ^ n10032 ^ 1'b0 ;
  assign n10249 = ( n10032 & n10247 ) | ( n10032 & ~n10248 ) | ( n10247 & ~n10248 ) ;
  assign n10250 = n10113 ^ n10035 ^ x105 ;
  assign n10251 = n10130 ^ n10035 ^ 1'b0 ;
  assign n10252 = ( n10035 & n10250 ) | ( n10035 & ~n10251 ) | ( n10250 & ~n10251 ) ;
  assign n10253 = n10112 ^ n10038 ^ x104 ;
  assign n10254 = n10130 ^ n10038 ^ 1'b0 ;
  assign n10255 = ( n10038 & n10253 ) | ( n10038 & ~n10254 ) | ( n10253 & ~n10254 ) ;
  assign n10256 = n10111 ^ n10041 ^ x103 ;
  assign n10257 = n10130 ^ n10041 ^ 1'b0 ;
  assign n10258 = ( n10041 & n10256 ) | ( n10041 & ~n10257 ) | ( n10256 & ~n10257 ) ;
  assign n10259 = n10110 ^ n10044 ^ x102 ;
  assign n10260 = n10130 ^ n10044 ^ 1'b0 ;
  assign n10261 = ( n10044 & n10259 ) | ( n10044 & ~n10260 ) | ( n10259 & ~n10260 ) ;
  assign n10262 = n10109 ^ n10047 ^ x101 ;
  assign n10263 = n10130 ^ n10047 ^ 1'b0 ;
  assign n10264 = ( n10047 & n10262 ) | ( n10047 & ~n10263 ) | ( n10262 & ~n10263 ) ;
  assign n10265 = n10107 ^ n9963 ^ x99 ;
  assign n10266 = n10130 ^ n9963 ^ 1'b0 ;
  assign n10267 = ( n9963 & n10265 ) | ( n9963 & ~n10266 ) | ( n10265 & ~n10266 ) ;
  assign n10268 = x64 & n10130 ;
  assign n10269 = n10268 ^ x64 ^ x10 ;
  assign n10270 = n10130 ^ n10054 ^ 1'b0 ;
  assign n10271 = ( n10052 & n10054 ) | ( n10052 & n10270 ) | ( n10054 & n10270 ) ;
  assign n10272 = n10269 ^ n7381 ^ x65 ;
  assign n10273 = ( x65 & n7381 ) | ( x65 & n10272 ) | ( n7381 & n10272 ) ;
  assign n10274 = n10273 ^ n10271 ^ x66 ;
  assign n10275 = ( x66 & n10273 ) | ( x66 & n10274 ) | ( n10273 & n10274 ) ;
  assign n10276 = ( x67 & ~n10169 ) | ( x67 & n10275 ) | ( ~n10169 & n10275 ) ;
  assign n10277 = ( x68 & ~n10167 ) | ( x68 & n10276 ) | ( ~n10167 & n10276 ) ;
  assign n10278 = ( x69 & ~n10225 ) | ( x69 & n10277 ) | ( ~n10225 & n10277 ) ;
  assign n10279 = ( x70 & ~n10222 ) | ( x70 & n10278 ) | ( ~n10222 & n10278 ) ;
  assign n10280 = ( x71 & ~n10219 ) | ( x71 & n10279 ) | ( ~n10219 & n10279 ) ;
  assign n10281 = ( x72 & ~n10216 ) | ( x72 & n10280 ) | ( ~n10216 & n10280 ) ;
  assign n10282 = ( x73 & ~n10213 ) | ( x73 & n10281 ) | ( ~n10213 & n10281 ) ;
  assign n10283 = ( x74 & ~n10165 ) | ( x74 & n10282 ) | ( ~n10165 & n10282 ) ;
  assign n10284 = ( x75 & ~n10163 ) | ( x75 & n10283 ) | ( ~n10163 & n10283 ) ;
  assign n10285 = ( x76 & ~n10210 ) | ( x76 & n10284 ) | ( ~n10210 & n10284 ) ;
  assign n10286 = ( x77 & ~n10207 ) | ( x77 & n10285 ) | ( ~n10207 & n10285 ) ;
  assign n10287 = ( x78 & ~n10161 ) | ( x78 & n10286 ) | ( ~n10161 & n10286 ) ;
  assign n10288 = ( x79 & ~n10159 ) | ( x79 & n10287 ) | ( ~n10159 & n10287 ) ;
  assign n10289 = ( x80 & ~n10204 ) | ( x80 & n10288 ) | ( ~n10204 & n10288 ) ;
  assign n10290 = ( x81 & ~n10157 ) | ( x81 & n10289 ) | ( ~n10157 & n10289 ) ;
  assign n10291 = ( x82 & ~n10155 ) | ( x82 & n10290 ) | ( ~n10155 & n10290 ) ;
  assign n10292 = ( x83 & ~n10153 ) | ( x83 & n10291 ) | ( ~n10153 & n10291 ) ;
  assign n10293 = ( x84 & ~n10151 ) | ( x84 & n10292 ) | ( ~n10151 & n10292 ) ;
  assign n10294 = ( x85 & ~n10201 ) | ( x85 & n10293 ) | ( ~n10201 & n10293 ) ;
  assign n10295 = ( x86 & ~n10149 ) | ( x86 & n10294 ) | ( ~n10149 & n10294 ) ;
  assign n10296 = ( x87 & ~n10198 ) | ( x87 & n10295 ) | ( ~n10198 & n10295 ) ;
  assign n10297 = ( x88 & ~n10147 ) | ( x88 & n10296 ) | ( ~n10147 & n10296 ) ;
  assign n10298 = ( x89 & ~n10195 ) | ( x89 & n10297 ) | ( ~n10195 & n10297 ) ;
  assign n10299 = ( x90 & ~n10145 ) | ( x90 & n10298 ) | ( ~n10145 & n10298 ) ;
  assign n10300 = ( x91 & ~n10192 ) | ( x91 & n10299 ) | ( ~n10192 & n10299 ) ;
  assign n10301 = ( x92 & ~n10143 ) | ( x92 & n10300 ) | ( ~n10143 & n10300 ) ;
  assign n10302 = ( x93 & ~n10189 ) | ( x93 & n10301 ) | ( ~n10189 & n10301 ) ;
  assign n10303 = ( x94 & ~n10141 ) | ( x94 & n10302 ) | ( ~n10141 & n10302 ) ;
  assign n10304 = ( x95 & ~n10186 ) | ( x95 & n10303 ) | ( ~n10186 & n10303 ) ;
  assign n10305 = ( x96 & ~n10139 ) | ( x96 & n10304 ) | ( ~n10139 & n10304 ) ;
  assign n10306 = ( x97 & ~n10137 ) | ( x97 & n10305 ) | ( ~n10137 & n10305 ) ;
  assign n10307 = n10295 ^ n10198 ^ x87 ;
  assign n10308 = ( x98 & ~n10135 ) | ( x98 & n10306 ) | ( ~n10135 & n10306 ) ;
  assign n10309 = ( x99 & ~n10183 ) | ( x99 & n10308 ) | ( ~n10183 & n10308 ) ;
  assign n10310 = ( x100 & ~n10267 ) | ( x100 & n10309 ) | ( ~n10267 & n10309 ) ;
  assign n10311 = n10299 ^ n10192 ^ x91 ;
  assign n10312 = n10300 ^ n10143 ^ x92 ;
  assign n10313 = n10301 ^ n10189 ^ x93 ;
  assign n10314 = ( x101 & ~n10133 ) | ( x101 & n10310 ) | ( ~n10133 & n10310 ) ;
  assign n10315 = n10293 ^ n10201 ^ x85 ;
  assign n10316 = n10304 ^ n10139 ^ x96 ;
  assign n10317 = n10309 ^ n10267 ^ x100 ;
  assign n10318 = n10289 ^ n10157 ^ x81 ;
  assign n10319 = n10287 ^ n10159 ^ x79 ;
  assign n10320 = n10292 ^ n10151 ^ x84 ;
  assign n10321 = n10283 ^ n10163 ^ x75 ;
  assign n10322 = n10280 ^ n10216 ^ x72 ;
  assign n10323 = ( x102 & ~n10264 ) | ( x102 & n10314 ) | ( ~n10264 & n10314 ) ;
  assign n10324 = ( x103 & ~n10261 ) | ( x103 & n10323 ) | ( ~n10261 & n10323 ) ;
  assign n10325 = ( x104 & ~n10258 ) | ( x104 & n10324 ) | ( ~n10258 & n10324 ) ;
  assign n10326 = ( x105 & ~n10255 ) | ( x105 & n10325 ) | ( ~n10255 & n10325 ) ;
  assign n10327 = ( x106 & ~n10252 ) | ( x106 & n10326 ) | ( ~n10252 & n10326 ) ;
  assign n10328 = ( x107 & ~n10249 ) | ( x107 & n10327 ) | ( ~n10249 & n10327 ) ;
  assign n10329 = ( x108 & ~n10246 ) | ( x108 & n10328 ) | ( ~n10246 & n10328 ) ;
  assign n10330 = ( x109 & ~n10243 ) | ( x109 & n10329 ) | ( ~n10243 & n10329 ) ;
  assign n10331 = ( x110 & ~n10240 ) | ( x110 & n10330 ) | ( ~n10240 & n10330 ) ;
  assign n10332 = ( x111 & ~n10237 ) | ( x111 & n10331 ) | ( ~n10237 & n10331 ) ;
  assign n10333 = ( x112 & ~n10234 ) | ( x112 & n10332 ) | ( ~n10234 & n10332 ) ;
  assign n10334 = ( x113 & ~n10231 ) | ( x113 & n10333 ) | ( ~n10231 & n10333 ) ;
  assign n10335 = ( x114 & ~n10228 ) | ( x114 & n10334 ) | ( ~n10228 & n10334 ) ;
  assign n10336 = ( x115 & ~n10180 ) | ( x115 & n10335 ) | ( ~n10180 & n10335 ) ;
  assign n10337 = ( x116 & ~n10177 ) | ( x116 & n10336 ) | ( ~n10177 & n10336 ) ;
  assign n10338 = ( x117 & ~n10174 ) | ( x117 & n10337 ) | ( ~n10174 & n10337 ) ;
  assign n10339 = ( x118 & ~n10171 ) | ( x118 & n10338 ) | ( ~n10171 & n10338 ) ;
  assign n10340 = n10324 ^ n10258 ^ x104 ;
  assign n10341 = n7632 | n10339 ;
  assign n10342 = ( x9 & ~n10339 ) | ( x9 & n10341 ) | ( ~n10339 & n10341 ) ;
  assign n10343 = ~n7631 & n10342 ;
  assign n10344 = ( n10341 & n10342 ) | ( n10341 & n10343 ) | ( n10342 & n10343 ) ;
  assign n10345 = n1296 | n10339 ;
  assign n10346 = n10345 ^ n10143 ^ 1'b0 ;
  assign n10347 = n10345 ^ n10272 ^ 1'b0 ;
  assign n10348 = ( n10269 & n10272 ) | ( n10269 & n10347 ) | ( n10272 & n10347 ) ;
  assign n10349 = n10345 ^ n10151 ^ 1'b0 ;
  assign n10350 = ( n10151 & n10320 ) | ( n10151 & ~n10349 ) | ( n10320 & ~n10349 ) ;
  assign n10351 = n10345 ^ n10198 ^ 1'b0 ;
  assign n10352 = n10325 ^ n10255 ^ x105 ;
  assign n10353 = n10323 ^ n10261 ^ x103 ;
  assign n10354 = n10345 ^ n10139 ^ 1'b0 ;
  assign n10355 = n10345 ^ n10163 ^ 1'b0 ;
  assign n10356 = ( n10143 & n10312 ) | ( n10143 & ~n10346 ) | ( n10312 & ~n10346 ) ;
  assign n10357 = n10345 ^ n10261 ^ 1'b0 ;
  assign n10358 = n10345 ^ n10192 ^ 1'b0 ;
  assign n10359 = ( n10192 & n10311 ) | ( n10192 & ~n10358 ) | ( n10311 & ~n10358 ) ;
  assign n10360 = n10345 ^ n10258 ^ 1'b0 ;
  assign n10361 = n10345 ^ n10189 ^ 1'b0 ;
  assign n10362 = ( n10163 & n10321 ) | ( n10163 & ~n10355 ) | ( n10321 & ~n10355 ) ;
  assign n10363 = n10345 ^ n10157 ^ 1'b0 ;
  assign n10364 = n10345 ^ n10255 ^ 1'b0 ;
  assign n10365 = ( n10261 & n10353 ) | ( n10261 & ~n10357 ) | ( n10353 & ~n10357 ) ;
  assign n10366 = n10345 ^ n10216 ^ 1'b0 ;
  assign n10367 = ( n10216 & n10322 ) | ( n10216 & ~n10366 ) | ( n10322 & ~n10366 ) ;
  assign n10368 = ( n10189 & n10313 ) | ( n10189 & ~n10361 ) | ( n10313 & ~n10361 ) ;
  assign n10369 = ( n10258 & n10340 ) | ( n10258 & ~n10360 ) | ( n10340 & ~n10360 ) ;
  assign n10370 = ( n10255 & n10352 ) | ( n10255 & ~n10364 ) | ( n10352 & ~n10364 ) ;
  assign n10371 = n10345 ^ n10267 ^ 1'b0 ;
  assign n10372 = n10345 ^ n10274 ^ 1'b0 ;
  assign n10373 = n10345 ^ n10201 ^ 1'b0 ;
  assign n10374 = n10345 ^ n10159 ^ 1'b0 ;
  assign n10375 = n10314 ^ n10264 ^ x102 ;
  assign n10376 = ( n10159 & n10319 ) | ( n10159 & ~n10374 ) | ( n10319 & ~n10374 ) ;
  assign n10377 = ( n10201 & n10315 ) | ( n10201 & ~n10373 ) | ( n10315 & ~n10373 ) ;
  assign n10378 = ( n10139 & n10316 ) | ( n10139 & ~n10354 ) | ( n10316 & ~n10354 ) ;
  assign n10379 = ( n10198 & n10307 ) | ( n10198 & ~n10351 ) | ( n10307 & ~n10351 ) ;
  assign n10380 = n10345 ^ n10264 ^ 1'b0 ;
  assign n10381 = ( n10264 & n10375 ) | ( n10264 & ~n10380 ) | ( n10375 & ~n10380 ) ;
  assign n10382 = ( n10271 & n10274 ) | ( n10271 & n10372 ) | ( n10274 & n10372 ) ;
  assign n10383 = ( n10157 & n10318 ) | ( n10157 & ~n10363 ) | ( n10318 & ~n10363 ) ;
  assign n10384 = ( n10267 & n10317 ) | ( n10267 & ~n10371 ) | ( n10317 & ~n10371 ) ;
  assign n10385 = n10337 ^ n10174 ^ x117 ;
  assign n10386 = n10345 ^ n10174 ^ 1'b0 ;
  assign n10387 = ( n10174 & n10385 ) | ( n10174 & ~n10386 ) | ( n10385 & ~n10386 ) ;
  assign n10388 = n10336 ^ n10177 ^ x116 ;
  assign n10389 = n10345 ^ n10177 ^ 1'b0 ;
  assign n10390 = ( n10177 & n10388 ) | ( n10177 & ~n10389 ) | ( n10388 & ~n10389 ) ;
  assign n10391 = n10302 ^ n10141 ^ x94 ;
  assign n10392 = n10345 ^ n10141 ^ 1'b0 ;
  assign n10393 = ( n10141 & n10391 ) | ( n10141 & ~n10392 ) | ( n10391 & ~n10392 ) ;
  assign n10394 = n10298 ^ n10145 ^ x90 ;
  assign n10395 = n10345 ^ n10145 ^ 1'b0 ;
  assign n10396 = ( n10145 & n10394 ) | ( n10145 & ~n10395 ) | ( n10394 & ~n10395 ) ;
  assign n10397 = n10297 ^ n10195 ^ x89 ;
  assign n10398 = n10345 ^ n10195 ^ 1'b0 ;
  assign n10399 = ( n10195 & n10397 ) | ( n10195 & ~n10398 ) | ( n10397 & ~n10398 ) ;
  assign n10400 = n10296 ^ n10147 ^ x88 ;
  assign n10401 = n10345 ^ n10147 ^ 1'b0 ;
  assign n10402 = ( n10147 & n10400 ) | ( n10147 & ~n10401 ) | ( n10400 & ~n10401 ) ;
  assign n10403 = n10294 ^ n10149 ^ x86 ;
  assign n10404 = n10345 ^ n10149 ^ 1'b0 ;
  assign n10405 = ( n10149 & n10403 ) | ( n10149 & ~n10404 ) | ( n10403 & ~n10404 ) ;
  assign n10406 = n10291 ^ n10153 ^ x83 ;
  assign n10407 = n10345 ^ n10153 ^ 1'b0 ;
  assign n10408 = ( n10153 & n10406 ) | ( n10153 & ~n10407 ) | ( n10406 & ~n10407 ) ;
  assign n10409 = n10290 ^ n10155 ^ x82 ;
  assign n10410 = n10345 ^ n10155 ^ 1'b0 ;
  assign n10411 = ( n10155 & n10409 ) | ( n10155 & ~n10410 ) | ( n10409 & ~n10410 ) ;
  assign n10412 = n10288 ^ n10204 ^ x80 ;
  assign n10413 = n10345 ^ n10204 ^ 1'b0 ;
  assign n10414 = ( n10204 & n10412 ) | ( n10204 & ~n10413 ) | ( n10412 & ~n10413 ) ;
  assign n10415 = n10286 ^ n10161 ^ x78 ;
  assign n10416 = n10345 ^ n10161 ^ 1'b0 ;
  assign n10417 = ( n10161 & n10415 ) | ( n10161 & ~n10416 ) | ( n10415 & ~n10416 ) ;
  assign n10418 = n10285 ^ n10207 ^ x77 ;
  assign n10419 = n10345 ^ n10207 ^ 1'b0 ;
  assign n10420 = ( n10207 & n10418 ) | ( n10207 & ~n10419 ) | ( n10418 & ~n10419 ) ;
  assign n10421 = n10284 ^ n10210 ^ x76 ;
  assign n10422 = n10345 ^ n10210 ^ 1'b0 ;
  assign n10423 = ( n10210 & n10421 ) | ( n10210 & ~n10422 ) | ( n10421 & ~n10422 ) ;
  assign n10424 = n10282 ^ n10165 ^ x74 ;
  assign n10425 = n10345 ^ n10165 ^ 1'b0 ;
  assign n10426 = ( n10165 & n10424 ) | ( n10165 & ~n10425 ) | ( n10424 & ~n10425 ) ;
  assign n10427 = n10281 ^ n10213 ^ x73 ;
  assign n10428 = n10345 ^ n10213 ^ 1'b0 ;
  assign n10429 = ( n10213 & n10427 ) | ( n10213 & ~n10428 ) | ( n10427 & ~n10428 ) ;
  assign n10430 = n10279 ^ n10219 ^ x71 ;
  assign n10431 = n10345 ^ n10219 ^ 1'b0 ;
  assign n10432 = ( n10219 & n10430 ) | ( n10219 & ~n10431 ) | ( n10430 & ~n10431 ) ;
  assign n10433 = n10276 ^ n10167 ^ x68 ;
  assign n10434 = n10345 ^ n10167 ^ 1'b0 ;
  assign n10435 = ( n10167 & n10433 ) | ( n10167 & ~n10434 ) | ( n10433 & ~n10434 ) ;
  assign n10436 = n10335 ^ n10180 ^ x115 ;
  assign n10437 = n10345 ^ n10180 ^ 1'b0 ;
  assign n10438 = ( n10180 & n10436 ) | ( n10180 & ~n10437 ) | ( n10436 & ~n10437 ) ;
  assign n10439 = n10334 ^ n10228 ^ x114 ;
  assign n10440 = n10345 ^ n10228 ^ 1'b0 ;
  assign n10441 = ( n10228 & n10439 ) | ( n10228 & ~n10440 ) | ( n10439 & ~n10440 ) ;
  assign n10442 = n10333 ^ n10231 ^ x113 ;
  assign n10443 = n10345 ^ n10231 ^ 1'b0 ;
  assign n10444 = ( n10231 & n10442 ) | ( n10231 & ~n10443 ) | ( n10442 & ~n10443 ) ;
  assign n10445 = n10332 ^ n10234 ^ x112 ;
  assign n10446 = n10345 ^ n10234 ^ 1'b0 ;
  assign n10447 = ( n10234 & n10445 ) | ( n10234 & ~n10446 ) | ( n10445 & ~n10446 ) ;
  assign n10448 = n10331 ^ n10237 ^ x111 ;
  assign n10449 = n10345 ^ n10237 ^ 1'b0 ;
  assign n10450 = ( n10237 & n10448 ) | ( n10237 & ~n10449 ) | ( n10448 & ~n10449 ) ;
  assign n10451 = n10330 ^ n10240 ^ x110 ;
  assign n10452 = n10345 ^ n10240 ^ 1'b0 ;
  assign n10453 = ( n10240 & n10451 ) | ( n10240 & ~n10452 ) | ( n10451 & ~n10452 ) ;
  assign n10454 = n10329 ^ n10243 ^ x109 ;
  assign n10455 = n10345 ^ n10243 ^ 1'b0 ;
  assign n10456 = ( n10243 & n10454 ) | ( n10243 & ~n10455 ) | ( n10454 & ~n10455 ) ;
  assign n10457 = n10328 ^ n10246 ^ x108 ;
  assign n10458 = n10345 ^ n10246 ^ 1'b0 ;
  assign n10459 = ( n10246 & n10457 ) | ( n10246 & ~n10458 ) | ( n10457 & ~n10458 ) ;
  assign n10460 = n10327 ^ n10249 ^ x107 ;
  assign n10461 = n10345 ^ n10249 ^ 1'b0 ;
  assign n10462 = ( n10249 & n10460 ) | ( n10249 & ~n10461 ) | ( n10460 & ~n10461 ) ;
  assign n10463 = n10326 ^ n10252 ^ x106 ;
  assign n10464 = n10345 ^ n10252 ^ 1'b0 ;
  assign n10465 = ( n10252 & n10463 ) | ( n10252 & ~n10464 ) | ( n10463 & ~n10464 ) ;
  assign n10466 = n10310 ^ n10133 ^ x101 ;
  assign n10467 = n10345 ^ n10133 ^ 1'b0 ;
  assign n10468 = ( n10133 & n10466 ) | ( n10133 & ~n10467 ) | ( n10466 & ~n10467 ) ;
  assign n10469 = n10308 ^ n10183 ^ x99 ;
  assign n10470 = n10345 ^ n10183 ^ 1'b0 ;
  assign n10471 = ( n10183 & n10469 ) | ( n10183 & ~n10470 ) | ( n10469 & ~n10470 ) ;
  assign n10472 = n10306 ^ n10135 ^ x98 ;
  assign n10473 = n10345 ^ n10135 ^ 1'b0 ;
  assign n10474 = ( n10135 & n10472 ) | ( n10135 & ~n10473 ) | ( n10472 & ~n10473 ) ;
  assign n10475 = n10305 ^ n10137 ^ x97 ;
  assign n10476 = n10345 ^ n10137 ^ 1'b0 ;
  assign n10477 = ( n10137 & n10475 ) | ( n10137 & ~n10476 ) | ( n10475 & ~n10476 ) ;
  assign n10478 = n10303 ^ n10186 ^ x95 ;
  assign n10479 = n10345 ^ n10186 ^ 1'b0 ;
  assign n10480 = ( n10186 & n10478 ) | ( n10186 & ~n10479 ) | ( n10478 & ~n10479 ) ;
  assign n10481 = n10278 ^ n10222 ^ x70 ;
  assign n10482 = n10345 ^ n10222 ^ 1'b0 ;
  assign n10483 = ( n10222 & n10481 ) | ( n10222 & ~n10482 ) | ( n10481 & ~n10482 ) ;
  assign n10484 = n10277 ^ n10225 ^ x69 ;
  assign n10485 = n10345 ^ n10225 ^ 1'b0 ;
  assign n10486 = n10275 ^ n10169 ^ x67 ;
  assign n10487 = n10345 ^ n10169 ^ 1'b0 ;
  assign n10488 = ( n10169 & n10486 ) | ( n10169 & ~n10487 ) | ( n10486 & ~n10487 ) ;
  assign n10489 = n10344 ^ n7629 ^ x65 ;
  assign n10490 = n10171 & n10345 ;
  assign n10491 = n322 | n10490 ;
  assign n10492 = n1296 & n10491 ;
  assign n10493 = n1296 & n10171 ;
  assign n10494 = ( n10225 & n10484 ) | ( n10225 & ~n10485 ) | ( n10484 & ~n10485 ) ;
  assign n10495 = ( x65 & n7629 ) | ( x65 & n10489 ) | ( n7629 & n10489 ) ;
  assign n10496 = n10495 ^ n10348 ^ x66 ;
  assign n10497 = ( x66 & n10495 ) | ( x66 & n10496 ) | ( n10495 & n10496 ) ;
  assign n10498 = ( x67 & ~n10382 ) | ( x67 & n10497 ) | ( ~n10382 & n10497 ) ;
  assign n10499 = ( x68 & ~n10488 ) | ( x68 & n10498 ) | ( ~n10488 & n10498 ) ;
  assign n10500 = ( x69 & ~n10435 ) | ( x69 & n10499 ) | ( ~n10435 & n10499 ) ;
  assign n10501 = ( x70 & ~n10494 ) | ( x70 & n10500 ) | ( ~n10494 & n10500 ) ;
  assign n10502 = ( x71 & ~n10483 ) | ( x71 & n10501 ) | ( ~n10483 & n10501 ) ;
  assign n10503 = ( x72 & ~n10432 ) | ( x72 & n10502 ) | ( ~n10432 & n10502 ) ;
  assign n10504 = ( x73 & ~n10367 ) | ( x73 & n10503 ) | ( ~n10367 & n10503 ) ;
  assign n10505 = ( x74 & ~n10429 ) | ( x74 & n10504 ) | ( ~n10429 & n10504 ) ;
  assign n10506 = ( x75 & ~n10426 ) | ( x75 & n10505 ) | ( ~n10426 & n10505 ) ;
  assign n10507 = n10501 ^ n10483 ^ x71 ;
  assign n10508 = ( x76 & ~n10362 ) | ( x76 & n10506 ) | ( ~n10362 & n10506 ) ;
  assign n10509 = ( x77 & ~n10423 ) | ( x77 & n10508 ) | ( ~n10423 & n10508 ) ;
  assign n10510 = ( x78 & ~n10420 ) | ( x78 & n10509 ) | ( ~n10420 & n10509 ) ;
  assign n10511 = n10505 ^ n10426 ^ x75 ;
  assign n10512 = n10506 ^ n10362 ^ x76 ;
  assign n10513 = ( x79 & ~n10417 ) | ( x79 & n10510 ) | ( ~n10417 & n10510 ) ;
  assign n10514 = ( x80 & ~n10376 ) | ( x80 & n10513 ) | ( ~n10376 & n10513 ) ;
  assign n10515 = ( x81 & ~n10414 ) | ( x81 & n10514 ) | ( ~n10414 & n10514 ) ;
  assign n10516 = ( x82 & ~n10383 ) | ( x82 & n10515 ) | ( ~n10383 & n10515 ) ;
  assign n10517 = ( x83 & ~n10411 ) | ( x83 & n10516 ) | ( ~n10411 & n10516 ) ;
  assign n10518 = ( x84 & ~n10408 ) | ( x84 & n10517 ) | ( ~n10408 & n10517 ) ;
  assign n10519 = ( x85 & ~n10350 ) | ( x85 & n10518 ) | ( ~n10350 & n10518 ) ;
  assign n10520 = ( x86 & ~n10377 ) | ( x86 & n10519 ) | ( ~n10377 & n10519 ) ;
  assign n10521 = ( x87 & ~n10405 ) | ( x87 & n10520 ) | ( ~n10405 & n10520 ) ;
  assign n10522 = ( x88 & ~n10379 ) | ( x88 & n10521 ) | ( ~n10379 & n10521 ) ;
  assign n10523 = ( x89 & ~n10402 ) | ( x89 & n10522 ) | ( ~n10402 & n10522 ) ;
  assign n10524 = ( x90 & ~n10399 ) | ( x90 & n10523 ) | ( ~n10399 & n10523 ) ;
  assign n10525 = ( x91 & ~n10396 ) | ( x91 & n10524 ) | ( ~n10396 & n10524 ) ;
  assign n10526 = ( x92 & ~n10359 ) | ( x92 & n10525 ) | ( ~n10359 & n10525 ) ;
  assign n10527 = ( ~x119 & n163 ) | ( ~x119 & n10491 ) | ( n163 & n10491 ) ;
  assign n10528 = n10498 ^ n10488 ^ x68 ;
  assign n10529 = ( x119 & n163 ) | ( x119 & ~n10490 ) | ( n163 & ~n10490 ) ;
  assign n10530 = ( x93 & ~n10356 ) | ( x93 & n10526 ) | ( ~n10356 & n10526 ) ;
  assign n10531 = ( x94 & ~n10368 ) | ( x94 & n10530 ) | ( ~n10368 & n10530 ) ;
  assign n10532 = ( x95 & ~n10393 ) | ( x95 & n10531 ) | ( ~n10393 & n10531 ) ;
  assign n10533 = ( x96 & ~n10480 ) | ( x96 & n10532 ) | ( ~n10480 & n10532 ) ;
  assign n10534 = ( x97 & ~n10378 ) | ( x97 & n10533 ) | ( ~n10378 & n10533 ) ;
  assign n10535 = ( x98 & ~n10477 ) | ( x98 & n10534 ) | ( ~n10477 & n10534 ) ;
  assign n10536 = ( x99 & ~n10474 ) | ( x99 & n10535 ) | ( ~n10474 & n10535 ) ;
  assign n10537 = ( x100 & ~n10471 ) | ( x100 & n10536 ) | ( ~n10471 & n10536 ) ;
  assign n10538 = ( x101 & ~n10384 ) | ( x101 & n10537 ) | ( ~n10384 & n10537 ) ;
  assign n10539 = ( x102 & ~n10468 ) | ( x102 & n10538 ) | ( ~n10468 & n10538 ) ;
  assign n10540 = ( x103 & ~n10381 ) | ( x103 & n10539 ) | ( ~n10381 & n10539 ) ;
  assign n10541 = ( x104 & ~n10365 ) | ( x104 & n10540 ) | ( ~n10365 & n10540 ) ;
  assign n10542 = ( x105 & ~n10369 ) | ( x105 & n10541 ) | ( ~n10369 & n10541 ) ;
  assign n10543 = ( x106 & ~n10370 ) | ( x106 & n10542 ) | ( ~n10370 & n10542 ) ;
  assign n10544 = ( x107 & ~n10465 ) | ( x107 & n10543 ) | ( ~n10465 & n10543 ) ;
  assign n10545 = ( x108 & ~n10462 ) | ( x108 & n10544 ) | ( ~n10462 & n10544 ) ;
  assign n10546 = ( x109 & ~n10459 ) | ( x109 & n10545 ) | ( ~n10459 & n10545 ) ;
  assign n10547 = ( x110 & ~n10456 ) | ( x110 & n10546 ) | ( ~n10456 & n10546 ) ;
  assign n10548 = ( x111 & ~n10453 ) | ( x111 & n10547 ) | ( ~n10453 & n10547 ) ;
  assign n10549 = ( x112 & ~n10450 ) | ( x112 & n10548 ) | ( ~n10450 & n10548 ) ;
  assign n10550 = ( x113 & ~n10447 ) | ( x113 & n10549 ) | ( ~n10447 & n10549 ) ;
  assign n10551 = ( x114 & ~n10444 ) | ( x114 & n10550 ) | ( ~n10444 & n10550 ) ;
  assign n10552 = ( x115 & ~n10441 ) | ( x115 & n10551 ) | ( ~n10441 & n10551 ) ;
  assign n10553 = ( x116 & ~n10438 ) | ( x116 & n10552 ) | ( ~n10438 & n10552 ) ;
  assign n10554 = ( x117 & ~n10390 ) | ( x117 & n10553 ) | ( ~n10390 & n10553 ) ;
  assign n10555 = ( x118 & ~n10387 ) | ( x118 & n10554 ) | ( ~n10387 & n10554 ) ;
  assign n10556 = ( n10527 & n10529 ) | ( n10527 & ~n10555 ) | ( n10529 & ~n10555 ) ;
  assign n10557 = n10555 | n10556 ;
  assign n10558 = ( ~n10491 & n10492 ) | ( ~n10491 & n10557 ) | ( n10492 & n10557 ) ;
  assign n10559 = n10553 ^ n10390 ^ x117 ;
  assign n10560 = n10558 ^ n10390 ^ 1'b0 ;
  assign n10561 = ( n10390 & n10559 ) | ( n10390 & ~n10560 ) | ( n10559 & ~n10560 ) ;
  assign n10562 = n10552 ^ n10438 ^ x116 ;
  assign n10563 = n10558 ^ n10438 ^ 1'b0 ;
  assign n10564 = ( n10438 & n10562 ) | ( n10438 & ~n10563 ) | ( n10562 & ~n10563 ) ;
  assign n10565 = n10551 ^ n10441 ^ x115 ;
  assign n10566 = n10558 ^ n10441 ^ 1'b0 ;
  assign n10567 = ( n10441 & n10565 ) | ( n10441 & ~n10566 ) | ( n10565 & ~n10566 ) ;
  assign n10568 = n10550 ^ n10444 ^ x114 ;
  assign n10569 = n10558 ^ n10444 ^ 1'b0 ;
  assign n10570 = ( n10444 & n10568 ) | ( n10444 & ~n10569 ) | ( n10568 & ~n10569 ) ;
  assign n10571 = n10549 ^ n10447 ^ x113 ;
  assign n10572 = n10548 ^ n10450 ^ x112 ;
  assign n10573 = n10558 ^ n10450 ^ 1'b0 ;
  assign n10574 = ( n10450 & n10572 ) | ( n10450 & ~n10573 ) | ( n10572 & ~n10573 ) ;
  assign n10575 = n10547 ^ n10453 ^ x111 ;
  assign n10576 = n10558 ^ n10453 ^ 1'b0 ;
  assign n10577 = ( n10453 & n10575 ) | ( n10453 & ~n10576 ) | ( n10575 & ~n10576 ) ;
  assign n10578 = n10545 ^ n10459 ^ x109 ;
  assign n10579 = n10558 ^ n10459 ^ 1'b0 ;
  assign n10580 = ( n10459 & n10578 ) | ( n10459 & ~n10579 ) | ( n10578 & ~n10579 ) ;
  assign n10581 = n10558 ^ n10447 ^ 1'b0 ;
  assign n10582 = ( n10447 & n10571 ) | ( n10447 & ~n10581 ) | ( n10571 & ~n10581 ) ;
  assign n10583 = n10558 ^ n10362 ^ 1'b0 ;
  assign n10584 = ( n10362 & n10512 ) | ( n10362 & ~n10583 ) | ( n10512 & ~n10583 ) ;
  assign n10585 = n10558 ^ n10426 ^ 1'b0 ;
  assign n10586 = ( n10426 & n10511 ) | ( n10426 & ~n10585 ) | ( n10511 & ~n10585 ) ;
  assign n10587 = n10558 ^ n10483 ^ 1'b0 ;
  assign n10588 = ( n10483 & n10507 ) | ( n10483 & ~n10587 ) | ( n10507 & ~n10587 ) ;
  assign n10589 = n10558 ^ n10488 ^ 1'b0 ;
  assign n10590 = ( n10488 & n10528 ) | ( n10488 & ~n10589 ) | ( n10528 & ~n10589 ) ;
  assign n10591 = n10558 ^ n10496 ^ 1'b0 ;
  assign n10592 = ( n10348 & n10496 ) | ( n10348 & n10591 ) | ( n10496 & n10591 ) ;
  assign n10593 = n10493 & n10557 ;
  assign n10594 = n10544 ^ n10462 ^ x108 ;
  assign n10595 = n10558 ^ n10462 ^ 1'b0 ;
  assign n10596 = ( n10462 & n10594 ) | ( n10462 & ~n10595 ) | ( n10594 & ~n10595 ) ;
  assign n10597 = n10543 ^ n10465 ^ x107 ;
  assign n10598 = n10558 ^ n10465 ^ 1'b0 ;
  assign n10599 = ( n10465 & n10597 ) | ( n10465 & ~n10598 ) | ( n10597 & ~n10598 ) ;
  assign n10600 = n10522 ^ n10402 ^ x89 ;
  assign n10601 = n10558 ^ n10402 ^ 1'b0 ;
  assign n10602 = ( n10402 & n10600 ) | ( n10402 & ~n10601 ) | ( n10600 & ~n10601 ) ;
  assign n10603 = n10521 ^ n10379 ^ x88 ;
  assign n10604 = n10558 ^ n10379 ^ 1'b0 ;
  assign n10605 = ( n10379 & n10603 ) | ( n10379 & ~n10604 ) | ( n10603 & ~n10604 ) ;
  assign n10606 = n10520 ^ n10405 ^ x87 ;
  assign n10607 = n10558 ^ n10405 ^ 1'b0 ;
  assign n10608 = ( n10405 & n10606 ) | ( n10405 & ~n10607 ) | ( n10606 & ~n10607 ) ;
  assign n10609 = n10519 ^ n10377 ^ x86 ;
  assign n10610 = n10558 ^ n10377 ^ 1'b0 ;
  assign n10611 = ( n10377 & n10609 ) | ( n10377 & ~n10610 ) | ( n10609 & ~n10610 ) ;
  assign n10612 = n10517 ^ n10408 ^ x84 ;
  assign n10613 = n10558 ^ n10408 ^ 1'b0 ;
  assign n10614 = ( n10408 & n10612 ) | ( n10408 & ~n10613 ) | ( n10612 & ~n10613 ) ;
  assign n10615 = n10516 ^ n10411 ^ x83 ;
  assign n10616 = n10558 ^ n10411 ^ 1'b0 ;
  assign n10617 = ( n10411 & n10615 ) | ( n10411 & ~n10616 ) | ( n10615 & ~n10616 ) ;
  assign n10618 = n10515 ^ n10383 ^ x82 ;
  assign n10619 = n10558 ^ n10383 ^ 1'b0 ;
  assign n10620 = ( n10383 & n10618 ) | ( n10383 & ~n10619 ) | ( n10618 & ~n10619 ) ;
  assign n10621 = n10513 ^ n10376 ^ x80 ;
  assign n10622 = n10558 ^ n10376 ^ 1'b0 ;
  assign n10623 = ( n10376 & n10621 ) | ( n10376 & ~n10622 ) | ( n10621 & ~n10622 ) ;
  assign n10624 = n10510 ^ n10417 ^ x79 ;
  assign n10625 = n10558 ^ n10417 ^ 1'b0 ;
  assign n10626 = ( n10417 & n10624 ) | ( n10417 & ~n10625 ) | ( n10624 & ~n10625 ) ;
  assign n10627 = n10509 ^ n10420 ^ x78 ;
  assign n10628 = n10558 ^ n10420 ^ 1'b0 ;
  assign n10629 = ( n10420 & n10627 ) | ( n10420 & ~n10628 ) | ( n10627 & ~n10628 ) ;
  assign n10630 = n10508 ^ n10423 ^ x77 ;
  assign n10631 = n10558 ^ n10423 ^ 1'b0 ;
  assign n10632 = ( n10423 & n10630 ) | ( n10423 & ~n10631 ) | ( n10630 & ~n10631 ) ;
  assign n10633 = n10504 ^ n10429 ^ x74 ;
  assign n10634 = n10558 ^ n10429 ^ 1'b0 ;
  assign n10635 = ( n10429 & n10633 ) | ( n10429 & ~n10634 ) | ( n10633 & ~n10634 ) ;
  assign n10636 = n10502 ^ n10432 ^ x72 ;
  assign n10637 = n10558 ^ n10432 ^ 1'b0 ;
  assign n10638 = ( n10432 & n10636 ) | ( n10432 & ~n10637 ) | ( n10636 & ~n10637 ) ;
  assign n10639 = n10500 ^ n10494 ^ x70 ;
  assign n10640 = n10558 ^ n10494 ^ 1'b0 ;
  assign n10641 = ( n10494 & n10639 ) | ( n10494 & ~n10640 ) | ( n10639 & ~n10640 ) ;
  assign n10642 = n10497 ^ n10382 ^ x67 ;
  assign n10643 = n10558 ^ n10382 ^ 1'b0 ;
  assign n10644 = ( n10382 & n10642 ) | ( n10382 & ~n10643 ) | ( n10642 & ~n10643 ) ;
  assign n10645 = n10542 ^ n10370 ^ x106 ;
  assign n10646 = n10558 ^ n10370 ^ 1'b0 ;
  assign n10647 = ( n10370 & n10645 ) | ( n10370 & ~n10646 ) | ( n10645 & ~n10646 ) ;
  assign n10648 = n10541 ^ n10369 ^ x105 ;
  assign n10649 = n10558 ^ n10369 ^ 1'b0 ;
  assign n10650 = ( n10369 & n10648 ) | ( n10369 & ~n10649 ) | ( n10648 & ~n10649 ) ;
  assign n10651 = n10540 ^ n10365 ^ x104 ;
  assign n10652 = n10558 ^ n10365 ^ 1'b0 ;
  assign n10653 = ( n10365 & n10651 ) | ( n10365 & ~n10652 ) | ( n10651 & ~n10652 ) ;
  assign n10654 = n10539 ^ n10381 ^ x103 ;
  assign n10655 = n10558 ^ n10381 ^ 1'b0 ;
  assign n10656 = ( n10381 & n10654 ) | ( n10381 & ~n10655 ) | ( n10654 & ~n10655 ) ;
  assign n10657 = n10538 ^ n10468 ^ x102 ;
  assign n10658 = n10558 ^ n10468 ^ 1'b0 ;
  assign n10659 = ( n10468 & n10657 ) | ( n10468 & ~n10658 ) | ( n10657 & ~n10658 ) ;
  assign n10660 = n10537 ^ n10384 ^ x101 ;
  assign n10661 = n10558 ^ n10384 ^ 1'b0 ;
  assign n10662 = ( n10384 & n10660 ) | ( n10384 & ~n10661 ) | ( n10660 & ~n10661 ) ;
  assign n10663 = n10535 ^ n10474 ^ x99 ;
  assign n10664 = n10558 ^ n10474 ^ 1'b0 ;
  assign n10665 = ( n10474 & n10663 ) | ( n10474 & ~n10664 ) | ( n10663 & ~n10664 ) ;
  assign n10666 = n10534 ^ n10477 ^ x98 ;
  assign n10667 = n10558 ^ n10477 ^ 1'b0 ;
  assign n10668 = ( n10477 & n10666 ) | ( n10477 & ~n10667 ) | ( n10666 & ~n10667 ) ;
  assign n10669 = n10533 ^ n10378 ^ x97 ;
  assign n10670 = n10558 ^ n10378 ^ 1'b0 ;
  assign n10671 = ( n10378 & n10669 ) | ( n10378 & ~n10670 ) | ( n10669 & ~n10670 ) ;
  assign n10672 = n10532 ^ n10480 ^ x96 ;
  assign n10673 = n10558 ^ n10480 ^ 1'b0 ;
  assign n10674 = ( n10480 & n10672 ) | ( n10480 & ~n10673 ) | ( n10672 & ~n10673 ) ;
  assign n10675 = n10531 ^ n10393 ^ x95 ;
  assign n10676 = n10558 ^ n10393 ^ 1'b0 ;
  assign n10677 = ( n10393 & n10675 ) | ( n10393 & ~n10676 ) | ( n10675 & ~n10676 ) ;
  assign n10678 = n10530 ^ n10368 ^ x94 ;
  assign n10679 = n10558 ^ n10368 ^ 1'b0 ;
  assign n10680 = ( n10368 & n10678 ) | ( n10368 & ~n10679 ) | ( n10678 & ~n10679 ) ;
  assign n10681 = n10526 ^ n10356 ^ x93 ;
  assign n10682 = n10558 ^ n10356 ^ 1'b0 ;
  assign n10683 = ( n10356 & n10681 ) | ( n10356 & ~n10682 ) | ( n10681 & ~n10682 ) ;
  assign n10684 = n10524 ^ n10396 ^ x91 ;
  assign n10685 = n10558 ^ n10396 ^ 1'b0 ;
  assign n10686 = ( n10396 & n10684 ) | ( n10396 & ~n10685 ) | ( n10684 & ~n10685 ) ;
  assign n10687 = n10523 ^ n10399 ^ x90 ;
  assign n10688 = n10558 ^ n10399 ^ 1'b0 ;
  assign n10689 = ( n10399 & n10687 ) | ( n10399 & ~n10688 ) | ( n10687 & ~n10688 ) ;
  assign n10690 = n10546 ^ n10456 ^ x110 ;
  assign n10691 = n10558 ^ n10387 ^ 1'b0 ;
  assign n10692 = n10536 ^ n10471 ^ x100 ;
  assign n10693 = n10558 ^ n10367 ^ 1'b0 ;
  assign n10694 = n10558 ^ n10456 ^ 1'b0 ;
  assign n10695 = n10558 ^ n10414 ^ 1'b0 ;
  assign n10696 = n10518 ^ n10350 ^ x85 ;
  assign n10697 = n10499 ^ n10435 ^ x69 ;
  assign n10698 = n10558 ^ n10489 ^ 1'b0 ;
  assign n10699 = n10558 ^ n10435 ^ 1'b0 ;
  assign n10700 = ( n10344 & n10489 ) | ( n10344 & n10698 ) | ( n10489 & n10698 ) ;
  assign n10701 = n10558 ^ n10350 ^ 1'b0 ;
  assign n10702 = x64 & n10558 ;
  assign n10703 = n10702 ^ x64 ^ x8 ;
  assign n10704 = n10703 ^ n7863 ^ x65 ;
  assign n10705 = ( n10435 & n10697 ) | ( n10435 & ~n10699 ) | ( n10697 & ~n10699 ) ;
  assign n10706 = ( x65 & n7863 ) | ( x65 & n10704 ) | ( n7863 & n10704 ) ;
  assign n10707 = n10706 ^ n10700 ^ x66 ;
  assign n10708 = ( x66 & n10706 ) | ( x66 & n10707 ) | ( n10706 & n10707 ) ;
  assign n10709 = ( x67 & ~n10592 ) | ( x67 & n10708 ) | ( ~n10592 & n10708 ) ;
  assign n10710 = ( x68 & ~n10644 ) | ( x68 & n10709 ) | ( ~n10644 & n10709 ) ;
  assign n10711 = ( x69 & ~n10590 ) | ( x69 & n10710 ) | ( ~n10590 & n10710 ) ;
  assign n10712 = ( x70 & ~n10705 ) | ( x70 & n10711 ) | ( ~n10705 & n10711 ) ;
  assign n10713 = ( x71 & ~n10641 ) | ( x71 & n10712 ) | ( ~n10641 & n10712 ) ;
  assign n10714 = n10713 ^ n10588 ^ x72 ;
  assign n10715 = ( n10456 & n10690 ) | ( n10456 & ~n10694 ) | ( n10690 & ~n10694 ) ;
  assign n10716 = n10554 ^ n10387 ^ x118 ;
  assign n10717 = n10503 ^ n10367 ^ x73 ;
  assign n10718 = n10514 ^ n10414 ^ x81 ;
  assign n10719 = n322 | n10593 ;
  assign n10720 = ( x72 & ~n10588 ) | ( x72 & n10713 ) | ( ~n10588 & n10713 ) ;
  assign n10721 = ( x73 & ~n10638 ) | ( x73 & n10720 ) | ( ~n10638 & n10720 ) ;
  assign n10722 = ( n10367 & ~n10693 ) | ( n10367 & n10717 ) | ( ~n10693 & n10717 ) ;
  assign n10723 = ( x74 & n10721 ) | ( x74 & ~n10722 ) | ( n10721 & ~n10722 ) ;
  assign n10724 = ( x75 & ~n10635 ) | ( x75 & n10723 ) | ( ~n10635 & n10723 ) ;
  assign n10725 = ( x76 & ~n10586 ) | ( x76 & n10724 ) | ( ~n10586 & n10724 ) ;
  assign n10726 = ( x77 & ~n10584 ) | ( x77 & n10725 ) | ( ~n10584 & n10725 ) ;
  assign n10727 = n10726 ^ n10632 ^ x78 ;
  assign n10728 = n10725 ^ n10584 ^ x77 ;
  assign n10729 = ( x78 & ~n10632 ) | ( x78 & n10726 ) | ( ~n10632 & n10726 ) ;
  assign n10730 = n10729 ^ n10629 ^ x79 ;
  assign n10731 = ( x79 & ~n10629 ) | ( x79 & n10729 ) | ( ~n10629 & n10729 ) ;
  assign n10732 = ( x80 & ~n10626 ) | ( x80 & n10731 ) | ( ~n10626 & n10731 ) ;
  assign n10733 = ( x81 & ~n10623 ) | ( x81 & n10732 ) | ( ~n10623 & n10732 ) ;
  assign n10734 = n10732 ^ n10623 ^ x81 ;
  assign n10735 = ( n10350 & n10696 ) | ( n10350 & ~n10701 ) | ( n10696 & ~n10701 ) ;
  assign n10736 = ( n10414 & ~n10695 ) | ( n10414 & n10718 ) | ( ~n10695 & n10718 ) ;
  assign n10737 = n10558 ^ n10471 ^ 1'b0 ;
  assign n10738 = n10736 ^ n10733 ^ x82 ;
  assign n10739 = ( n10471 & n10692 ) | ( n10471 & ~n10737 ) | ( n10692 & ~n10737 ) ;
  assign n10740 = ( x82 & n10733 ) | ( x82 & ~n10736 ) | ( n10733 & ~n10736 ) ;
  assign n10741 = n10740 ^ n10620 ^ x83 ;
  assign n10742 = ( x83 & ~n10620 ) | ( x83 & n10740 ) | ( ~n10620 & n10740 ) ;
  assign n10743 = ( x84 & ~n10617 ) | ( x84 & n10742 ) | ( ~n10617 & n10742 ) ;
  assign n10744 = ( x85 & ~n10614 ) | ( x85 & n10743 ) | ( ~n10614 & n10743 ) ;
  assign n10745 = ( x86 & ~n10735 ) | ( x86 & n10744 ) | ( ~n10735 & n10744 ) ;
  assign n10746 = n10745 ^ n10611 ^ x87 ;
  assign n10747 = ( x87 & ~n10611 ) | ( x87 & n10745 ) | ( ~n10611 & n10745 ) ;
  assign n10748 = ( x88 & ~n10608 ) | ( x88 & n10747 ) | ( ~n10608 & n10747 ) ;
  assign n10749 = n10748 ^ n10605 ^ x89 ;
  assign n10750 = ( x89 & ~n10605 ) | ( x89 & n10748 ) | ( ~n10605 & n10748 ) ;
  assign n10751 = ( x90 & ~n10602 ) | ( x90 & n10750 ) | ( ~n10602 & n10750 ) ;
  assign n10752 = ( x91 & ~n10689 ) | ( x91 & n10751 ) | ( ~n10689 & n10751 ) ;
  assign n10753 = ( x92 & ~n10686 ) | ( x92 & n10752 ) | ( ~n10686 & n10752 ) ;
  assign n10754 = n10751 ^ n10689 ^ x91 ;
  assign n10755 = n10558 ^ n10359 ^ 1'b0 ;
  assign n10756 = n10525 ^ n10359 ^ x92 ;
  assign n10757 = ( x120 & n156 ) | ( x120 & ~n10593 ) | ( n156 & ~n10593 ) ;
  assign n10758 = ( n10387 & ~n10691 ) | ( n10387 & n10716 ) | ( ~n10691 & n10716 ) ;
  assign n10759 = ( n10359 & ~n10755 ) | ( n10359 & n10756 ) | ( ~n10755 & n10756 ) ;
  assign n10760 = ( x93 & n10753 ) | ( x93 & ~n10759 ) | ( n10753 & ~n10759 ) ;
  assign n10761 = ( x94 & ~n10683 ) | ( x94 & n10760 ) | ( ~n10683 & n10760 ) ;
  assign n10762 = ( x95 & ~n10680 ) | ( x95 & n10761 ) | ( ~n10680 & n10761 ) ;
  assign n10763 = n10762 ^ n10677 ^ x96 ;
  assign n10764 = n163 & n10719 ;
  assign n10765 = ( ~x120 & n156 ) | ( ~x120 & n10719 ) | ( n156 & n10719 ) ;
  assign n10766 = n10759 ^ n10753 ^ x93 ;
  assign n10767 = ( x96 & ~n10677 ) | ( x96 & n10762 ) | ( ~n10677 & n10762 ) ;
  assign n10768 = ( x97 & ~n10674 ) | ( x97 & n10767 ) | ( ~n10674 & n10767 ) ;
  assign n10769 = ( x98 & ~n10671 ) | ( x98 & n10768 ) | ( ~n10671 & n10768 ) ;
  assign n10770 = ( x99 & ~n10668 ) | ( x99 & n10769 ) | ( ~n10668 & n10769 ) ;
  assign n10771 = ( x100 & ~n10665 ) | ( x100 & n10770 ) | ( ~n10665 & n10770 ) ;
  assign n10772 = ( x101 & ~n10739 ) | ( x101 & n10771 ) | ( ~n10739 & n10771 ) ;
  assign n10773 = ( x102 & ~n10662 ) | ( x102 & n10772 ) | ( ~n10662 & n10772 ) ;
  assign n10774 = ( x103 & ~n10659 ) | ( x103 & n10773 ) | ( ~n10659 & n10773 ) ;
  assign n10775 = ( x104 & ~n10656 ) | ( x104 & n10774 ) | ( ~n10656 & n10774 ) ;
  assign n10776 = ( x105 & ~n10653 ) | ( x105 & n10775 ) | ( ~n10653 & n10775 ) ;
  assign n10777 = ( x106 & ~n10650 ) | ( x106 & n10776 ) | ( ~n10650 & n10776 ) ;
  assign n10778 = ( x107 & ~n10647 ) | ( x107 & n10777 ) | ( ~n10647 & n10777 ) ;
  assign n10779 = ( x108 & ~n10599 ) | ( x108 & n10778 ) | ( ~n10599 & n10778 ) ;
  assign n10780 = ( x109 & ~n10596 ) | ( x109 & n10779 ) | ( ~n10596 & n10779 ) ;
  assign n10781 = ( x110 & ~n10580 ) | ( x110 & n10780 ) | ( ~n10580 & n10780 ) ;
  assign n10782 = ( x111 & ~n10715 ) | ( x111 & n10781 ) | ( ~n10715 & n10781 ) ;
  assign n10783 = ( x112 & ~n10577 ) | ( x112 & n10782 ) | ( ~n10577 & n10782 ) ;
  assign n10784 = ( x113 & ~n10574 ) | ( x113 & n10783 ) | ( ~n10574 & n10783 ) ;
  assign n10785 = ( x114 & ~n10582 ) | ( x114 & n10784 ) | ( ~n10582 & n10784 ) ;
  assign n10786 = ( x115 & ~n10570 ) | ( x115 & n10785 ) | ( ~n10570 & n10785 ) ;
  assign n10787 = ( x116 & ~n10567 ) | ( x116 & n10786 ) | ( ~n10567 & n10786 ) ;
  assign n10788 = ( x117 & ~n10564 ) | ( x117 & n10787 ) | ( ~n10564 & n10787 ) ;
  assign n10789 = ( x118 & ~n10561 ) | ( x118 & n10788 ) | ( ~n10561 & n10788 ) ;
  assign n10790 = ( x119 & ~n10758 ) | ( x119 & n10789 ) | ( ~n10758 & n10789 ) ;
  assign n10791 = ( n10757 & n10765 ) | ( n10757 & ~n10790 ) | ( n10765 & ~n10790 ) ;
  assign n10792 = n10790 | n10791 ;
  assign n10793 = ( ~n10719 & n10764 ) | ( ~n10719 & n10792 ) | ( n10764 & n10792 ) ;
  assign n10794 = n10793 ^ n10677 ^ 1'b0 ;
  assign n10795 = ( n10677 & n10763 ) | ( n10677 & ~n10794 ) | ( n10763 & ~n10794 ) ;
  assign n10796 = n10793 ^ n10759 ^ 1'b0 ;
  assign n10797 = ( n10759 & n10766 ) | ( n10759 & ~n10796 ) | ( n10766 & ~n10796 ) ;
  assign n10798 = n10793 ^ n10689 ^ 1'b0 ;
  assign n10799 = ( n10689 & n10754 ) | ( n10689 & ~n10798 ) | ( n10754 & ~n10798 ) ;
  assign n10800 = n10793 ^ n10605 ^ 1'b0 ;
  assign n10801 = ( n10605 & n10749 ) | ( n10605 & ~n10800 ) | ( n10749 & ~n10800 ) ;
  assign n10802 = n10793 ^ n10620 ^ 1'b0 ;
  assign n10803 = ( n10620 & n10741 ) | ( n10620 & ~n10802 ) | ( n10741 & ~n10802 ) ;
  assign n10804 = n10793 ^ n10736 ^ 1'b0 ;
  assign n10805 = ( n10736 & n10738 ) | ( n10736 & ~n10804 ) | ( n10738 & ~n10804 ) ;
  assign n10806 = n10793 ^ n10623 ^ 1'b0 ;
  assign n10807 = ( n10623 & n10734 ) | ( n10623 & ~n10806 ) | ( n10734 & ~n10806 ) ;
  assign n10808 = n10793 ^ n10629 ^ 1'b0 ;
  assign n10809 = ( n10629 & n10730 ) | ( n10629 & ~n10808 ) | ( n10730 & ~n10808 ) ;
  assign n10810 = n10793 ^ n10632 ^ 1'b0 ;
  assign n10811 = ( n10632 & n10727 ) | ( n10632 & ~n10810 ) | ( n10727 & ~n10810 ) ;
  assign n10812 = n10793 ^ n10584 ^ 1'b0 ;
  assign n10813 = ( n10584 & n10728 ) | ( n10584 & ~n10812 ) | ( n10728 & ~n10812 ) ;
  assign n10814 = n10793 ^ n10588 ^ 1'b0 ;
  assign n10815 = ( n10588 & n10714 ) | ( n10588 & ~n10814 ) | ( n10714 & ~n10814 ) ;
  assign n10816 = n10793 ^ n10707 ^ 1'b0 ;
  assign n10817 = ( n10700 & n10707 ) | ( n10700 & n10816 ) | ( n10707 & n10816 ) ;
  assign n10818 = n10764 & ~n10792 ;
  assign n10819 = ( n322 & n10764 ) | ( n322 & ~n10818 ) | ( n10764 & ~n10818 ) ;
  assign n10820 = n10789 ^ n10758 ^ x119 ;
  assign n10821 = n10793 ^ n10758 ^ 1'b0 ;
  assign n10822 = ( n10758 & n10820 ) | ( n10758 & ~n10821 ) | ( n10820 & ~n10821 ) ;
  assign n10823 = n10787 ^ n10564 ^ x117 ;
  assign n10824 = n10793 ^ n10564 ^ 1'b0 ;
  assign n10825 = ( n10564 & n10823 ) | ( n10564 & ~n10824 ) | ( n10823 & ~n10824 ) ;
  assign n10826 = n10786 ^ n10567 ^ x116 ;
  assign n10827 = n10793 ^ n10567 ^ 1'b0 ;
  assign n10828 = ( n10567 & n10826 ) | ( n10567 & ~n10827 ) | ( n10826 & ~n10827 ) ;
  assign n10829 = n10782 ^ n10577 ^ x112 ;
  assign n10830 = n10793 ^ n10577 ^ 1'b0 ;
  assign n10831 = ( n10577 & n10829 ) | ( n10577 & ~n10830 ) | ( n10829 & ~n10830 ) ;
  assign n10832 = n10780 ^ n10580 ^ x110 ;
  assign n10833 = n10793 ^ n10580 ^ 1'b0 ;
  assign n10834 = ( n10580 & n10832 ) | ( n10580 & ~n10833 ) | ( n10832 & ~n10833 ) ;
  assign n10835 = n10779 ^ n10596 ^ x109 ;
  assign n10836 = n10793 ^ n10596 ^ 1'b0 ;
  assign n10837 = ( n10596 & n10835 ) | ( n10596 & ~n10836 ) | ( n10835 & ~n10836 ) ;
  assign n10838 = n10778 ^ n10599 ^ x108 ;
  assign n10839 = n10793 ^ n10599 ^ 1'b0 ;
  assign n10840 = ( n10599 & n10838 ) | ( n10599 & ~n10839 ) | ( n10838 & ~n10839 ) ;
  assign n10841 = n10777 ^ n10647 ^ x107 ;
  assign n10842 = n10793 ^ n10647 ^ 1'b0 ;
  assign n10843 = ( n10647 & n10841 ) | ( n10647 & ~n10842 ) | ( n10841 & ~n10842 ) ;
  assign n10844 = n10776 ^ n10650 ^ x106 ;
  assign n10845 = n10793 ^ n10650 ^ 1'b0 ;
  assign n10846 = ( n10650 & n10844 ) | ( n10650 & ~n10845 ) | ( n10844 & ~n10845 ) ;
  assign n10847 = n10775 ^ n10653 ^ x105 ;
  assign n10848 = n10793 ^ n10653 ^ 1'b0 ;
  assign n10849 = ( n10653 & n10847 ) | ( n10653 & ~n10848 ) | ( n10847 & ~n10848 ) ;
  assign n10850 = n10774 ^ n10656 ^ x104 ;
  assign n10851 = n10793 ^ n10656 ^ 1'b0 ;
  assign n10852 = ( n10656 & n10850 ) | ( n10656 & ~n10851 ) | ( n10850 & ~n10851 ) ;
  assign n10853 = n10773 ^ n10659 ^ x103 ;
  assign n10854 = n10793 ^ n10659 ^ 1'b0 ;
  assign n10855 = ( n10659 & n10853 ) | ( n10659 & ~n10854 ) | ( n10853 & ~n10854 ) ;
  assign n10856 = n10767 ^ n10674 ^ x97 ;
  assign n10857 = n10793 ^ n10674 ^ 1'b0 ;
  assign n10858 = ( n10674 & n10856 ) | ( n10674 & ~n10857 ) | ( n10856 & ~n10857 ) ;
  assign n10859 = n10793 ^ n10611 ^ 1'b0 ;
  assign n10860 = ( n10611 & n10746 ) | ( n10611 & ~n10859 ) | ( n10746 & ~n10859 ) ;
  assign n10861 = n10793 ^ n10704 ^ 1'b0 ;
  assign n10862 = ( n10703 & n10704 ) | ( n10703 & n10861 ) | ( n10704 & n10861 ) ;
  assign n10863 = n10788 ^ n10561 ^ x118 ;
  assign n10864 = n10785 ^ n10570 ^ x115 ;
  assign n10865 = n10793 ^ n10570 ^ 1'b0 ;
  assign n10866 = ( n10570 & n10864 ) | ( n10570 & ~n10865 ) | ( n10864 & ~n10865 ) ;
  assign n10867 = n10784 ^ n10582 ^ x114 ;
  assign n10868 = n10793 ^ n10582 ^ 1'b0 ;
  assign n10869 = ( n10582 & n10867 ) | ( n10582 & ~n10868 ) | ( n10867 & ~n10868 ) ;
  assign n10870 = n10781 ^ n10715 ^ x111 ;
  assign n10871 = n10793 ^ n10715 ^ 1'b0 ;
  assign n10872 = ( n10715 & n10870 ) | ( n10715 & ~n10871 ) | ( n10870 & ~n10871 ) ;
  assign n10873 = n10772 ^ n10662 ^ x102 ;
  assign n10874 = n10793 ^ n10662 ^ 1'b0 ;
  assign n10875 = ( n10662 & n10873 ) | ( n10662 & ~n10874 ) | ( n10873 & ~n10874 ) ;
  assign n10876 = n10771 ^ n10739 ^ x101 ;
  assign n10877 = n10793 ^ n10739 ^ 1'b0 ;
  assign n10878 = ( n10739 & n10876 ) | ( n10739 & ~n10877 ) | ( n10876 & ~n10877 ) ;
  assign n10879 = n10770 ^ n10665 ^ x100 ;
  assign n10880 = n10793 ^ n10665 ^ 1'b0 ;
  assign n10881 = ( n10665 & n10879 ) | ( n10665 & ~n10880 ) | ( n10879 & ~n10880 ) ;
  assign n10882 = n10769 ^ n10668 ^ x99 ;
  assign n10883 = n10793 ^ n10668 ^ 1'b0 ;
  assign n10884 = ( n10668 & n10882 ) | ( n10668 & ~n10883 ) | ( n10882 & ~n10883 ) ;
  assign n10885 = n10768 ^ n10671 ^ x98 ;
  assign n10886 = n10793 ^ n10671 ^ 1'b0 ;
  assign n10887 = ( n10671 & n10885 ) | ( n10671 & ~n10886 ) | ( n10885 & ~n10886 ) ;
  assign n10888 = n10760 ^ n10683 ^ x94 ;
  assign n10889 = n10793 ^ n10683 ^ 1'b0 ;
  assign n10890 = ( n10683 & n10888 ) | ( n10683 & ~n10889 ) | ( n10888 & ~n10889 ) ;
  assign n10891 = n10752 ^ n10686 ^ x92 ;
  assign n10892 = n10793 ^ n10686 ^ 1'b0 ;
  assign n10893 = ( n10686 & n10891 ) | ( n10686 & ~n10892 ) | ( n10891 & ~n10892 ) ;
  assign n10894 = n10750 ^ n10602 ^ x90 ;
  assign n10895 = n10793 ^ n10602 ^ 1'b0 ;
  assign n10896 = ( n10602 & n10894 ) | ( n10602 & ~n10895 ) | ( n10894 & ~n10895 ) ;
  assign n10897 = n10747 ^ n10608 ^ x88 ;
  assign n10898 = n10793 ^ n10608 ^ 1'b0 ;
  assign n10899 = ( n10608 & n10897 ) | ( n10608 & ~n10898 ) | ( n10897 & ~n10898 ) ;
  assign n10900 = n10744 ^ n10735 ^ x86 ;
  assign n10901 = n10793 ^ n10735 ^ 1'b0 ;
  assign n10902 = ( n10735 & n10900 ) | ( n10735 & ~n10901 ) | ( n10900 & ~n10901 ) ;
  assign n10903 = n10743 ^ n10614 ^ x85 ;
  assign n10904 = n10793 ^ n10614 ^ 1'b0 ;
  assign n10905 = ( n10614 & n10903 ) | ( n10614 & ~n10904 ) | ( n10903 & ~n10904 ) ;
  assign n10906 = n10742 ^ n10617 ^ x84 ;
  assign n10907 = n10793 ^ n10617 ^ 1'b0 ;
  assign n10908 = ( n10617 & n10906 ) | ( n10617 & ~n10907 ) | ( n10906 & ~n10907 ) ;
  assign n10909 = n10731 ^ n10626 ^ x80 ;
  assign n10910 = n10793 ^ n10626 ^ 1'b0 ;
  assign n10911 = ( n10626 & n10909 ) | ( n10626 & ~n10910 ) | ( n10909 & ~n10910 ) ;
  assign n10912 = n10724 ^ n10586 ^ x76 ;
  assign n10913 = n10793 ^ n10586 ^ 1'b0 ;
  assign n10914 = ( n10586 & n10912 ) | ( n10586 & ~n10913 ) | ( n10912 & ~n10913 ) ;
  assign n10915 = n10723 ^ n10635 ^ x75 ;
  assign n10916 = n10793 ^ n10561 ^ 1'b0 ;
  assign n10917 = ( n10561 & n10863 ) | ( n10561 & ~n10916 ) | ( n10863 & ~n10916 ) ;
  assign n10918 = n10793 ^ n10635 ^ 1'b0 ;
  assign n10919 = ( n10635 & n10915 ) | ( n10635 & ~n10918 ) | ( n10915 & ~n10918 ) ;
  assign n10920 = n10722 ^ n10721 ^ x74 ;
  assign n10921 = n10793 ^ n10722 ^ 1'b0 ;
  assign n10922 = ( n10722 & n10920 ) | ( n10722 & ~n10921 ) | ( n10920 & ~n10921 ) ;
  assign n10923 = n10720 ^ n10638 ^ x73 ;
  assign n10924 = n10793 ^ n10638 ^ 1'b0 ;
  assign n10925 = ( n10638 & n10923 ) | ( n10638 & ~n10924 ) | ( n10923 & ~n10924 ) ;
  assign n10926 = n10712 ^ n10641 ^ x71 ;
  assign n10927 = n10793 ^ n10641 ^ 1'b0 ;
  assign n10928 = ( n10641 & n10926 ) | ( n10641 & ~n10927 ) | ( n10926 & ~n10927 ) ;
  assign n10929 = n10711 ^ n10705 ^ x70 ;
  assign n10930 = n10793 ^ n10705 ^ 1'b0 ;
  assign n10931 = ( n10705 & n10929 ) | ( n10705 & ~n10930 ) | ( n10929 & ~n10930 ) ;
  assign n10932 = n10710 ^ n10590 ^ x69 ;
  assign n10933 = n10793 ^ n10590 ^ 1'b0 ;
  assign n10934 = ( n10590 & n10932 ) | ( n10590 & ~n10933 ) | ( n10932 & ~n10933 ) ;
  assign n10935 = n10709 ^ n10644 ^ x68 ;
  assign n10936 = n10793 ^ n10644 ^ 1'b0 ;
  assign n10937 = ( n10644 & n10935 ) | ( n10644 & ~n10936 ) | ( n10935 & ~n10936 ) ;
  assign n10938 = n10708 ^ n10592 ^ x67 ;
  assign n10939 = n10793 ^ n10592 ^ 1'b0 ;
  assign n10940 = ( n10592 & n10938 ) | ( n10592 & ~n10939 ) | ( n10938 & ~n10939 ) ;
  assign n10941 = x64 & n10793 ;
  assign n10942 = n10941 ^ x64 ^ x7 ;
  assign n10943 = n10942 ^ n8096 ^ x65 ;
  assign n10944 = ( x65 & n8096 ) | ( x65 & n10943 ) | ( n8096 & n10943 ) ;
  assign n10945 = n10761 ^ n10680 ^ x95 ;
  assign n10946 = n10793 ^ n10574 ^ 1'b0 ;
  assign n10947 = n10944 ^ n10862 ^ x66 ;
  assign n10948 = ( x66 & n10944 ) | ( x66 & n10947 ) | ( n10944 & n10947 ) ;
  assign n10949 = ( x67 & ~n10817 ) | ( x67 & n10948 ) | ( ~n10817 & n10948 ) ;
  assign n10950 = ( x68 & ~n10940 ) | ( x68 & n10949 ) | ( ~n10940 & n10949 ) ;
  assign n10951 = x6 & ~n8332 ;
  assign n10952 = ( x69 & ~n10937 ) | ( x69 & n10950 ) | ( ~n10937 & n10950 ) ;
  assign n10953 = n10949 ^ n10940 ^ x68 ;
  assign n10954 = ( x70 & ~n10934 ) | ( x70 & n10952 ) | ( ~n10934 & n10952 ) ;
  assign n10955 = ( x71 & ~n10931 ) | ( x71 & n10954 ) | ( ~n10931 & n10954 ) ;
  assign n10956 = n10955 ^ n10928 ^ x72 ;
  assign n10957 = ( x72 & ~n10928 ) | ( x72 & n10955 ) | ( ~n10928 & n10955 ) ;
  assign n10958 = ( x73 & ~n10815 ) | ( x73 & n10957 ) | ( ~n10815 & n10957 ) ;
  assign n10959 = n10950 ^ n10937 ^ x69 ;
  assign n10960 = ( x74 & ~n10925 ) | ( x74 & n10958 ) | ( ~n10925 & n10958 ) ;
  assign n10961 = ( x75 & ~n10922 ) | ( x75 & n10960 ) | ( ~n10922 & n10960 ) ;
  assign n10962 = ( x76 & ~n10919 ) | ( x76 & n10961 ) | ( ~n10919 & n10961 ) ;
  assign n10963 = ( x77 & ~n10914 ) | ( x77 & n10962 ) | ( ~n10914 & n10962 ) ;
  assign n10964 = ( x78 & ~n10813 ) | ( x78 & n10963 ) | ( ~n10813 & n10963 ) ;
  assign n10965 = ( x79 & ~n10811 ) | ( x79 & n10964 ) | ( ~n10811 & n10964 ) ;
  assign n10966 = ( x80 & ~n10809 ) | ( x80 & n10965 ) | ( ~n10809 & n10965 ) ;
  assign n10967 = ( x81 & ~n10911 ) | ( x81 & n10966 ) | ( ~n10911 & n10966 ) ;
  assign n10968 = ( x82 & ~n10807 ) | ( x82 & n10967 ) | ( ~n10807 & n10967 ) ;
  assign n10969 = n10968 ^ n10805 ^ x83 ;
  assign n10970 = n10965 ^ n10809 ^ x80 ;
  assign n10971 = ( x83 & ~n10805 ) | ( x83 & n10968 ) | ( ~n10805 & n10968 ) ;
  assign n10972 = ( x84 & ~n10803 ) | ( x84 & n10971 ) | ( ~n10803 & n10971 ) ;
  assign n10973 = n10948 ^ n10817 ^ x67 ;
  assign n10974 = n10971 ^ n10803 ^ x84 ;
  assign n10975 = n10966 ^ n10911 ^ x81 ;
  assign n10976 = n10952 ^ n10934 ^ x70 ;
  assign n10977 = n10783 ^ n10574 ^ x113 ;
  assign n10978 = ( x85 & ~n10908 ) | ( x85 & n10972 ) | ( ~n10908 & n10972 ) ;
  assign n10979 = ( n10574 & ~n10946 ) | ( n10574 & n10977 ) | ( ~n10946 & n10977 ) ;
  assign n10980 = ( x86 & ~n10905 ) | ( x86 & n10978 ) | ( ~n10905 & n10978 ) ;
  assign n10981 = ( x87 & ~n10902 ) | ( x87 & n10980 ) | ( ~n10902 & n10980 ) ;
  assign n10982 = n10793 ^ n10680 ^ 1'b0 ;
  assign n10983 = n10981 ^ n10860 ^ x88 ;
  assign n10984 = n10972 ^ n10908 ^ x85 ;
  assign n10985 = n10962 ^ n10914 ^ x77 ;
  assign n10986 = n10960 ^ n10922 ^ x75 ;
  assign n10987 = n10963 ^ n10813 ^ x78 ;
  assign n10988 = n10957 ^ n10815 ^ x73 ;
  assign n10989 = n10954 ^ n10931 ^ x71 ;
  assign n10990 = n10978 ^ n10905 ^ x86 ;
  assign n10991 = ( n10680 & n10945 ) | ( n10680 & ~n10982 ) | ( n10945 & ~n10982 ) ;
  assign n10992 = n10964 ^ n10811 ^ x79 ;
  assign n10993 = n10961 ^ n10919 ^ x76 ;
  assign n10994 = n10958 ^ n10925 ^ x74 ;
  assign n10995 = ( x88 & ~n10860 ) | ( x88 & n10981 ) | ( ~n10860 & n10981 ) ;
  assign n10996 = ( x89 & ~n10899 ) | ( x89 & n10995 ) | ( ~n10899 & n10995 ) ;
  assign n10997 = ( x90 & ~n10801 ) | ( x90 & n10996 ) | ( ~n10801 & n10996 ) ;
  assign n10998 = ( x91 & ~n10896 ) | ( x91 & n10997 ) | ( ~n10896 & n10997 ) ;
  assign n10999 = n10967 ^ n10807 ^ x82 ;
  assign n11000 = n10997 ^ n10896 ^ x91 ;
  assign n11001 = n10995 ^ n10899 ^ x89 ;
  assign n11002 = n10996 ^ n10801 ^ x90 ;
  assign n11003 = n10980 ^ n10902 ^ x87 ;
  assign n11004 = n10998 ^ n10799 ^ x92 ;
  assign n11005 = ( x92 & ~n10799 ) | ( x92 & n10998 ) | ( ~n10799 & n10998 ) ;
  assign n11006 = ( x93 & ~n10893 ) | ( x93 & n11005 ) | ( ~n10893 & n11005 ) ;
  assign n11007 = ( x94 & ~n10797 ) | ( x94 & n11006 ) | ( ~n10797 & n11006 ) ;
  assign n11008 = ( x95 & ~n10890 ) | ( x95 & n11007 ) | ( ~n10890 & n11007 ) ;
  assign n11009 = ( x96 & ~n10991 ) | ( x96 & n11008 ) | ( ~n10991 & n11008 ) ;
  assign n11010 = ( x97 & ~n10795 ) | ( x97 & n11009 ) | ( ~n10795 & n11009 ) ;
  assign n11011 = ( x98 & ~n10858 ) | ( x98 & n11010 ) | ( ~n10858 & n11010 ) ;
  assign n11012 = ( x99 & ~n10887 ) | ( x99 & n11011 ) | ( ~n10887 & n11011 ) ;
  assign n11013 = ( x100 & ~n10884 ) | ( x100 & n11012 ) | ( ~n10884 & n11012 ) ;
  assign n11014 = ( x101 & ~n10881 ) | ( x101 & n11013 ) | ( ~n10881 & n11013 ) ;
  assign n11015 = ( x102 & ~n10878 ) | ( x102 & n11014 ) | ( ~n10878 & n11014 ) ;
  assign n11016 = ( x103 & ~n10875 ) | ( x103 & n11015 ) | ( ~n10875 & n11015 ) ;
  assign n11017 = ( x104 & ~n10855 ) | ( x104 & n11016 ) | ( ~n10855 & n11016 ) ;
  assign n11018 = ( x105 & ~n10852 ) | ( x105 & n11017 ) | ( ~n10852 & n11017 ) ;
  assign n11019 = ( x106 & ~n10849 ) | ( x106 & n11018 ) | ( ~n10849 & n11018 ) ;
  assign n11020 = ( x107 & ~n10846 ) | ( x107 & n11019 ) | ( ~n10846 & n11019 ) ;
  assign n11021 = ( x108 & ~n10843 ) | ( x108 & n11020 ) | ( ~n10843 & n11020 ) ;
  assign n11022 = ( x109 & ~n10840 ) | ( x109 & n11021 ) | ( ~n10840 & n11021 ) ;
  assign n11023 = ( x110 & ~n10837 ) | ( x110 & n11022 ) | ( ~n10837 & n11022 ) ;
  assign n11024 = ( x111 & ~n10834 ) | ( x111 & n11023 ) | ( ~n10834 & n11023 ) ;
  assign n11025 = ( x112 & ~n10872 ) | ( x112 & n11024 ) | ( ~n10872 & n11024 ) ;
  assign n11026 = ( x113 & ~n10831 ) | ( x113 & n11025 ) | ( ~n10831 & n11025 ) ;
  assign n11027 = ( x114 & ~n10979 ) | ( x114 & n11026 ) | ( ~n10979 & n11026 ) ;
  assign n11028 = ( x115 & ~n10869 ) | ( x115 & n11027 ) | ( ~n10869 & n11027 ) ;
  assign n11029 = ( x116 & ~n10866 ) | ( x116 & n11028 ) | ( ~n10866 & n11028 ) ;
  assign n11030 = ( x117 & ~n10828 ) | ( x117 & n11029 ) | ( ~n10828 & n11029 ) ;
  assign n11031 = ( x118 & ~n10825 ) | ( x118 & n11030 ) | ( ~n10825 & n11030 ) ;
  assign n11032 = ( x119 & ~n10917 ) | ( x119 & n11031 ) | ( ~n10917 & n11031 ) ;
  assign n11033 = ( x120 & ~n10822 ) | ( x120 & n11032 ) | ( ~n10822 & n11032 ) ;
  assign n11034 = ( x121 & ~n10819 ) | ( x121 & n11033 ) | ( ~n10819 & n11033 ) ;
  assign n11035 = n155 | n11034 ;
  assign n11036 = n8327 | n11034 ;
  assign n11037 = ( x6 & ~n11034 ) | ( x6 & n11036 ) | ( ~n11034 & n11036 ) ;
  assign n11038 = ( n10951 & n11036 ) | ( n10951 & n11037 ) | ( n11036 & n11037 ) ;
  assign n11039 = n11035 ^ n10937 ^ 1'b0 ;
  assign n11040 = n11035 ^ n10947 ^ 1'b0 ;
  assign n11041 = ( n10862 & n10947 ) | ( n10862 & n11040 ) | ( n10947 & n11040 ) ;
  assign n11042 = n11035 ^ n10928 ^ 1'b0 ;
  assign n11043 = ( n10928 & n10956 ) | ( n10928 & ~n11042 ) | ( n10956 & ~n11042 ) ;
  assign n11044 = ( n10937 & n10959 ) | ( n10937 & ~n11039 ) | ( n10959 & ~n11039 ) ;
  assign n11045 = n11035 ^ n10934 ^ 1'b0 ;
  assign n11046 = n11035 ^ n10817 ^ 1'b0 ;
  assign n11047 = n11035 ^ n10931 ^ 1'b0 ;
  assign n11048 = n11035 ^ n10925 ^ 1'b0 ;
  assign n11049 = ( n10931 & n10989 ) | ( n10931 & ~n11047 ) | ( n10989 & ~n11047 ) ;
  assign n11050 = ( n10925 & n10994 ) | ( n10925 & ~n11048 ) | ( n10994 & ~n11048 ) ;
  assign n11051 = ( n10934 & n10976 ) | ( n10934 & ~n11045 ) | ( n10976 & ~n11045 ) ;
  assign n11052 = ( n10817 & n10973 ) | ( n10817 & ~n11046 ) | ( n10973 & ~n11046 ) ;
  assign n11053 = n11035 ^ n10815 ^ 1'b0 ;
  assign n11054 = n11035 ^ n10940 ^ 1'b0 ;
  assign n11055 = ( n10815 & n10988 ) | ( n10815 & ~n11053 ) | ( n10988 & ~n11053 ) ;
  assign n11056 = ( n10940 & n10953 ) | ( n10940 & ~n11054 ) | ( n10953 & ~n11054 ) ;
  assign n11057 = n11031 ^ n10917 ^ x119 ;
  assign n11058 = n11035 ^ n10917 ^ 1'b0 ;
  assign n11059 = ( n10917 & n11057 ) | ( n10917 & ~n11058 ) | ( n11057 & ~n11058 ) ;
  assign n11060 = n11030 ^ n10825 ^ x118 ;
  assign n11061 = n11035 ^ n10799 ^ 1'b0 ;
  assign n11062 = ( n10799 & n11004 ) | ( n10799 & ~n11061 ) | ( n11004 & ~n11061 ) ;
  assign n11063 = n11035 ^ n10896 ^ 1'b0 ;
  assign n11064 = ( n10896 & n11000 ) | ( n10896 & ~n11063 ) | ( n11000 & ~n11063 ) ;
  assign n11065 = n11035 ^ n10801 ^ 1'b0 ;
  assign n11066 = ( n10801 & n11002 ) | ( n10801 & ~n11065 ) | ( n11002 & ~n11065 ) ;
  assign n11067 = n11035 ^ n10899 ^ 1'b0 ;
  assign n11068 = ( n10899 & n11001 ) | ( n10899 & ~n11067 ) | ( n11001 & ~n11067 ) ;
  assign n11069 = n11035 ^ n10860 ^ 1'b0 ;
  assign n11070 = ( n10860 & n10983 ) | ( n10860 & ~n11069 ) | ( n10983 & ~n11069 ) ;
  assign n11071 = n11035 ^ n10902 ^ 1'b0 ;
  assign n11072 = ( n10902 & n11003 ) | ( n10902 & ~n11071 ) | ( n11003 & ~n11071 ) ;
  assign n11073 = n11035 ^ n10905 ^ 1'b0 ;
  assign n11074 = ( n10905 & n10990 ) | ( n10905 & ~n11073 ) | ( n10990 & ~n11073 ) ;
  assign n11075 = n11035 ^ n10908 ^ 1'b0 ;
  assign n11076 = ( n10908 & n10984 ) | ( n10908 & ~n11075 ) | ( n10984 & ~n11075 ) ;
  assign n11077 = n11035 ^ n10803 ^ 1'b0 ;
  assign n11078 = ( n10803 & n10974 ) | ( n10803 & ~n11077 ) | ( n10974 & ~n11077 ) ;
  assign n11079 = n11035 ^ n10805 ^ 1'b0 ;
  assign n11080 = ( n10805 & n10969 ) | ( n10805 & ~n11079 ) | ( n10969 & ~n11079 ) ;
  assign n11081 = n11035 ^ n10807 ^ 1'b0 ;
  assign n11082 = ( n10807 & n10999 ) | ( n10807 & ~n11081 ) | ( n10999 & ~n11081 ) ;
  assign n11083 = n11035 ^ n10911 ^ 1'b0 ;
  assign n11084 = ( n10911 & n10975 ) | ( n10911 & ~n11083 ) | ( n10975 & ~n11083 ) ;
  assign n11085 = n11035 ^ n10809 ^ 1'b0 ;
  assign n11086 = ( n10809 & n10970 ) | ( n10809 & ~n11085 ) | ( n10970 & ~n11085 ) ;
  assign n11087 = n11035 ^ n10825 ^ 1'b0 ;
  assign n11088 = ( n10825 & n11060 ) | ( n10825 & ~n11087 ) | ( n11060 & ~n11087 ) ;
  assign n11089 = n11035 ^ n10811 ^ 1'b0 ;
  assign n11090 = ( n10811 & n10992 ) | ( n10811 & ~n11089 ) | ( n10992 & ~n11089 ) ;
  assign n11091 = n11035 ^ n10813 ^ 1'b0 ;
  assign n11092 = ( n10813 & n10987 ) | ( n10813 & ~n11091 ) | ( n10987 & ~n11091 ) ;
  assign n11093 = n11035 ^ n10914 ^ 1'b0 ;
  assign n11094 = ( n10914 & n10985 ) | ( n10914 & ~n11093 ) | ( n10985 & ~n11093 ) ;
  assign n11095 = n11035 ^ n10919 ^ 1'b0 ;
  assign n11096 = ( n10919 & n10993 ) | ( n10919 & ~n11095 ) | ( n10993 & ~n11095 ) ;
  assign n11097 = n11035 ^ n10922 ^ 1'b0 ;
  assign n11098 = ( n10922 & n10986 ) | ( n10922 & ~n11097 ) | ( n10986 & ~n11097 ) ;
  assign n11099 = n11035 ^ n10943 ^ 1'b0 ;
  assign n11100 = ( n10942 & n10943 ) | ( n10942 & n11099 ) | ( n10943 & n11099 ) ;
  assign n11101 = n11032 ^ n10822 ^ x120 ;
  assign n11102 = n11035 ^ n10822 ^ 1'b0 ;
  assign n11103 = ( n10822 & n11101 ) | ( n10822 & ~n11102 ) | ( n11101 & ~n11102 ) ;
  assign n11104 = n11029 ^ n10828 ^ x117 ;
  assign n11105 = n11035 ^ n10828 ^ 1'b0 ;
  assign n11106 = ( n10828 & n11104 ) | ( n10828 & ~n11105 ) | ( n11104 & ~n11105 ) ;
  assign n11107 = n11028 ^ n10866 ^ x116 ;
  assign n11108 = n11035 ^ n10866 ^ 1'b0 ;
  assign n11109 = ( n10866 & n11107 ) | ( n10866 & ~n11108 ) | ( n11107 & ~n11108 ) ;
  assign n11110 = n11027 ^ n10869 ^ x115 ;
  assign n11111 = n11035 ^ n10869 ^ 1'b0 ;
  assign n11112 = ( n10869 & n11110 ) | ( n10869 & ~n11111 ) | ( n11110 & ~n11111 ) ;
  assign n11113 = n11026 ^ n10979 ^ x114 ;
  assign n11114 = n11035 ^ n10979 ^ 1'b0 ;
  assign n11115 = ( n10979 & n11113 ) | ( n10979 & ~n11114 ) | ( n11113 & ~n11114 ) ;
  assign n11116 = n11025 ^ n10831 ^ x113 ;
  assign n11117 = n11035 ^ n10831 ^ 1'b0 ;
  assign n11118 = ( n10831 & n11116 ) | ( n10831 & ~n11117 ) | ( n11116 & ~n11117 ) ;
  assign n11119 = n11024 ^ n10872 ^ x112 ;
  assign n11120 = n11035 ^ n10872 ^ 1'b0 ;
  assign n11121 = ( n10872 & n11119 ) | ( n10872 & ~n11120 ) | ( n11119 & ~n11120 ) ;
  assign n11122 = n11023 ^ n10834 ^ x111 ;
  assign n11123 = n11035 ^ n10834 ^ 1'b0 ;
  assign n11124 = ( n10834 & n11122 ) | ( n10834 & ~n11123 ) | ( n11122 & ~n11123 ) ;
  assign n11125 = n11022 ^ n10837 ^ x110 ;
  assign n11126 = n11035 ^ n10837 ^ 1'b0 ;
  assign n11127 = ( n10837 & n11125 ) | ( n10837 & ~n11126 ) | ( n11125 & ~n11126 ) ;
  assign n11128 = n11021 ^ n10840 ^ x109 ;
  assign n11129 = n11035 ^ n10840 ^ 1'b0 ;
  assign n11130 = ( n10840 & n11128 ) | ( n10840 & ~n11129 ) | ( n11128 & ~n11129 ) ;
  assign n11131 = n11020 ^ n10843 ^ x108 ;
  assign n11132 = n11035 ^ n10843 ^ 1'b0 ;
  assign n11133 = ( n10843 & n11131 ) | ( n10843 & ~n11132 ) | ( n11131 & ~n11132 ) ;
  assign n11134 = n11019 ^ n10846 ^ x107 ;
  assign n11135 = n11035 ^ n10846 ^ 1'b0 ;
  assign n11136 = ( n10846 & n11134 ) | ( n10846 & ~n11135 ) | ( n11134 & ~n11135 ) ;
  assign n11137 = n11018 ^ n10849 ^ x106 ;
  assign n11138 = n11035 ^ n10849 ^ 1'b0 ;
  assign n11139 = ( n10849 & n11137 ) | ( n10849 & ~n11138 ) | ( n11137 & ~n11138 ) ;
  assign n11140 = n11017 ^ n10852 ^ x105 ;
  assign n11141 = n11035 ^ n10852 ^ 1'b0 ;
  assign n11142 = ( n10852 & n11140 ) | ( n10852 & ~n11141 ) | ( n11140 & ~n11141 ) ;
  assign n11143 = n11016 ^ n10855 ^ x104 ;
  assign n11144 = n11035 ^ n10855 ^ 1'b0 ;
  assign n11145 = ( n10855 & n11143 ) | ( n10855 & ~n11144 ) | ( n11143 & ~n11144 ) ;
  assign n11146 = n11015 ^ n10875 ^ x103 ;
  assign n11147 = n11035 ^ n10875 ^ 1'b0 ;
  assign n11148 = ( n10875 & n11146 ) | ( n10875 & ~n11147 ) | ( n11146 & ~n11147 ) ;
  assign n11149 = n11014 ^ n10878 ^ x102 ;
  assign n11150 = n11035 ^ n10878 ^ 1'b0 ;
  assign n11151 = ( n10878 & n11149 ) | ( n10878 & ~n11150 ) | ( n11149 & ~n11150 ) ;
  assign n11152 = n11013 ^ n10881 ^ x101 ;
  assign n11153 = n11035 ^ n10881 ^ 1'b0 ;
  assign n11154 = ( n10881 & n11152 ) | ( n10881 & ~n11153 ) | ( n11152 & ~n11153 ) ;
  assign n11155 = n11012 ^ n10884 ^ x100 ;
  assign n11156 = n11035 ^ n10884 ^ 1'b0 ;
  assign n11157 = ( n10884 & n11155 ) | ( n10884 & ~n11156 ) | ( n11155 & ~n11156 ) ;
  assign n11158 = n11011 ^ n10887 ^ x99 ;
  assign n11159 = n11035 ^ n10887 ^ 1'b0 ;
  assign n11160 = ( n10887 & n11158 ) | ( n10887 & ~n11159 ) | ( n11158 & ~n11159 ) ;
  assign n11161 = n11010 ^ n10858 ^ x98 ;
  assign n11162 = n11035 ^ n10858 ^ 1'b0 ;
  assign n11163 = ( n10858 & n11161 ) | ( n10858 & ~n11162 ) | ( n11161 & ~n11162 ) ;
  assign n11164 = n11009 ^ n10795 ^ x97 ;
  assign n11165 = n11035 ^ n10795 ^ 1'b0 ;
  assign n11166 = ( n10795 & n11164 ) | ( n10795 & ~n11165 ) | ( n11164 & ~n11165 ) ;
  assign n11167 = n11008 ^ n10991 ^ x96 ;
  assign n11168 = n11035 ^ n10991 ^ 1'b0 ;
  assign n11169 = ( n10991 & n11167 ) | ( n10991 & ~n11168 ) | ( n11167 & ~n11168 ) ;
  assign n11170 = n11007 ^ n10890 ^ x95 ;
  assign n11171 = n11035 ^ n10890 ^ 1'b0 ;
  assign n11172 = ( n10890 & n11170 ) | ( n10890 & ~n11171 ) | ( n11170 & ~n11171 ) ;
  assign n11173 = n11006 ^ n10797 ^ x94 ;
  assign n11174 = n11035 ^ n10797 ^ 1'b0 ;
  assign n11175 = ( n10797 & n11173 ) | ( n10797 & ~n11174 ) | ( n11173 & ~n11174 ) ;
  assign n11176 = n11005 ^ n10893 ^ x93 ;
  assign n11177 = n11035 ^ n10893 ^ 1'b0 ;
  assign n11178 = ( n10893 & n11176 ) | ( n10893 & ~n11177 ) | ( n11176 & ~n11177 ) ;
  assign n11179 = n11038 ^ n8326 ^ x65 ;
  assign n11180 = ( x65 & n8326 ) | ( x65 & n11179 ) | ( n8326 & n11179 ) ;
  assign n11181 = n11180 ^ n11100 ^ x66 ;
  assign n11182 = ( x66 & n11180 ) | ( x66 & n11181 ) | ( n11180 & n11181 ) ;
  assign n11183 = ( x67 & ~n11041 ) | ( x67 & n11182 ) | ( ~n11041 & n11182 ) ;
  assign n11184 = ( x68 & ~n11052 ) | ( x68 & n11183 ) | ( ~n11052 & n11183 ) ;
  assign n11185 = ( x69 & ~n11056 ) | ( x69 & n11184 ) | ( ~n11056 & n11184 ) ;
  assign n11186 = ( x70 & ~n11044 ) | ( x70 & n11185 ) | ( ~n11044 & n11185 ) ;
  assign n11187 = ( x71 & ~n11051 ) | ( x71 & n11186 ) | ( ~n11051 & n11186 ) ;
  assign n11188 = ( x72 & ~n11049 ) | ( x72 & n11187 ) | ( ~n11049 & n11187 ) ;
  assign n11189 = ( x73 & ~n11043 ) | ( x73 & n11188 ) | ( ~n11043 & n11188 ) ;
  assign n11190 = ( x74 & ~n11055 ) | ( x74 & n11189 ) | ( ~n11055 & n11189 ) ;
  assign n11191 = ( x75 & ~n11050 ) | ( x75 & n11190 ) | ( ~n11050 & n11190 ) ;
  assign n11192 = ( x76 & ~n11098 ) | ( x76 & n11191 ) | ( ~n11098 & n11191 ) ;
  assign n11193 = ( x77 & ~n11096 ) | ( x77 & n11192 ) | ( ~n11096 & n11192 ) ;
  assign n11194 = ( x78 & ~n11094 ) | ( x78 & n11193 ) | ( ~n11094 & n11193 ) ;
  assign n11195 = ( x79 & ~n11092 ) | ( x79 & n11194 ) | ( ~n11092 & n11194 ) ;
  assign n11196 = ( x80 & ~n11090 ) | ( x80 & n11195 ) | ( ~n11090 & n11195 ) ;
  assign n11197 = ( x81 & ~n11086 ) | ( x81 & n11196 ) | ( ~n11086 & n11196 ) ;
  assign n11198 = ( x82 & ~n11084 ) | ( x82 & n11197 ) | ( ~n11084 & n11197 ) ;
  assign n11199 = ( x83 & ~n11082 ) | ( x83 & n11198 ) | ( ~n11082 & n11198 ) ;
  assign n11200 = n10819 & n11035 ;
  assign n11201 = ( x84 & ~n11080 ) | ( x84 & n11199 ) | ( ~n11080 & n11199 ) ;
  assign n11202 = ( x85 & ~n11078 ) | ( x85 & n11201 ) | ( ~n11078 & n11201 ) ;
  assign n11203 = ( x86 & ~n11076 ) | ( x86 & n11202 ) | ( ~n11076 & n11202 ) ;
  assign n11204 = ( x87 & ~n11074 ) | ( x87 & n11203 ) | ( ~n11074 & n11203 ) ;
  assign n11205 = ( x88 & ~n11072 ) | ( x88 & n11204 ) | ( ~n11072 & n11204 ) ;
  assign n11206 = ( x89 & ~n11070 ) | ( x89 & n11205 ) | ( ~n11070 & n11205 ) ;
  assign n11207 = ( x90 & ~n11068 ) | ( x90 & n11206 ) | ( ~n11068 & n11206 ) ;
  assign n11208 = ( x91 & ~n11066 ) | ( x91 & n11207 ) | ( ~n11066 & n11207 ) ;
  assign n11209 = ( x92 & ~n11064 ) | ( x92 & n11208 ) | ( ~n11064 & n11208 ) ;
  assign n11210 = ( x93 & ~n11062 ) | ( x93 & n11209 ) | ( ~n11062 & n11209 ) ;
  assign n11211 = ( x94 & ~n11178 ) | ( x94 & n11210 ) | ( ~n11178 & n11210 ) ;
  assign n11212 = ( x95 & ~n11175 ) | ( x95 & n11211 ) | ( ~n11175 & n11211 ) ;
  assign n11213 = n322 | n11200 ;
  assign n11214 = n155 & n11213 ;
  assign n11215 = n155 & n10819 ;
  assign n11216 = ( x96 & ~n11172 ) | ( x96 & n11212 ) | ( ~n11172 & n11212 ) ;
  assign n11217 = ( x97 & ~n11169 ) | ( x97 & n11216 ) | ( ~n11169 & n11216 ) ;
  assign n11218 = ( x98 & ~n11166 ) | ( x98 & n11217 ) | ( ~n11166 & n11217 ) ;
  assign n11219 = ( x99 & ~n11163 ) | ( x99 & n11218 ) | ( ~n11163 & n11218 ) ;
  assign n11220 = n11192 ^ n11096 ^ x77 ;
  assign n11221 = n11191 ^ n11098 ^ x76 ;
  assign n11222 = n11190 ^ n11050 ^ x75 ;
  assign n11223 = n11189 ^ n11055 ^ x74 ;
  assign n11224 = n11188 ^ n11043 ^ x73 ;
  assign n11225 = n11187 ^ n11049 ^ x72 ;
  assign n11226 = n11186 ^ n11051 ^ x71 ;
  assign n11227 = n11185 ^ n11044 ^ x70 ;
  assign n11228 = n11184 ^ n11056 ^ x69 ;
  assign n11229 = n11182 ^ n11041 ^ x67 ;
  assign n11230 = ( x122 & n8330 ) | ( x122 & ~n11200 ) | ( n8330 & ~n11200 ) ;
  assign n11231 = ( x100 & ~n11160 ) | ( x100 & n11219 ) | ( ~n11160 & n11219 ) ;
  assign n11232 = ( x101 & ~n11157 ) | ( x101 & n11231 ) | ( ~n11157 & n11231 ) ;
  assign n11233 = ( x102 & ~n11154 ) | ( x102 & n11232 ) | ( ~n11154 & n11232 ) ;
  assign n11234 = ( x103 & ~n11151 ) | ( x103 & n11233 ) | ( ~n11151 & n11233 ) ;
  assign n11235 = ( x104 & ~n11148 ) | ( x104 & n11234 ) | ( ~n11148 & n11234 ) ;
  assign n11236 = ( x105 & ~n11145 ) | ( x105 & n11235 ) | ( ~n11145 & n11235 ) ;
  assign n11237 = ( x106 & ~n11142 ) | ( x106 & n11236 ) | ( ~n11142 & n11236 ) ;
  assign n11238 = ( x107 & ~n11139 ) | ( x107 & n11237 ) | ( ~n11139 & n11237 ) ;
  assign n11239 = ( x108 & ~n11136 ) | ( x108 & n11238 ) | ( ~n11136 & n11238 ) ;
  assign n11240 = ( x109 & ~n11133 ) | ( x109 & n11239 ) | ( ~n11133 & n11239 ) ;
  assign n11241 = ( x110 & ~n11130 ) | ( x110 & n11240 ) | ( ~n11130 & n11240 ) ;
  assign n11242 = ( x111 & ~n11127 ) | ( x111 & n11241 ) | ( ~n11127 & n11241 ) ;
  assign n11243 = ( x112 & ~n11124 ) | ( x112 & n11242 ) | ( ~n11124 & n11242 ) ;
  assign n11244 = ( x113 & ~n11121 ) | ( x113 & n11243 ) | ( ~n11121 & n11243 ) ;
  assign n11245 = ( x114 & ~n11118 ) | ( x114 & n11244 ) | ( ~n11118 & n11244 ) ;
  assign n11246 = ( x115 & ~n11115 ) | ( x115 & n11245 ) | ( ~n11115 & n11245 ) ;
  assign n11247 = ( x116 & ~n11112 ) | ( x116 & n11246 ) | ( ~n11112 & n11246 ) ;
  assign n11248 = ( x117 & ~n11109 ) | ( x117 & n11247 ) | ( ~n11109 & n11247 ) ;
  assign n11249 = ( x118 & ~n11106 ) | ( x118 & n11248 ) | ( ~n11106 & n11248 ) ;
  assign n11250 = ( x119 & ~n11088 ) | ( x119 & n11249 ) | ( ~n11088 & n11249 ) ;
  assign n11251 = ( x120 & ~n11059 ) | ( x120 & n11250 ) | ( ~n11059 & n11250 ) ;
  assign n11252 = ( x121 & ~n11103 ) | ( x121 & n11251 ) | ( ~n11103 & n11251 ) ;
  assign n11253 = ( ~x122 & n8330 ) | ( ~x122 & n11213 ) | ( n8330 & n11213 ) ;
  assign n11254 = ( n11230 & ~n11252 ) | ( n11230 & n11253 ) | ( ~n11252 & n11253 ) ;
  assign n11255 = n11252 | n11254 ;
  assign n11256 = ( ~n11213 & n11214 ) | ( ~n11213 & n11255 ) | ( n11214 & n11255 ) ;
  assign n11257 = n11250 ^ n11059 ^ x120 ;
  assign n11258 = n11256 ^ n11059 ^ 1'b0 ;
  assign n11259 = ( n11059 & n11257 ) | ( n11059 & ~n11258 ) | ( n11257 & ~n11258 ) ;
  assign n11260 = n11249 ^ n11088 ^ x119 ;
  assign n11261 = n11256 ^ n11088 ^ 1'b0 ;
  assign n11262 = ( n11088 & n11260 ) | ( n11088 & ~n11261 ) | ( n11260 & ~n11261 ) ;
  assign n11263 = n11247 ^ n11109 ^ x117 ;
  assign n11264 = n11256 ^ n11109 ^ 1'b0 ;
  assign n11265 = ( n11109 & n11263 ) | ( n11109 & ~n11264 ) | ( n11263 & ~n11264 ) ;
  assign n11266 = n11246 ^ n11112 ^ x116 ;
  assign n11267 = n11256 ^ n11112 ^ 1'b0 ;
  assign n11268 = n11245 ^ n11115 ^ x115 ;
  assign n11269 = n11256 ^ n11115 ^ 1'b0 ;
  assign n11270 = ( n11115 & n11268 ) | ( n11115 & ~n11269 ) | ( n11268 & ~n11269 ) ;
  assign n11271 = n11244 ^ n11118 ^ x114 ;
  assign n11272 = n11256 ^ n11118 ^ 1'b0 ;
  assign n11273 = ( n11118 & n11271 ) | ( n11118 & ~n11272 ) | ( n11271 & ~n11272 ) ;
  assign n11274 = n11256 ^ n11096 ^ 1'b0 ;
  assign n11275 = ( n11096 & n11220 ) | ( n11096 & ~n11274 ) | ( n11220 & ~n11274 ) ;
  assign n11276 = n11256 ^ n11098 ^ 1'b0 ;
  assign n11277 = ( n11098 & n11221 ) | ( n11098 & ~n11276 ) | ( n11221 & ~n11276 ) ;
  assign n11278 = n11256 ^ n11050 ^ 1'b0 ;
  assign n11279 = ( n11050 & n11222 ) | ( n11050 & ~n11278 ) | ( n11222 & ~n11278 ) ;
  assign n11280 = n11256 ^ n11055 ^ 1'b0 ;
  assign n11281 = ( n11055 & n11223 ) | ( n11055 & ~n11280 ) | ( n11223 & ~n11280 ) ;
  assign n11282 = n11256 ^ n11043 ^ 1'b0 ;
  assign n11283 = ( n11043 & n11224 ) | ( n11043 & ~n11282 ) | ( n11224 & ~n11282 ) ;
  assign n11284 = n11256 ^ n11049 ^ 1'b0 ;
  assign n11285 = ( n11049 & n11225 ) | ( n11049 & ~n11284 ) | ( n11225 & ~n11284 ) ;
  assign n11286 = n11256 ^ n11051 ^ 1'b0 ;
  assign n11287 = ( n11051 & n11226 ) | ( n11051 & ~n11286 ) | ( n11226 & ~n11286 ) ;
  assign n11288 = n11256 ^ n11044 ^ 1'b0 ;
  assign n11289 = ( n11044 & n11227 ) | ( n11044 & ~n11288 ) | ( n11227 & ~n11288 ) ;
  assign n11290 = n11256 ^ n11056 ^ 1'b0 ;
  assign n11291 = ( n11056 & n11228 ) | ( n11056 & ~n11290 ) | ( n11228 & ~n11290 ) ;
  assign n11292 = n11256 ^ n11041 ^ 1'b0 ;
  assign n11293 = ( n11041 & n11229 ) | ( n11041 & ~n11292 ) | ( n11229 & ~n11292 ) ;
  assign n11294 = ( n11112 & n11266 ) | ( n11112 & ~n11267 ) | ( n11266 & ~n11267 ) ;
  assign n11295 = n11256 ^ n11179 ^ 1'b0 ;
  assign n11296 = ( n11038 & n11179 ) | ( n11038 & n11295 ) | ( n11179 & n11295 ) ;
  assign n11297 = n11215 & n11255 ;
  assign n11298 = n11251 ^ n11103 ^ x121 ;
  assign n11299 = n11256 ^ n11103 ^ 1'b0 ;
  assign n11300 = ( n11103 & n11298 ) | ( n11103 & ~n11299 ) | ( n11298 & ~n11299 ) ;
  assign n11301 = n11248 ^ n11106 ^ x118 ;
  assign n11302 = n11256 ^ n11106 ^ 1'b0 ;
  assign n11303 = ( n11106 & n11301 ) | ( n11106 & ~n11302 ) | ( n11301 & ~n11302 ) ;
  assign n11304 = n11243 ^ n11121 ^ x113 ;
  assign n11305 = n11256 ^ n11121 ^ 1'b0 ;
  assign n11306 = ( n11121 & n11304 ) | ( n11121 & ~n11305 ) | ( n11304 & ~n11305 ) ;
  assign n11307 = n11212 ^ n11172 ^ x96 ;
  assign n11308 = n11256 ^ n11172 ^ 1'b0 ;
  assign n11309 = ( n11172 & n11307 ) | ( n11172 & ~n11308 ) | ( n11307 & ~n11308 ) ;
  assign n11310 = n11211 ^ n11175 ^ x95 ;
  assign n11311 = n11256 ^ n11175 ^ 1'b0 ;
  assign n11312 = ( n11175 & n11310 ) | ( n11175 & ~n11311 ) | ( n11310 & ~n11311 ) ;
  assign n11313 = n11209 ^ n11062 ^ x93 ;
  assign n11314 = n11256 ^ n11062 ^ 1'b0 ;
  assign n11315 = ( n11062 & n11313 ) | ( n11062 & ~n11314 ) | ( n11313 & ~n11314 ) ;
  assign n11316 = n11208 ^ n11064 ^ x92 ;
  assign n11317 = n11256 ^ n11064 ^ 1'b0 ;
  assign n11318 = ( n11064 & n11316 ) | ( n11064 & ~n11317 ) | ( n11316 & ~n11317 ) ;
  assign n11319 = n11207 ^ n11066 ^ x91 ;
  assign n11320 = n11256 ^ n11066 ^ 1'b0 ;
  assign n11321 = ( n11066 & n11319 ) | ( n11066 & ~n11320 ) | ( n11319 & ~n11320 ) ;
  assign n11322 = n11206 ^ n11068 ^ x90 ;
  assign n11323 = n11256 ^ n11068 ^ 1'b0 ;
  assign n11324 = ( n11068 & n11322 ) | ( n11068 & ~n11323 ) | ( n11322 & ~n11323 ) ;
  assign n11325 = n11204 ^ n11072 ^ x88 ;
  assign n11326 = n11256 ^ n11072 ^ 1'b0 ;
  assign n11327 = ( n11072 & n11325 ) | ( n11072 & ~n11326 ) | ( n11325 & ~n11326 ) ;
  assign n11328 = n11203 ^ n11074 ^ x87 ;
  assign n11329 = n11256 ^ n11074 ^ 1'b0 ;
  assign n11330 = ( n11074 & n11328 ) | ( n11074 & ~n11329 ) | ( n11328 & ~n11329 ) ;
  assign n11331 = n11201 ^ n11078 ^ x85 ;
  assign n11332 = n11256 ^ n11078 ^ 1'b0 ;
  assign n11333 = ( n11078 & n11331 ) | ( n11078 & ~n11332 ) | ( n11331 & ~n11332 ) ;
  assign n11334 = n11198 ^ n11082 ^ x83 ;
  assign n11335 = n11256 ^ n11082 ^ 1'b0 ;
  assign n11336 = ( n11082 & n11334 ) | ( n11082 & ~n11335 ) | ( n11334 & ~n11335 ) ;
  assign n11337 = n11197 ^ n11084 ^ x82 ;
  assign n11338 = n11256 ^ n11084 ^ 1'b0 ;
  assign n11339 = ( n11084 & n11337 ) | ( n11084 & ~n11338 ) | ( n11337 & ~n11338 ) ;
  assign n11340 = n11196 ^ n11086 ^ x81 ;
  assign n11341 = n11256 ^ n11086 ^ 1'b0 ;
  assign n11342 = ( n11086 & n11340 ) | ( n11086 & ~n11341 ) | ( n11340 & ~n11341 ) ;
  assign n11343 = n11195 ^ n11090 ^ x80 ;
  assign n11344 = n11256 ^ n11090 ^ 1'b0 ;
  assign n11345 = ( n11090 & n11343 ) | ( n11090 & ~n11344 ) | ( n11343 & ~n11344 ) ;
  assign n11346 = n11194 ^ n11092 ^ x79 ;
  assign n11347 = n11256 ^ n11092 ^ 1'b0 ;
  assign n11348 = ( n11092 & n11346 ) | ( n11092 & ~n11347 ) | ( n11346 & ~n11347 ) ;
  assign n11349 = n11193 ^ n11094 ^ x78 ;
  assign n11350 = n11256 ^ n11094 ^ 1'b0 ;
  assign n11351 = ( n11094 & n11349 ) | ( n11094 & ~n11350 ) | ( n11349 & ~n11350 ) ;
  assign n11352 = n11242 ^ n11124 ^ x112 ;
  assign n11353 = n11256 ^ n11124 ^ 1'b0 ;
  assign n11354 = ( n11124 & n11352 ) | ( n11124 & ~n11353 ) | ( n11352 & ~n11353 ) ;
  assign n11355 = n11241 ^ n11127 ^ x111 ;
  assign n11356 = n11256 ^ n11127 ^ 1'b0 ;
  assign n11357 = ( n11127 & n11355 ) | ( n11127 & ~n11356 ) | ( n11355 & ~n11356 ) ;
  assign n11358 = n11240 ^ n11130 ^ x110 ;
  assign n11359 = n11256 ^ n11130 ^ 1'b0 ;
  assign n11360 = ( n11130 & n11358 ) | ( n11130 & ~n11359 ) | ( n11358 & ~n11359 ) ;
  assign n11361 = n11239 ^ n11133 ^ x109 ;
  assign n11362 = n11256 ^ n11133 ^ 1'b0 ;
  assign n11363 = ( n11133 & n11361 ) | ( n11133 & ~n11362 ) | ( n11361 & ~n11362 ) ;
  assign n11364 = n11238 ^ n11136 ^ x108 ;
  assign n11365 = n11256 ^ n11136 ^ 1'b0 ;
  assign n11366 = ( n11136 & n11364 ) | ( n11136 & ~n11365 ) | ( n11364 & ~n11365 ) ;
  assign n11367 = n11237 ^ n11139 ^ x107 ;
  assign n11368 = n11256 ^ n11139 ^ 1'b0 ;
  assign n11369 = ( n11139 & n11367 ) | ( n11139 & ~n11368 ) | ( n11367 & ~n11368 ) ;
  assign n11370 = n11235 ^ n11145 ^ x105 ;
  assign n11371 = n11256 ^ n11145 ^ 1'b0 ;
  assign n11372 = ( n11145 & n11370 ) | ( n11145 & ~n11371 ) | ( n11370 & ~n11371 ) ;
  assign n11373 = n11234 ^ n11148 ^ x104 ;
  assign n11374 = n11256 ^ n11148 ^ 1'b0 ;
  assign n11375 = ( n11148 & n11373 ) | ( n11148 & ~n11374 ) | ( n11373 & ~n11374 ) ;
  assign n11376 = n11233 ^ n11151 ^ x103 ;
  assign n11377 = n11256 ^ n11151 ^ 1'b0 ;
  assign n11378 = ( n11151 & n11376 ) | ( n11151 & ~n11377 ) | ( n11376 & ~n11377 ) ;
  assign n11379 = n11232 ^ n11154 ^ x102 ;
  assign n11380 = n11256 ^ n11154 ^ 1'b0 ;
  assign n11381 = ( n11154 & n11379 ) | ( n11154 & ~n11380 ) | ( n11379 & ~n11380 ) ;
  assign n11382 = n11231 ^ n11157 ^ x101 ;
  assign n11383 = n11256 ^ n11157 ^ 1'b0 ;
  assign n11384 = ( n11157 & n11382 ) | ( n11157 & ~n11383 ) | ( n11382 & ~n11383 ) ;
  assign n11385 = n11219 ^ n11160 ^ x100 ;
  assign n11386 = n11256 ^ n11160 ^ 1'b0 ;
  assign n11387 = ( n11160 & n11385 ) | ( n11160 & ~n11386 ) | ( n11385 & ~n11386 ) ;
  assign n11388 = n11218 ^ n11163 ^ x99 ;
  assign n11389 = n11256 ^ n11163 ^ 1'b0 ;
  assign n11390 = ( n11163 & n11388 ) | ( n11163 & ~n11389 ) | ( n11388 & ~n11389 ) ;
  assign n11391 = n11217 ^ n11166 ^ x98 ;
  assign n11392 = n11256 ^ n11166 ^ 1'b0 ;
  assign n11393 = ( n11166 & n11391 ) | ( n11166 & ~n11392 ) | ( n11391 & ~n11392 ) ;
  assign n11394 = n11216 ^ n11169 ^ x97 ;
  assign n11395 = n11256 ^ n11169 ^ 1'b0 ;
  assign n11396 = ( n11169 & n11394 ) | ( n11169 & ~n11395 ) | ( n11394 & ~n11395 ) ;
  assign n11397 = n11236 ^ n11142 ^ x106 ;
  assign n11398 = n11256 ^ n11142 ^ 1'b0 ;
  assign n11399 = ( n11142 & n11397 ) | ( n11142 & ~n11398 ) | ( n11397 & ~n11398 ) ;
  assign n11400 = n11210 ^ n11178 ^ x94 ;
  assign n11401 = n11256 ^ n11178 ^ 1'b0 ;
  assign n11402 = ( n11178 & n11400 ) | ( n11178 & ~n11401 ) | ( n11400 & ~n11401 ) ;
  assign n11403 = n11205 ^ n11070 ^ x89 ;
  assign n11404 = n11256 ^ n11070 ^ 1'b0 ;
  assign n11405 = ( n11070 & n11403 ) | ( n11070 & ~n11404 ) | ( n11403 & ~n11404 ) ;
  assign n11406 = n11202 ^ n11076 ^ x86 ;
  assign n11407 = n11256 ^ n11076 ^ 1'b0 ;
  assign n11408 = ( n11076 & n11406 ) | ( n11076 & ~n11407 ) | ( n11406 & ~n11407 ) ;
  assign n11409 = n11199 ^ n11080 ^ x84 ;
  assign n11410 = n11256 ^ n11080 ^ 1'b0 ;
  assign n11411 = ( n11080 & n11409 ) | ( n11080 & ~n11410 ) | ( n11409 & ~n11410 ) ;
  assign n11412 = n11183 ^ n11052 ^ x68 ;
  assign n11413 = n11256 ^ n11052 ^ 1'b0 ;
  assign n11414 = ( n11052 & n11412 ) | ( n11052 & ~n11413 ) | ( n11412 & ~n11413 ) ;
  assign n11415 = n11256 ^ n11181 ^ 1'b0 ;
  assign n11416 = ( n11100 & n11181 ) | ( n11100 & n11415 ) | ( n11181 & n11415 ) ;
  assign n11417 = x64 & n11256 ;
  assign n11418 = n11417 ^ x64 ^ x5 ;
  assign n11419 = n11418 ^ n8575 ^ x65 ;
  assign n11420 = ( x65 & n8575 ) | ( x65 & n11419 ) | ( n8575 & n11419 ) ;
  assign n11421 = n11420 ^ n11296 ^ x66 ;
  assign n11422 = ( x66 & n11420 ) | ( x66 & n11421 ) | ( n11420 & n11421 ) ;
  assign n11423 = ( x67 & ~n11416 ) | ( x67 & n11422 ) | ( ~n11416 & n11422 ) ;
  assign n11424 = ( x68 & ~n11293 ) | ( x68 & n11423 ) | ( ~n11293 & n11423 ) ;
  assign n11425 = ( x69 & ~n11414 ) | ( x69 & n11424 ) | ( ~n11414 & n11424 ) ;
  assign n11426 = ( x70 & ~n11291 ) | ( x70 & n11425 ) | ( ~n11291 & n11425 ) ;
  assign n11427 = n322 | n11297 ;
  assign n11428 = ( x123 & n154 ) | ( x123 & ~n11297 ) | ( n154 & ~n11297 ) ;
  assign n11429 = n8330 & n11427 ;
  assign n11430 = n11425 ^ n11291 ^ x70 ;
  assign n11431 = n11424 ^ n11414 ^ x69 ;
  assign n11432 = n11423 ^ n11293 ^ x68 ;
  assign n11433 = n11422 ^ n11416 ^ x67 ;
  assign n11434 = ( x71 & ~n11289 ) | ( x71 & n11426 ) | ( ~n11289 & n11426 ) ;
  assign n11435 = ( x72 & ~n11287 ) | ( x72 & n11434 ) | ( ~n11287 & n11434 ) ;
  assign n11436 = ( x73 & ~n11285 ) | ( x73 & n11435 ) | ( ~n11285 & n11435 ) ;
  assign n11437 = ( x74 & ~n11283 ) | ( x74 & n11436 ) | ( ~n11283 & n11436 ) ;
  assign n11438 = ( x75 & ~n11281 ) | ( x75 & n11437 ) | ( ~n11281 & n11437 ) ;
  assign n11439 = ( x76 & ~n11279 ) | ( x76 & n11438 ) | ( ~n11279 & n11438 ) ;
  assign n11440 = ( x77 & ~n11277 ) | ( x77 & n11439 ) | ( ~n11277 & n11439 ) ;
  assign n11441 = ( x78 & ~n11275 ) | ( x78 & n11440 ) | ( ~n11275 & n11440 ) ;
  assign n11442 = ( x79 & ~n11351 ) | ( x79 & n11441 ) | ( ~n11351 & n11441 ) ;
  assign n11443 = ( x80 & ~n11348 ) | ( x80 & n11442 ) | ( ~n11348 & n11442 ) ;
  assign n11444 = ( x81 & ~n11345 ) | ( x81 & n11443 ) | ( ~n11345 & n11443 ) ;
  assign n11445 = ( x82 & ~n11342 ) | ( x82 & n11444 ) | ( ~n11342 & n11444 ) ;
  assign n11446 = ( x83 & ~n11339 ) | ( x83 & n11445 ) | ( ~n11339 & n11445 ) ;
  assign n11447 = ( x84 & ~n11336 ) | ( x84 & n11446 ) | ( ~n11336 & n11446 ) ;
  assign n11448 = ( x85 & ~n11411 ) | ( x85 & n11447 ) | ( ~n11411 & n11447 ) ;
  assign n11449 = ( x86 & ~n11333 ) | ( x86 & n11448 ) | ( ~n11333 & n11448 ) ;
  assign n11450 = ( x87 & ~n11408 ) | ( x87 & n11449 ) | ( ~n11408 & n11449 ) ;
  assign n11451 = ( x88 & ~n11330 ) | ( x88 & n11450 ) | ( ~n11330 & n11450 ) ;
  assign n11452 = ( x89 & ~n11327 ) | ( x89 & n11451 ) | ( ~n11327 & n11451 ) ;
  assign n11453 = ( x90 & ~n11405 ) | ( x90 & n11452 ) | ( ~n11405 & n11452 ) ;
  assign n11454 = ( x91 & ~n11324 ) | ( x91 & n11453 ) | ( ~n11324 & n11453 ) ;
  assign n11455 = ( x92 & ~n11321 ) | ( x92 & n11454 ) | ( ~n11321 & n11454 ) ;
  assign n11456 = ( x93 & ~n11318 ) | ( x93 & n11455 ) | ( ~n11318 & n11455 ) ;
  assign n11457 = ( x94 & ~n11315 ) | ( x94 & n11456 ) | ( ~n11315 & n11456 ) ;
  assign n11458 = ( x95 & ~n11402 ) | ( x95 & n11457 ) | ( ~n11402 & n11457 ) ;
  assign n11459 = ( x96 & ~n11312 ) | ( x96 & n11458 ) | ( ~n11312 & n11458 ) ;
  assign n11460 = ( x97 & ~n11309 ) | ( x97 & n11459 ) | ( ~n11309 & n11459 ) ;
  assign n11461 = ( x98 & ~n11396 ) | ( x98 & n11460 ) | ( ~n11396 & n11460 ) ;
  assign n11462 = ( x99 & ~n11393 ) | ( x99 & n11461 ) | ( ~n11393 & n11461 ) ;
  assign n11463 = ( x100 & ~n11390 ) | ( x100 & n11462 ) | ( ~n11390 & n11462 ) ;
  assign n11464 = ( x101 & ~n11387 ) | ( x101 & n11463 ) | ( ~n11387 & n11463 ) ;
  assign n11465 = ( x102 & ~n11384 ) | ( x102 & n11464 ) | ( ~n11384 & n11464 ) ;
  assign n11466 = ( x103 & ~n11381 ) | ( x103 & n11465 ) | ( ~n11381 & n11465 ) ;
  assign n11467 = ( x104 & ~n11378 ) | ( x104 & n11466 ) | ( ~n11378 & n11466 ) ;
  assign n11468 = ( x105 & ~n11375 ) | ( x105 & n11467 ) | ( ~n11375 & n11467 ) ;
  assign n11469 = n11452 ^ n11405 ^ x90 ;
  assign n11470 = n11448 ^ n11333 ^ x86 ;
  assign n11471 = n11437 ^ n11281 ^ x75 ;
  assign n11472 = n11435 ^ n11285 ^ x73 ;
  assign n11473 = n11466 ^ n11378 ^ x104 ;
  assign n11474 = n11434 ^ n11287 ^ x72 ;
  assign n11475 = n11426 ^ n11289 ^ x71 ;
  assign n11476 = n11468 ^ n11372 ^ x106 ;
  assign n11477 = n11467 ^ n11375 ^ x105 ;
  assign n11478 = ( x106 & ~n11372 ) | ( x106 & n11468 ) | ( ~n11372 & n11468 ) ;
  assign n11479 = ( x107 & ~n11399 ) | ( x107 & n11478 ) | ( ~n11399 & n11478 ) ;
  assign n11480 = ( x108 & ~n11369 ) | ( x108 & n11479 ) | ( ~n11369 & n11479 ) ;
  assign n11481 = ( x109 & ~n11366 ) | ( x109 & n11480 ) | ( ~n11366 & n11480 ) ;
  assign n11482 = ( x110 & ~n11363 ) | ( x110 & n11481 ) | ( ~n11363 & n11481 ) ;
  assign n11483 = ( x111 & ~n11360 ) | ( x111 & n11482 ) | ( ~n11360 & n11482 ) ;
  assign n11484 = ( x112 & ~n11357 ) | ( x112 & n11483 ) | ( ~n11357 & n11483 ) ;
  assign n11485 = ( x113 & ~n11354 ) | ( x113 & n11484 ) | ( ~n11354 & n11484 ) ;
  assign n11486 = ( x114 & ~n11306 ) | ( x114 & n11485 ) | ( ~n11306 & n11485 ) ;
  assign n11487 = ( x115 & ~n11273 ) | ( x115 & n11486 ) | ( ~n11273 & n11486 ) ;
  assign n11488 = ( x116 & ~n11270 ) | ( x116 & n11487 ) | ( ~n11270 & n11487 ) ;
  assign n11489 = ( x117 & ~n11294 ) | ( x117 & n11488 ) | ( ~n11294 & n11488 ) ;
  assign n11490 = ( x118 & ~n11265 ) | ( x118 & n11489 ) | ( ~n11265 & n11489 ) ;
  assign n11491 = ( x119 & ~n11303 ) | ( x119 & n11490 ) | ( ~n11303 & n11490 ) ;
  assign n11492 = ( x120 & ~n11262 ) | ( x120 & n11491 ) | ( ~n11262 & n11491 ) ;
  assign n11493 = ( x121 & ~n11259 ) | ( x121 & n11492 ) | ( ~n11259 & n11492 ) ;
  assign n11494 = ( x122 & ~n11300 ) | ( x122 & n11493 ) | ( ~n11300 & n11493 ) ;
  assign n11495 = ( ~x123 & n154 ) | ( ~x123 & n11427 ) | ( n154 & n11427 ) ;
  assign n11496 = ( n11428 & ~n11494 ) | ( n11428 & n11495 ) | ( ~n11494 & n11495 ) ;
  assign n11497 = n11494 | n11496 ;
  assign n11498 = ( ~n11427 & n11429 ) | ( ~n11427 & n11497 ) | ( n11429 & n11497 ) ;
  assign n11499 = n11492 ^ n11259 ^ x121 ;
  assign n11500 = n11498 ^ n11259 ^ 1'b0 ;
  assign n11501 = ( n11259 & n11499 ) | ( n11259 & ~n11500 ) | ( n11499 & ~n11500 ) ;
  assign n11502 = n11498 ^ n11372 ^ 1'b0 ;
  assign n11503 = ( n11372 & n11476 ) | ( n11372 & ~n11502 ) | ( n11476 & ~n11502 ) ;
  assign n11504 = n11498 ^ n11375 ^ 1'b0 ;
  assign n11505 = n11498 ^ n11378 ^ 1'b0 ;
  assign n11506 = ( n11378 & n11473 ) | ( n11378 & ~n11505 ) | ( n11473 & ~n11505 ) ;
  assign n11507 = n11498 ^ n11405 ^ 1'b0 ;
  assign n11508 = ( n11405 & n11469 ) | ( n11405 & ~n11507 ) | ( n11469 & ~n11507 ) ;
  assign n11509 = n11498 ^ n11333 ^ 1'b0 ;
  assign n11510 = ( n11333 & n11470 ) | ( n11333 & ~n11509 ) | ( n11470 & ~n11509 ) ;
  assign n11511 = n11498 ^ n11281 ^ 1'b0 ;
  assign n11512 = ( n11281 & n11471 ) | ( n11281 & ~n11511 ) | ( n11471 & ~n11511 ) ;
  assign n11513 = n11498 ^ n11285 ^ 1'b0 ;
  assign n11514 = ( n11285 & n11472 ) | ( n11285 & ~n11513 ) | ( n11472 & ~n11513 ) ;
  assign n11515 = ( n11375 & n11477 ) | ( n11375 & ~n11504 ) | ( n11477 & ~n11504 ) ;
  assign n11516 = n11498 ^ n11287 ^ 1'b0 ;
  assign n11517 = ( n11287 & n11474 ) | ( n11287 & ~n11516 ) | ( n11474 & ~n11516 ) ;
  assign n11518 = n11498 ^ n11289 ^ 1'b0 ;
  assign n11519 = ( n11289 & n11475 ) | ( n11289 & ~n11518 ) | ( n11475 & ~n11518 ) ;
  assign n11520 = n11498 ^ n11291 ^ 1'b0 ;
  assign n11521 = ( n11291 & n11430 ) | ( n11291 & ~n11520 ) | ( n11430 & ~n11520 ) ;
  assign n11522 = n11498 ^ n11414 ^ 1'b0 ;
  assign n11523 = ( n11414 & n11431 ) | ( n11414 & ~n11522 ) | ( n11431 & ~n11522 ) ;
  assign n11524 = n11498 ^ n11293 ^ 1'b0 ;
  assign n11525 = ( n11293 & n11432 ) | ( n11293 & ~n11524 ) | ( n11432 & ~n11524 ) ;
  assign n11526 = n11498 ^ n11416 ^ 1'b0 ;
  assign n11527 = ( n11416 & n11433 ) | ( n11416 & ~n11526 ) | ( n11433 & ~n11526 ) ;
  assign n11528 = n11498 ^ n11421 ^ 1'b0 ;
  assign n11529 = ( n11296 & n11421 ) | ( n11296 & n11528 ) | ( n11421 & n11528 ) ;
  assign n11530 = n11498 ^ n11419 ^ 1'b0 ;
  assign n11531 = ( n11418 & n11419 ) | ( n11418 & n11530 ) | ( n11419 & n11530 ) ;
  assign n11532 = n11429 & n11497 ;
  assign n11533 = n11493 ^ n11300 ^ x122 ;
  assign n11534 = n11498 ^ n11300 ^ 1'b0 ;
  assign n11535 = ( n11300 & n11533 ) | ( n11300 & ~n11534 ) | ( n11533 & ~n11534 ) ;
  assign n11536 = n11491 ^ n11262 ^ x120 ;
  assign n11537 = n11498 ^ n11262 ^ 1'b0 ;
  assign n11538 = ( n11262 & n11536 ) | ( n11262 & ~n11537 ) | ( n11536 & ~n11537 ) ;
  assign n11539 = n11490 ^ n11303 ^ x119 ;
  assign n11540 = n11498 ^ n11303 ^ 1'b0 ;
  assign n11541 = ( n11303 & n11539 ) | ( n11303 & ~n11540 ) | ( n11539 & ~n11540 ) ;
  assign n11542 = n11489 ^ n11265 ^ x118 ;
  assign n11543 = n11498 ^ n11265 ^ 1'b0 ;
  assign n11544 = ( n11265 & n11542 ) | ( n11265 & ~n11543 ) | ( n11542 & ~n11543 ) ;
  assign n11545 = n11488 ^ n11294 ^ x117 ;
  assign n11546 = n11498 ^ n11294 ^ 1'b0 ;
  assign n11547 = ( n11294 & n11545 ) | ( n11294 & ~n11546 ) | ( n11545 & ~n11546 ) ;
  assign n11548 = n11487 ^ n11270 ^ x116 ;
  assign n11549 = n11498 ^ n11270 ^ 1'b0 ;
  assign n11550 = ( n11270 & n11548 ) | ( n11270 & ~n11549 ) | ( n11548 & ~n11549 ) ;
  assign n11551 = n11486 ^ n11273 ^ x115 ;
  assign n11552 = n11498 ^ n11273 ^ 1'b0 ;
  assign n11553 = ( n11273 & n11551 ) | ( n11273 & ~n11552 ) | ( n11551 & ~n11552 ) ;
  assign n11554 = n11485 ^ n11306 ^ x114 ;
  assign n11555 = n11498 ^ n11306 ^ 1'b0 ;
  assign n11556 = ( n11306 & n11554 ) | ( n11306 & ~n11555 ) | ( n11554 & ~n11555 ) ;
  assign n11557 = n11484 ^ n11354 ^ x113 ;
  assign n11558 = n11498 ^ n11354 ^ 1'b0 ;
  assign n11559 = ( n11354 & n11557 ) | ( n11354 & ~n11558 ) | ( n11557 & ~n11558 ) ;
  assign n11560 = n11483 ^ n11357 ^ x112 ;
  assign n11561 = n11498 ^ n11357 ^ 1'b0 ;
  assign n11562 = ( n11357 & n11560 ) | ( n11357 & ~n11561 ) | ( n11560 & ~n11561 ) ;
  assign n11563 = n11482 ^ n11360 ^ x111 ;
  assign n11564 = n11498 ^ n11360 ^ 1'b0 ;
  assign n11565 = ( n11360 & n11563 ) | ( n11360 & ~n11564 ) | ( n11563 & ~n11564 ) ;
  assign n11566 = n11481 ^ n11363 ^ x110 ;
  assign n11567 = n11498 ^ n11363 ^ 1'b0 ;
  assign n11568 = ( n11363 & n11566 ) | ( n11363 & ~n11567 ) | ( n11566 & ~n11567 ) ;
  assign n11569 = n11480 ^ n11366 ^ x109 ;
  assign n11570 = n11498 ^ n11366 ^ 1'b0 ;
  assign n11571 = ( n11366 & n11569 ) | ( n11366 & ~n11570 ) | ( n11569 & ~n11570 ) ;
  assign n11572 = n11479 ^ n11369 ^ x108 ;
  assign n11573 = n11498 ^ n11369 ^ 1'b0 ;
  assign n11574 = ( n11369 & n11572 ) | ( n11369 & ~n11573 ) | ( n11572 & ~n11573 ) ;
  assign n11575 = n11478 ^ n11399 ^ x107 ;
  assign n11576 = n11498 ^ n11399 ^ 1'b0 ;
  assign n11577 = ( n11399 & n11575 ) | ( n11399 & ~n11576 ) | ( n11575 & ~n11576 ) ;
  assign n11578 = n11465 ^ n11381 ^ x103 ;
  assign n11579 = n11498 ^ n11381 ^ 1'b0 ;
  assign n11580 = ( n11381 & n11578 ) | ( n11381 & ~n11579 ) | ( n11578 & ~n11579 ) ;
  assign n11581 = n11450 ^ n11330 ^ x88 ;
  assign n11582 = n11498 ^ n11330 ^ 1'b0 ;
  assign n11583 = ( n11330 & n11581 ) | ( n11330 & ~n11582 ) | ( n11581 & ~n11582 ) ;
  assign n11584 = n11449 ^ n11408 ^ x87 ;
  assign n11585 = n11498 ^ n11408 ^ 1'b0 ;
  assign n11586 = ( n11408 & n11584 ) | ( n11408 & ~n11585 ) | ( n11584 & ~n11585 ) ;
  assign n11587 = n11447 ^ n11411 ^ x85 ;
  assign n11588 = n11498 ^ n11411 ^ 1'b0 ;
  assign n11589 = ( n11411 & n11587 ) | ( n11411 & ~n11588 ) | ( n11587 & ~n11588 ) ;
  assign n11590 = n11446 ^ n11336 ^ x84 ;
  assign n11591 = n11498 ^ n11336 ^ 1'b0 ;
  assign n11592 = ( n11336 & n11590 ) | ( n11336 & ~n11591 ) | ( n11590 & ~n11591 ) ;
  assign n11593 = n11445 ^ n11339 ^ x83 ;
  assign n11594 = n11498 ^ n11339 ^ 1'b0 ;
  assign n11595 = ( n11339 & n11593 ) | ( n11339 & ~n11594 ) | ( n11593 & ~n11594 ) ;
  assign n11596 = n11444 ^ n11342 ^ x82 ;
  assign n11597 = n11498 ^ n11342 ^ 1'b0 ;
  assign n11598 = ( n11342 & n11596 ) | ( n11342 & ~n11597 ) | ( n11596 & ~n11597 ) ;
  assign n11599 = n11443 ^ n11345 ^ x81 ;
  assign n11600 = n11498 ^ n11345 ^ 1'b0 ;
  assign n11601 = ( n11345 & n11599 ) | ( n11345 & ~n11600 ) | ( n11599 & ~n11600 ) ;
  assign n11602 = n11442 ^ n11348 ^ x80 ;
  assign n11603 = n11498 ^ n11348 ^ 1'b0 ;
  assign n11604 = ( n11348 & n11602 ) | ( n11348 & ~n11603 ) | ( n11602 & ~n11603 ) ;
  assign n11605 = n11441 ^ n11351 ^ x79 ;
  assign n11606 = n11498 ^ n11351 ^ 1'b0 ;
  assign n11607 = ( n11351 & n11605 ) | ( n11351 & ~n11606 ) | ( n11605 & ~n11606 ) ;
  assign n11608 = n11440 ^ n11275 ^ x78 ;
  assign n11609 = n11498 ^ n11275 ^ 1'b0 ;
  assign n11610 = ( n11275 & n11608 ) | ( n11275 & ~n11609 ) | ( n11608 & ~n11609 ) ;
  assign n11611 = n11439 ^ n11277 ^ x77 ;
  assign n11612 = n11498 ^ n11277 ^ 1'b0 ;
  assign n11613 = ( n11277 & n11611 ) | ( n11277 & ~n11612 ) | ( n11611 & ~n11612 ) ;
  assign n11614 = n11438 ^ n11279 ^ x76 ;
  assign n11615 = n11498 ^ n11279 ^ 1'b0 ;
  assign n11616 = ( n11279 & n11614 ) | ( n11279 & ~n11615 ) | ( n11614 & ~n11615 ) ;
  assign n11617 = n11436 ^ n11283 ^ x74 ;
  assign n11618 = n11498 ^ n11283 ^ 1'b0 ;
  assign n11619 = ( n11283 & n11617 ) | ( n11283 & ~n11618 ) | ( n11617 & ~n11618 ) ;
  assign n11620 = n11464 ^ n11384 ^ x102 ;
  assign n11621 = n11498 ^ n11384 ^ 1'b0 ;
  assign n11622 = ( n11384 & n11620 ) | ( n11384 & ~n11621 ) | ( n11620 & ~n11621 ) ;
  assign n11623 = n11463 ^ n11387 ^ x101 ;
  assign n11624 = n11498 ^ n11387 ^ 1'b0 ;
  assign n11625 = ( n11387 & n11623 ) | ( n11387 & ~n11624 ) | ( n11623 & ~n11624 ) ;
  assign n11626 = n11462 ^ n11390 ^ x100 ;
  assign n11627 = n11498 ^ n11390 ^ 1'b0 ;
  assign n11628 = ( n11390 & n11626 ) | ( n11390 & ~n11627 ) | ( n11626 & ~n11627 ) ;
  assign n11629 = n11461 ^ n11393 ^ x99 ;
  assign n11630 = n11498 ^ n11393 ^ 1'b0 ;
  assign n11631 = ( n11393 & n11629 ) | ( n11393 & ~n11630 ) | ( n11629 & ~n11630 ) ;
  assign n11632 = n11460 ^ n11396 ^ x98 ;
  assign n11633 = n11498 ^ n11396 ^ 1'b0 ;
  assign n11634 = ( n11396 & n11632 ) | ( n11396 & ~n11633 ) | ( n11632 & ~n11633 ) ;
  assign n11635 = n11459 ^ n11309 ^ x97 ;
  assign n11636 = n11498 ^ n11309 ^ 1'b0 ;
  assign n11637 = ( n11309 & n11635 ) | ( n11309 & ~n11636 ) | ( n11635 & ~n11636 ) ;
  assign n11638 = n11458 ^ n11312 ^ x96 ;
  assign n11639 = n11498 ^ n11312 ^ 1'b0 ;
  assign n11640 = ( n11312 & n11638 ) | ( n11312 & ~n11639 ) | ( n11638 & ~n11639 ) ;
  assign n11641 = n11457 ^ n11402 ^ x95 ;
  assign n11642 = n11498 ^ n11402 ^ 1'b0 ;
  assign n11643 = ( n11402 & n11641 ) | ( n11402 & ~n11642 ) | ( n11641 & ~n11642 ) ;
  assign n11644 = n11456 ^ n11315 ^ x94 ;
  assign n11645 = n11498 ^ n11315 ^ 1'b0 ;
  assign n11646 = ( n11315 & n11644 ) | ( n11315 & ~n11645 ) | ( n11644 & ~n11645 ) ;
  assign n11647 = n11455 ^ n11318 ^ x93 ;
  assign n11648 = n11498 ^ n11318 ^ 1'b0 ;
  assign n11649 = ( n11318 & n11647 ) | ( n11318 & ~n11648 ) | ( n11647 & ~n11648 ) ;
  assign n11650 = n11454 ^ n11321 ^ x92 ;
  assign n11651 = n11498 ^ n11321 ^ 1'b0 ;
  assign n11652 = ( n11321 & n11650 ) | ( n11321 & ~n11651 ) | ( n11650 & ~n11651 ) ;
  assign n11653 = n11453 ^ n11324 ^ x91 ;
  assign n11654 = n11498 ^ n11324 ^ 1'b0 ;
  assign n11655 = ( n11324 & n11653 ) | ( n11324 & ~n11654 ) | ( n11653 & ~n11654 ) ;
  assign n11656 = n11451 ^ n11327 ^ x89 ;
  assign n11657 = n11498 ^ n11327 ^ 1'b0 ;
  assign n11658 = ( n11327 & n11656 ) | ( n11327 & ~n11657 ) | ( n11656 & ~n11657 ) ;
  assign n11659 = x64 & n11498 ;
  assign n11660 = n11659 ^ x64 ^ x4 ;
  assign n11661 = n11660 ^ n8817 ^ x65 ;
  assign n11662 = ( x65 & n8817 ) | ( x65 & n11661 ) | ( n8817 & n11661 ) ;
  assign n11663 = n11662 ^ n11531 ^ x66 ;
  assign n11664 = ( x66 & n11662 ) | ( x66 & n11663 ) | ( n11662 & n11663 ) ;
  assign n11665 = ( x67 & ~n11529 ) | ( x67 & n11664 ) | ( ~n11529 & n11664 ) ;
  assign n11666 = ( x68 & ~n11527 ) | ( x68 & n11665 ) | ( ~n11527 & n11665 ) ;
  assign n11667 = ( x69 & ~n11525 ) | ( x69 & n11666 ) | ( ~n11525 & n11666 ) ;
  assign n11668 = ( x70 & ~n11523 ) | ( x70 & n11667 ) | ( ~n11523 & n11667 ) ;
  assign n11669 = ( x71 & ~n11521 ) | ( x71 & n11668 ) | ( ~n11521 & n11668 ) ;
  assign n11670 = ( x72 & ~n11519 ) | ( x72 & n11669 ) | ( ~n11519 & n11669 ) ;
  assign n11671 = ( x73 & ~n11517 ) | ( x73 & n11670 ) | ( ~n11517 & n11670 ) ;
  assign n11672 = ( x74 & ~n11514 ) | ( x74 & n11671 ) | ( ~n11514 & n11671 ) ;
  assign n11673 = ( x75 & ~n11619 ) | ( x75 & n11672 ) | ( ~n11619 & n11672 ) ;
  assign n11674 = ( x76 & ~n11512 ) | ( x76 & n11673 ) | ( ~n11512 & n11673 ) ;
  assign n11675 = ( x77 & ~n11616 ) | ( x77 & n11674 ) | ( ~n11616 & n11674 ) ;
  assign n11676 = ( x78 & ~n11613 ) | ( x78 & n11675 ) | ( ~n11613 & n11675 ) ;
  assign n11677 = ( x79 & ~n11610 ) | ( x79 & n11676 ) | ( ~n11610 & n11676 ) ;
  assign n11678 = ( x80 & ~n11607 ) | ( x80 & n11677 ) | ( ~n11607 & n11677 ) ;
  assign n11679 = ( x81 & ~n11604 ) | ( x81 & n11678 ) | ( ~n11604 & n11678 ) ;
  assign n11680 = ( x82 & ~n11601 ) | ( x82 & n11679 ) | ( ~n11601 & n11679 ) ;
  assign n11681 = n322 | n11532 ;
  assign n11682 = ( x83 & ~n11598 ) | ( x83 & n11680 ) | ( ~n11598 & n11680 ) ;
  assign n11683 = ( x84 & ~n11595 ) | ( x84 & n11682 ) | ( ~n11595 & n11682 ) ;
  assign n11684 = ( x85 & ~n11592 ) | ( x85 & n11683 ) | ( ~n11592 & n11683 ) ;
  assign n11685 = ( x86 & ~n11589 ) | ( x86 & n11684 ) | ( ~n11589 & n11684 ) ;
  assign n11686 = ( x87 & ~n11510 ) | ( x87 & n11685 ) | ( ~n11510 & n11685 ) ;
  assign n11687 = ( x88 & ~n11586 ) | ( x88 & n11686 ) | ( ~n11586 & n11686 ) ;
  assign n11688 = n11675 ^ n11613 ^ x78 ;
  assign n11689 = ( x89 & ~n11583 ) | ( x89 & n11687 ) | ( ~n11583 & n11687 ) ;
  assign n11690 = ( x90 & ~n11658 ) | ( x90 & n11689 ) | ( ~n11658 & n11689 ) ;
  assign n11691 = ( x91 & ~n11508 ) | ( x91 & n11690 ) | ( ~n11508 & n11690 ) ;
  assign n11692 = ( x92 & ~n11655 ) | ( x92 & n11691 ) | ( ~n11655 & n11691 ) ;
  assign n11693 = ( x93 & ~n11652 ) | ( x93 & n11692 ) | ( ~n11652 & n11692 ) ;
  assign n11694 = ( x94 & ~n11649 ) | ( x94 & n11693 ) | ( ~n11649 & n11693 ) ;
  assign n11695 = n154 & n11681 ;
  assign n11696 = n11664 ^ n11529 ^ x67 ;
  assign n11697 = n11665 ^ n11527 ^ x68 ;
  assign n11698 = n11666 ^ n11525 ^ x69 ;
  assign n11699 = n11667 ^ n11523 ^ x70 ;
  assign n11700 = n11668 ^ n11521 ^ x71 ;
  assign n11701 = n11669 ^ n11519 ^ x72 ;
  assign n11702 = n11670 ^ n11517 ^ x73 ;
  assign n11703 = n11671 ^ n11514 ^ x74 ;
  assign n11704 = n11672 ^ n11619 ^ x75 ;
  assign n11705 = n11673 ^ n11512 ^ x76 ;
  assign n11706 = n11674 ^ n11616 ^ x77 ;
  assign n11707 = n11694 ^ n11646 ^ x95 ;
  assign n11708 = n11676 ^ n11610 ^ x79 ;
  assign n11709 = n11677 ^ n11607 ^ x80 ;
  assign n11710 = n11678 ^ n11604 ^ x81 ;
  assign n11711 = n11679 ^ n11601 ^ x82 ;
  assign n11712 = n11680 ^ n11598 ^ x83 ;
  assign n11713 = n11682 ^ n11595 ^ x84 ;
  assign n11714 = n11683 ^ n11592 ^ x85 ;
  assign n11715 = n11684 ^ n11589 ^ x86 ;
  assign n11716 = n11685 ^ n11510 ^ x87 ;
  assign n11717 = n11686 ^ n11586 ^ x88 ;
  assign n11718 = n11687 ^ n11583 ^ x89 ;
  assign n11719 = n11689 ^ n11658 ^ x90 ;
  assign n11720 = n11690 ^ n11508 ^ x91 ;
  assign n11721 = n11691 ^ n11655 ^ x92 ;
  assign n11722 = n11692 ^ n11652 ^ x93 ;
  assign n11723 = ( x95 & ~n11646 ) | ( x95 & n11694 ) | ( ~n11646 & n11694 ) ;
  assign n11724 = ( x124 & n153 ) | ( x124 & ~n11532 ) | ( n153 & ~n11532 ) ;
  assign n11725 = n11693 ^ n11649 ^ x94 ;
  assign n11726 = ( x96 & ~n11643 ) | ( x96 & n11723 ) | ( ~n11643 & n11723 ) ;
  assign n11727 = ( x97 & ~n11640 ) | ( x97 & n11726 ) | ( ~n11640 & n11726 ) ;
  assign n11728 = ( x98 & ~n11637 ) | ( x98 & n11727 ) | ( ~n11637 & n11727 ) ;
  assign n11729 = ( x99 & ~n11634 ) | ( x99 & n11728 ) | ( ~n11634 & n11728 ) ;
  assign n11730 = ( x100 & ~n11631 ) | ( x100 & n11729 ) | ( ~n11631 & n11729 ) ;
  assign n11731 = ( x101 & ~n11628 ) | ( x101 & n11730 ) | ( ~n11628 & n11730 ) ;
  assign n11732 = ( x102 & ~n11625 ) | ( x102 & n11731 ) | ( ~n11625 & n11731 ) ;
  assign n11733 = ( x103 & ~n11622 ) | ( x103 & n11732 ) | ( ~n11622 & n11732 ) ;
  assign n11734 = ( x104 & ~n11580 ) | ( x104 & n11733 ) | ( ~n11580 & n11733 ) ;
  assign n11735 = ( x105 & ~n11506 ) | ( x105 & n11734 ) | ( ~n11506 & n11734 ) ;
  assign n11736 = ( x106 & ~n11515 ) | ( x106 & n11735 ) | ( ~n11515 & n11735 ) ;
  assign n11737 = ( x107 & ~n11503 ) | ( x107 & n11736 ) | ( ~n11503 & n11736 ) ;
  assign n11738 = ( x108 & ~n11577 ) | ( x108 & n11737 ) | ( ~n11577 & n11737 ) ;
  assign n11739 = ( x109 & ~n11574 ) | ( x109 & n11738 ) | ( ~n11574 & n11738 ) ;
  assign n11740 = ( x110 & ~n11571 ) | ( x110 & n11739 ) | ( ~n11571 & n11739 ) ;
  assign n11741 = ( x111 & ~n11568 ) | ( x111 & n11740 ) | ( ~n11568 & n11740 ) ;
  assign n11742 = ( x112 & ~n11565 ) | ( x112 & n11741 ) | ( ~n11565 & n11741 ) ;
  assign n11743 = ( x113 & ~n11562 ) | ( x113 & n11742 ) | ( ~n11562 & n11742 ) ;
  assign n11744 = ( x114 & ~n11559 ) | ( x114 & n11743 ) | ( ~n11559 & n11743 ) ;
  assign n11745 = ( x115 & ~n11556 ) | ( x115 & n11744 ) | ( ~n11556 & n11744 ) ;
  assign n11746 = ( x116 & ~n11553 ) | ( x116 & n11745 ) | ( ~n11553 & n11745 ) ;
  assign n11747 = ( x117 & ~n11550 ) | ( x117 & n11746 ) | ( ~n11550 & n11746 ) ;
  assign n11748 = ( x118 & ~n11547 ) | ( x118 & n11747 ) | ( ~n11547 & n11747 ) ;
  assign n11749 = ( x119 & ~n11544 ) | ( x119 & n11748 ) | ( ~n11544 & n11748 ) ;
  assign n11750 = ( x120 & ~n11541 ) | ( x120 & n11749 ) | ( ~n11541 & n11749 ) ;
  assign n11751 = ( x121 & ~n11538 ) | ( x121 & n11750 ) | ( ~n11538 & n11750 ) ;
  assign n11752 = ( x122 & ~n11501 ) | ( x122 & n11751 ) | ( ~n11501 & n11751 ) ;
  assign n11753 = ( x123 & ~n11535 ) | ( x123 & n11752 ) | ( ~n11535 & n11752 ) ;
  assign n11754 = ( ~x124 & n153 ) | ( ~x124 & n11681 ) | ( n153 & n11681 ) ;
  assign n11755 = ( n11724 & ~n11753 ) | ( n11724 & n11754 ) | ( ~n11753 & n11754 ) ;
  assign n11756 = n11753 | n11755 ;
  assign n11757 = ( ~n11681 & n11695 ) | ( ~n11681 & n11756 ) | ( n11695 & n11756 ) ;
  assign n11758 = n11757 ^ n11512 ^ 1'b0 ;
  assign n11759 = ( n11512 & n11705 ) | ( n11512 & ~n11758 ) | ( n11705 & ~n11758 ) ;
  assign n11760 = n11757 ^ n11619 ^ 1'b0 ;
  assign n11761 = ( n11619 & n11704 ) | ( n11619 & ~n11760 ) | ( n11704 & ~n11760 ) ;
  assign n11762 = n11757 ^ n11514 ^ 1'b0 ;
  assign n11763 = ( n11514 & n11703 ) | ( n11514 & ~n11762 ) | ( n11703 & ~n11762 ) ;
  assign n11764 = n11757 ^ n11517 ^ 1'b0 ;
  assign n11765 = ( n11517 & n11702 ) | ( n11517 & ~n11764 ) | ( n11702 & ~n11764 ) ;
  assign n11766 = n11757 ^ n11519 ^ 1'b0 ;
  assign n11767 = ( n11519 & n11701 ) | ( n11519 & ~n11766 ) | ( n11701 & ~n11766 ) ;
  assign n11768 = n11757 ^ n11521 ^ 1'b0 ;
  assign n11769 = ( n11521 & n11700 ) | ( n11521 & ~n11768 ) | ( n11700 & ~n11768 ) ;
  assign n11770 = n11757 ^ n11523 ^ 1'b0 ;
  assign n11771 = ( n11523 & n11699 ) | ( n11523 & ~n11770 ) | ( n11699 & ~n11770 ) ;
  assign n11772 = n11757 ^ n11525 ^ 1'b0 ;
  assign n11773 = ( n11525 & n11698 ) | ( n11525 & ~n11772 ) | ( n11698 & ~n11772 ) ;
  assign n11774 = n11757 ^ n11527 ^ 1'b0 ;
  assign n11775 = ( n11527 & n11697 ) | ( n11527 & ~n11774 ) | ( n11697 & ~n11774 ) ;
  assign n11776 = n11757 ^ n11529 ^ 1'b0 ;
  assign n11777 = ( n11529 & n11696 ) | ( n11529 & ~n11776 ) | ( n11696 & ~n11776 ) ;
  assign n11778 = n11695 & n11756 ;
  assign n11779 = n11751 ^ n11501 ^ x122 ;
  assign n11780 = n11757 ^ n11501 ^ 1'b0 ;
  assign n11781 = ( n11501 & n11779 ) | ( n11501 & ~n11780 ) | ( n11779 & ~n11780 ) ;
  assign n11782 = n11757 ^ n11646 ^ 1'b0 ;
  assign n11783 = ( n11646 & n11707 ) | ( n11646 & ~n11782 ) | ( n11707 & ~n11782 ) ;
  assign n11784 = n11757 ^ n11649 ^ 1'b0 ;
  assign n11785 = ( n11649 & n11725 ) | ( n11649 & ~n11784 ) | ( n11725 & ~n11784 ) ;
  assign n11786 = n11757 ^ n11652 ^ 1'b0 ;
  assign n11787 = ( n11652 & n11722 ) | ( n11652 & ~n11786 ) | ( n11722 & ~n11786 ) ;
  assign n11788 = n11757 ^ n11655 ^ 1'b0 ;
  assign n11789 = ( n11655 & n11721 ) | ( n11655 & ~n11788 ) | ( n11721 & ~n11788 ) ;
  assign n11790 = n11757 ^ n11508 ^ 1'b0 ;
  assign n11791 = ( n11508 & n11720 ) | ( n11508 & ~n11790 ) | ( n11720 & ~n11790 ) ;
  assign n11792 = n11757 ^ n11658 ^ 1'b0 ;
  assign n11793 = ( n11658 & n11719 ) | ( n11658 & ~n11792 ) | ( n11719 & ~n11792 ) ;
  assign n11794 = n11757 ^ n11583 ^ 1'b0 ;
  assign n11795 = ( n11583 & n11718 ) | ( n11583 & ~n11794 ) | ( n11718 & ~n11794 ) ;
  assign n11796 = n11757 ^ n11586 ^ 1'b0 ;
  assign n11797 = ( n11586 & n11717 ) | ( n11586 & ~n11796 ) | ( n11717 & ~n11796 ) ;
  assign n11798 = n11757 ^ n11510 ^ 1'b0 ;
  assign n11799 = ( n11510 & n11716 ) | ( n11510 & ~n11798 ) | ( n11716 & ~n11798 ) ;
  assign n11800 = n11757 ^ n11589 ^ 1'b0 ;
  assign n11801 = ( n11589 & n11715 ) | ( n11589 & ~n11800 ) | ( n11715 & ~n11800 ) ;
  assign n11802 = n11757 ^ n11592 ^ 1'b0 ;
  assign n11803 = ( n11592 & n11714 ) | ( n11592 & ~n11802 ) | ( n11714 & ~n11802 ) ;
  assign n11804 = n11757 ^ n11595 ^ 1'b0 ;
  assign n11805 = ( n11595 & n11713 ) | ( n11595 & ~n11804 ) | ( n11713 & ~n11804 ) ;
  assign n11806 = n11757 ^ n11598 ^ 1'b0 ;
  assign n11807 = ( n11598 & n11712 ) | ( n11598 & ~n11806 ) | ( n11712 & ~n11806 ) ;
  assign n11808 = n11757 ^ n11601 ^ 1'b0 ;
  assign n11809 = ( n11601 & n11711 ) | ( n11601 & ~n11808 ) | ( n11711 & ~n11808 ) ;
  assign n11810 = n11757 ^ n11604 ^ 1'b0 ;
  assign n11811 = ( n11604 & n11710 ) | ( n11604 & ~n11810 ) | ( n11710 & ~n11810 ) ;
  assign n11812 = n11757 ^ n11607 ^ 1'b0 ;
  assign n11813 = ( n11607 & n11709 ) | ( n11607 & ~n11812 ) | ( n11709 & ~n11812 ) ;
  assign n11814 = n11757 ^ n11610 ^ 1'b0 ;
  assign n11815 = ( n11610 & n11708 ) | ( n11610 & ~n11814 ) | ( n11708 & ~n11814 ) ;
  assign n11816 = n11757 ^ n11613 ^ 1'b0 ;
  assign n11817 = ( n11613 & n11688 ) | ( n11613 & ~n11816 ) | ( n11688 & ~n11816 ) ;
  assign n11818 = n11757 ^ n11616 ^ 1'b0 ;
  assign n11819 = ( n11616 & n11706 ) | ( n11616 & ~n11818 ) | ( n11706 & ~n11818 ) ;
  assign n11820 = n11757 ^ n11663 ^ 1'b0 ;
  assign n11821 = ( n11531 & n11663 ) | ( n11531 & n11820 ) | ( n11663 & n11820 ) ;
  assign n11822 = n11757 ^ n11661 ^ 1'b0 ;
  assign n11823 = ( n11660 & n11661 ) | ( n11660 & n11822 ) | ( n11661 & n11822 ) ;
  assign n11824 = n11752 ^ n11535 ^ x123 ;
  assign n11825 = n11757 ^ n11535 ^ 1'b0 ;
  assign n11826 = ( n11535 & n11824 ) | ( n11535 & ~n11825 ) | ( n11824 & ~n11825 ) ;
  assign n11827 = n11737 ^ n11577 ^ x108 ;
  assign n11828 = n11757 ^ n11577 ^ 1'b0 ;
  assign n11829 = ( n11577 & n11827 ) | ( n11577 & ~n11828 ) | ( n11827 & ~n11828 ) ;
  assign n11830 = n11736 ^ n11503 ^ x107 ;
  assign n11831 = n11757 ^ n11503 ^ 1'b0 ;
  assign n11832 = ( n11503 & n11830 ) | ( n11503 & ~n11831 ) | ( n11830 & ~n11831 ) ;
  assign n11833 = n11735 ^ n11515 ^ x106 ;
  assign n11834 = n11757 ^ n11515 ^ 1'b0 ;
  assign n11835 = ( n11515 & n11833 ) | ( n11515 & ~n11834 ) | ( n11833 & ~n11834 ) ;
  assign n11836 = n11734 ^ n11506 ^ x105 ;
  assign n11837 = n11757 ^ n11506 ^ 1'b0 ;
  assign n11838 = ( n11506 & n11836 ) | ( n11506 & ~n11837 ) | ( n11836 & ~n11837 ) ;
  assign n11839 = n11733 ^ n11580 ^ x104 ;
  assign n11840 = n11757 ^ n11580 ^ 1'b0 ;
  assign n11841 = ( n11580 & n11839 ) | ( n11580 & ~n11840 ) | ( n11839 & ~n11840 ) ;
  assign n11842 = n11732 ^ n11622 ^ x103 ;
  assign n11843 = n11757 ^ n11622 ^ 1'b0 ;
  assign n11844 = ( n11622 & n11842 ) | ( n11622 & ~n11843 ) | ( n11842 & ~n11843 ) ;
  assign n11845 = n11731 ^ n11625 ^ x102 ;
  assign n11846 = n11757 ^ n11625 ^ 1'b0 ;
  assign n11847 = ( n11625 & n11845 ) | ( n11625 & ~n11846 ) | ( n11845 & ~n11846 ) ;
  assign n11848 = n11730 ^ n11628 ^ x101 ;
  assign n11849 = n11757 ^ n11628 ^ 1'b0 ;
  assign n11850 = ( n11628 & n11848 ) | ( n11628 & ~n11849 ) | ( n11848 & ~n11849 ) ;
  assign n11851 = n11729 ^ n11631 ^ x100 ;
  assign n11852 = n11757 ^ n11631 ^ 1'b0 ;
  assign n11853 = ( n11631 & n11851 ) | ( n11631 & ~n11852 ) | ( n11851 & ~n11852 ) ;
  assign n11854 = n11728 ^ n11634 ^ x99 ;
  assign n11855 = n11757 ^ n11634 ^ 1'b0 ;
  assign n11856 = ( n11634 & n11854 ) | ( n11634 & ~n11855 ) | ( n11854 & ~n11855 ) ;
  assign n11857 = n11727 ^ n11637 ^ x98 ;
  assign n11858 = n11757 ^ n11637 ^ 1'b0 ;
  assign n11859 = ( n11637 & n11857 ) | ( n11637 & ~n11858 ) | ( n11857 & ~n11858 ) ;
  assign n11860 = n11726 ^ n11640 ^ x97 ;
  assign n11861 = n11757 ^ n11640 ^ 1'b0 ;
  assign n11862 = ( n11640 & n11860 ) | ( n11640 & ~n11861 ) | ( n11860 & ~n11861 ) ;
  assign n11863 = n11723 ^ n11643 ^ x96 ;
  assign n11864 = n11757 ^ n11643 ^ 1'b0 ;
  assign n11865 = ( n11643 & n11863 ) | ( n11643 & ~n11864 ) | ( n11863 & ~n11864 ) ;
  assign n11866 = n11750 ^ n11538 ^ x121 ;
  assign n11867 = n11757 ^ n11538 ^ 1'b0 ;
  assign n11868 = ( n11538 & n11866 ) | ( n11538 & ~n11867 ) | ( n11866 & ~n11867 ) ;
  assign n11869 = n11749 ^ n11541 ^ x120 ;
  assign n11870 = n11757 ^ n11541 ^ 1'b0 ;
  assign n11871 = ( n11541 & n11869 ) | ( n11541 & ~n11870 ) | ( n11869 & ~n11870 ) ;
  assign n11872 = n11748 ^ n11544 ^ x119 ;
  assign n11873 = n11757 ^ n11544 ^ 1'b0 ;
  assign n11874 = ( n11544 & n11872 ) | ( n11544 & ~n11873 ) | ( n11872 & ~n11873 ) ;
  assign n11875 = n11747 ^ n11547 ^ x118 ;
  assign n11876 = n11757 ^ n11547 ^ 1'b0 ;
  assign n11877 = ( n11547 & n11875 ) | ( n11547 & ~n11876 ) | ( n11875 & ~n11876 ) ;
  assign n11878 = n11746 ^ n11550 ^ x117 ;
  assign n11879 = n11757 ^ n11550 ^ 1'b0 ;
  assign n11880 = ( n11550 & n11878 ) | ( n11550 & ~n11879 ) | ( n11878 & ~n11879 ) ;
  assign n11881 = n11745 ^ n11553 ^ x116 ;
  assign n11882 = n11757 ^ n11553 ^ 1'b0 ;
  assign n11883 = ( n11553 & n11881 ) | ( n11553 & ~n11882 ) | ( n11881 & ~n11882 ) ;
  assign n11884 = n11744 ^ n11556 ^ x115 ;
  assign n11885 = n11757 ^ n11556 ^ 1'b0 ;
  assign n11886 = ( n11556 & n11884 ) | ( n11556 & ~n11885 ) | ( n11884 & ~n11885 ) ;
  assign n11887 = n11743 ^ n11559 ^ x114 ;
  assign n11888 = n11757 ^ n11559 ^ 1'b0 ;
  assign n11889 = ( n11559 & n11887 ) | ( n11559 & ~n11888 ) | ( n11887 & ~n11888 ) ;
  assign n11890 = n11742 ^ n11562 ^ x113 ;
  assign n11891 = n11757 ^ n11562 ^ 1'b0 ;
  assign n11892 = ( n11562 & n11890 ) | ( n11562 & ~n11891 ) | ( n11890 & ~n11891 ) ;
  assign n11893 = n11741 ^ n11565 ^ x112 ;
  assign n11894 = n11757 ^ n11565 ^ 1'b0 ;
  assign n11895 = ( n11565 & n11893 ) | ( n11565 & ~n11894 ) | ( n11893 & ~n11894 ) ;
  assign n11896 = n11740 ^ n11568 ^ x111 ;
  assign n11897 = n11757 ^ n11568 ^ 1'b0 ;
  assign n11898 = ( n11568 & n11896 ) | ( n11568 & ~n11897 ) | ( n11896 & ~n11897 ) ;
  assign n11899 = n11739 ^ n11571 ^ x110 ;
  assign n11900 = n11757 ^ n11571 ^ 1'b0 ;
  assign n11901 = ( n11571 & n11899 ) | ( n11571 & ~n11900 ) | ( n11899 & ~n11900 ) ;
  assign n11902 = n11738 ^ n11574 ^ x109 ;
  assign n11903 = n11757 ^ n11574 ^ 1'b0 ;
  assign n11904 = ( n11574 & n11902 ) | ( n11574 & ~n11903 ) | ( n11902 & ~n11903 ) ;
  assign n11905 = x64 & n11757 ;
  assign n11906 = n11905 ^ x64 ^ x3 ;
  assign n11907 = n11906 ^ n9064 ^ x65 ;
  assign n11908 = ( x65 & n9064 ) | ( x65 & n11907 ) | ( n9064 & n11907 ) ;
  assign n11909 = n11908 ^ n11823 ^ x66 ;
  assign n11910 = ( x66 & n11908 ) | ( x66 & n11909 ) | ( n11908 & n11909 ) ;
  assign n11911 = ( x67 & ~n11821 ) | ( x67 & n11910 ) | ( ~n11821 & n11910 ) ;
  assign n11912 = ( x68 & ~n11777 ) | ( x68 & n11911 ) | ( ~n11777 & n11911 ) ;
  assign n11913 = ( x69 & ~n11775 ) | ( x69 & n11912 ) | ( ~n11775 & n11912 ) ;
  assign n11914 = ( x70 & ~n11773 ) | ( x70 & n11913 ) | ( ~n11773 & n11913 ) ;
  assign n11915 = ( x71 & ~n11771 ) | ( x71 & n11914 ) | ( ~n11771 & n11914 ) ;
  assign n11916 = ( x72 & ~n11769 ) | ( x72 & n11915 ) | ( ~n11769 & n11915 ) ;
  assign n11917 = ( x73 & ~n11767 ) | ( x73 & n11916 ) | ( ~n11767 & n11916 ) ;
  assign n11918 = ( x74 & ~n11765 ) | ( x74 & n11917 ) | ( ~n11765 & n11917 ) ;
  assign n11919 = ( x75 & ~n11763 ) | ( x75 & n11918 ) | ( ~n11763 & n11918 ) ;
  assign n11920 = ( x76 & ~n11761 ) | ( x76 & n11919 ) | ( ~n11761 & n11919 ) ;
  assign n11921 = ( x77 & ~n11759 ) | ( x77 & n11920 ) | ( ~n11759 & n11920 ) ;
  assign n11922 = ( x78 & ~n11819 ) | ( x78 & n11921 ) | ( ~n11819 & n11921 ) ;
  assign n11923 = ( x79 & ~n11817 ) | ( x79 & n11922 ) | ( ~n11817 & n11922 ) ;
  assign n11924 = ( x80 & ~n11815 ) | ( x80 & n11923 ) | ( ~n11815 & n11923 ) ;
  assign n11925 = ( x81 & ~n11813 ) | ( x81 & n11924 ) | ( ~n11813 & n11924 ) ;
  assign n11926 = ( x82 & ~n11811 ) | ( x82 & n11925 ) | ( ~n11811 & n11925 ) ;
  assign n11927 = ( x83 & ~n11809 ) | ( x83 & n11926 ) | ( ~n11809 & n11926 ) ;
  assign n11928 = ( x84 & ~n11807 ) | ( x84 & n11927 ) | ( ~n11807 & n11927 ) ;
  assign n11929 = ( x85 & ~n11805 ) | ( x85 & n11928 ) | ( ~n11805 & n11928 ) ;
  assign n11930 = ( x86 & ~n11803 ) | ( x86 & n11929 ) | ( ~n11803 & n11929 ) ;
  assign n11931 = ( x87 & ~n11801 ) | ( x87 & n11930 ) | ( ~n11801 & n11930 ) ;
  assign n11932 = ( x88 & ~n11799 ) | ( x88 & n11931 ) | ( ~n11799 & n11931 ) ;
  assign n11933 = ( x89 & ~n11797 ) | ( x89 & n11932 ) | ( ~n11797 & n11932 ) ;
  assign n11934 = ( x90 & ~n11795 ) | ( x90 & n11933 ) | ( ~n11795 & n11933 ) ;
  assign n11935 = ( x91 & ~n11793 ) | ( x91 & n11934 ) | ( ~n11793 & n11934 ) ;
  assign n11936 = ( x92 & ~n11791 ) | ( x92 & n11935 ) | ( ~n11791 & n11935 ) ;
  assign n11937 = ( x93 & ~n11789 ) | ( x93 & n11936 ) | ( ~n11789 & n11936 ) ;
  assign n11938 = ( x94 & ~n11787 ) | ( x94 & n11937 ) | ( ~n11787 & n11937 ) ;
  assign n11939 = ( x95 & ~n11785 ) | ( x95 & n11938 ) | ( ~n11785 & n11938 ) ;
  assign n11940 = ( x96 & ~n11783 ) | ( x96 & n11939 ) | ( ~n11783 & n11939 ) ;
  assign n11941 = ( x97 & ~n11865 ) | ( x97 & n11940 ) | ( ~n11865 & n11940 ) ;
  assign n11942 = ( x98 & ~n11862 ) | ( x98 & n11941 ) | ( ~n11862 & n11941 ) ;
  assign n11943 = ( x99 & ~n11859 ) | ( x99 & n11942 ) | ( ~n11859 & n11942 ) ;
  assign n11944 = ( x100 & ~n11856 ) | ( x100 & n11943 ) | ( ~n11856 & n11943 ) ;
  assign n11945 = ( n147 & n153 ) | ( n147 & ~n11778 ) | ( n153 & ~n11778 ) ;
  assign n11946 = ( x101 & ~n11853 ) | ( x101 & n11944 ) | ( ~n11853 & n11944 ) ;
  assign n11947 = ( x102 & ~n11850 ) | ( x102 & n11946 ) | ( ~n11850 & n11946 ) ;
  assign n11948 = n11921 ^ n11819 ^ x78 ;
  assign n11949 = n11920 ^ n11759 ^ x77 ;
  assign n11950 = n11919 ^ n11761 ^ x76 ;
  assign n11951 = n11918 ^ n11763 ^ x75 ;
  assign n11952 = n11917 ^ n11765 ^ x74 ;
  assign n11953 = n11916 ^ n11767 ^ x73 ;
  assign n11954 = n11912 ^ n11775 ^ x69 ;
  assign n11955 = n11911 ^ n11777 ^ x68 ;
  assign n11956 = n322 | n11778 ;
  assign n11957 = x125 & n11956 ;
  assign n11958 = n153 & n11956 ;
  assign n11959 = ( n11945 & n11956 ) | ( n11945 & ~n11957 ) | ( n11956 & ~n11957 ) ;
  assign n11960 = ( x103 & ~n11847 ) | ( x103 & n11947 ) | ( ~n11847 & n11947 ) ;
  assign n11961 = ( x104 & ~n11844 ) | ( x104 & n11960 ) | ( ~n11844 & n11960 ) ;
  assign n11962 = ( x105 & ~n11841 ) | ( x105 & n11961 ) | ( ~n11841 & n11961 ) ;
  assign n11963 = ( x106 & ~n11838 ) | ( x106 & n11962 ) | ( ~n11838 & n11962 ) ;
  assign n11964 = ( x107 & ~n11835 ) | ( x107 & n11963 ) | ( ~n11835 & n11963 ) ;
  assign n11965 = ( x108 & ~n11832 ) | ( x108 & n11964 ) | ( ~n11832 & n11964 ) ;
  assign n11966 = ( x109 & ~n11829 ) | ( x109 & n11965 ) | ( ~n11829 & n11965 ) ;
  assign n11967 = ( x110 & ~n11904 ) | ( x110 & n11966 ) | ( ~n11904 & n11966 ) ;
  assign n11968 = ( x111 & ~n11901 ) | ( x111 & n11967 ) | ( ~n11901 & n11967 ) ;
  assign n11969 = ( x112 & ~n11898 ) | ( x112 & n11968 ) | ( ~n11898 & n11968 ) ;
  assign n11970 = ( x113 & ~n11895 ) | ( x113 & n11969 ) | ( ~n11895 & n11969 ) ;
  assign n11971 = ( x114 & ~n11892 ) | ( x114 & n11970 ) | ( ~n11892 & n11970 ) ;
  assign n11972 = ( x115 & ~n11889 ) | ( x115 & n11971 ) | ( ~n11889 & n11971 ) ;
  assign n11973 = ( x116 & ~n11886 ) | ( x116 & n11972 ) | ( ~n11886 & n11972 ) ;
  assign n11974 = ( x117 & ~n11883 ) | ( x117 & n11973 ) | ( ~n11883 & n11973 ) ;
  assign n11975 = ( x118 & ~n11880 ) | ( x118 & n11974 ) | ( ~n11880 & n11974 ) ;
  assign n11976 = ( x119 & ~n11877 ) | ( x119 & n11975 ) | ( ~n11877 & n11975 ) ;
  assign n11977 = ( x120 & ~n11874 ) | ( x120 & n11976 ) | ( ~n11874 & n11976 ) ;
  assign n11978 = ( x121 & ~n11871 ) | ( x121 & n11977 ) | ( ~n11871 & n11977 ) ;
  assign n11979 = ( x122 & ~n11868 ) | ( x122 & n11978 ) | ( ~n11868 & n11978 ) ;
  assign n11980 = ( x123 & ~n11781 ) | ( x123 & n11979 ) | ( ~n11781 & n11979 ) ;
  assign n11981 = n11980 ^ n11826 ^ x124 ;
  assign n11982 = ( x124 & ~n11826 ) | ( x124 & n11980 ) | ( ~n11826 & n11980 ) ;
  assign n11983 = n11959 | n11982 ;
  assign n11984 = ( ~n11956 & n11958 ) | ( ~n11956 & n11983 ) | ( n11958 & n11983 ) ;
  assign n11985 = n11984 ^ n11826 ^ 1'b0 ;
  assign n11986 = ( n11826 & n11981 ) | ( n11826 & ~n11985 ) | ( n11981 & ~n11985 ) ;
  assign n11987 = n11979 ^ n11781 ^ x123 ;
  assign n11988 = n11984 ^ n11781 ^ 1'b0 ;
  assign n11989 = ( n11781 & n11987 ) | ( n11781 & ~n11988 ) | ( n11987 & ~n11988 ) ;
  assign n11990 = n11977 ^ n11871 ^ x121 ;
  assign n11991 = n11984 ^ n11871 ^ 1'b0 ;
  assign n11992 = ( n11871 & n11990 ) | ( n11871 & ~n11991 ) | ( n11990 & ~n11991 ) ;
  assign n11993 = n11976 ^ n11874 ^ x120 ;
  assign n11994 = n11984 ^ n11874 ^ 1'b0 ;
  assign n11995 = ( n11874 & n11993 ) | ( n11874 & ~n11994 ) | ( n11993 & ~n11994 ) ;
  assign n11996 = n11975 ^ n11877 ^ x119 ;
  assign n11997 = n11984 ^ n11877 ^ 1'b0 ;
  assign n11998 = ( n11877 & n11996 ) | ( n11877 & ~n11997 ) | ( n11996 & ~n11997 ) ;
  assign n11999 = n11974 ^ n11880 ^ x118 ;
  assign n12000 = n11984 ^ n11880 ^ 1'b0 ;
  assign n12001 = ( n11880 & n11999 ) | ( n11880 & ~n12000 ) | ( n11999 & ~n12000 ) ;
  assign n12002 = n11973 ^ n11883 ^ x117 ;
  assign n12003 = n11984 ^ n11883 ^ 1'b0 ;
  assign n12004 = ( n11883 & n12002 ) | ( n11883 & ~n12003 ) | ( n12002 & ~n12003 ) ;
  assign n12005 = n11984 ^ n11886 ^ 1'b0 ;
  assign n12006 = n11984 ^ n11819 ^ 1'b0 ;
  assign n12007 = ( n11819 & n11948 ) | ( n11819 & ~n12006 ) | ( n11948 & ~n12006 ) ;
  assign n12008 = n11984 ^ n11759 ^ 1'b0 ;
  assign n12009 = n11972 ^ n11886 ^ x116 ;
  assign n12010 = ( n11886 & ~n12005 ) | ( n11886 & n12009 ) | ( ~n12005 & n12009 ) ;
  assign n12011 = ( n11759 & n11949 ) | ( n11759 & ~n12008 ) | ( n11949 & ~n12008 ) ;
  assign n12012 = n11984 ^ n11761 ^ 1'b0 ;
  assign n12013 = ( n11761 & n11950 ) | ( n11761 & ~n12012 ) | ( n11950 & ~n12012 ) ;
  assign n12014 = n11984 ^ n11763 ^ 1'b0 ;
  assign n12015 = ( n11763 & n11951 ) | ( n11763 & ~n12014 ) | ( n11951 & ~n12014 ) ;
  assign n12016 = n11984 ^ n11765 ^ 1'b0 ;
  assign n12017 = ( n11765 & n11952 ) | ( n11765 & ~n12016 ) | ( n11952 & ~n12016 ) ;
  assign n12018 = n11984 ^ n11767 ^ 1'b0 ;
  assign n12019 = ( n11767 & n11953 ) | ( n11767 & ~n12018 ) | ( n11953 & ~n12018 ) ;
  assign n12020 = n11984 ^ n11775 ^ 1'b0 ;
  assign n12021 = ( n11775 & n11954 ) | ( n11775 & ~n12020 ) | ( n11954 & ~n12020 ) ;
  assign n12022 = n11984 ^ n11777 ^ 1'b0 ;
  assign n12023 = ( n11777 & n11955 ) | ( n11777 & ~n12022 ) | ( n11955 & ~n12022 ) ;
  assign n12024 = n11984 ^ n11909 ^ 1'b0 ;
  assign n12025 = ( n11823 & n11909 ) | ( n11823 & n12024 ) | ( n11909 & n12024 ) ;
  assign n12026 = n11984 ^ n11907 ^ 1'b0 ;
  assign n12027 = ( n11906 & n11907 ) | ( n11906 & n12026 ) | ( n11907 & n12026 ) ;
  assign n12028 = n11958 & n11983 ;
  assign n12029 = n11971 ^ n11889 ^ x115 ;
  assign n12030 = n11984 ^ n11889 ^ 1'b0 ;
  assign n12031 = ( n11889 & n12029 ) | ( n11889 & ~n12030 ) | ( n12029 & ~n12030 ) ;
  assign n12032 = n11970 ^ n11892 ^ x114 ;
  assign n12033 = n11984 ^ n11892 ^ 1'b0 ;
  assign n12034 = ( n11892 & n12032 ) | ( n11892 & ~n12033 ) | ( n12032 & ~n12033 ) ;
  assign n12035 = n11969 ^ n11895 ^ x113 ;
  assign n12036 = n11984 ^ n11895 ^ 1'b0 ;
  assign n12037 = ( n11895 & n12035 ) | ( n11895 & ~n12036 ) | ( n12035 & ~n12036 ) ;
  assign n12038 = n11937 ^ n11787 ^ x94 ;
  assign n12039 = n11984 ^ n11787 ^ 1'b0 ;
  assign n12040 = ( n11787 & n12038 ) | ( n11787 & ~n12039 ) | ( n12038 & ~n12039 ) ;
  assign n12041 = n11936 ^ n11789 ^ x93 ;
  assign n12042 = n11984 ^ n11789 ^ 1'b0 ;
  assign n12043 = ( n11789 & n12041 ) | ( n11789 & ~n12042 ) | ( n12041 & ~n12042 ) ;
  assign n12044 = n11935 ^ n11791 ^ x92 ;
  assign n12045 = n11984 ^ n11791 ^ 1'b0 ;
  assign n12046 = ( n11791 & n12044 ) | ( n11791 & ~n12045 ) | ( n12044 & ~n12045 ) ;
  assign n12047 = n11934 ^ n11793 ^ x91 ;
  assign n12048 = n11984 ^ n11793 ^ 1'b0 ;
  assign n12049 = ( n11793 & n12047 ) | ( n11793 & ~n12048 ) | ( n12047 & ~n12048 ) ;
  assign n12050 = n11933 ^ n11795 ^ x90 ;
  assign n12051 = n11984 ^ n11795 ^ 1'b0 ;
  assign n12052 = ( n11795 & n12050 ) | ( n11795 & ~n12051 ) | ( n12050 & ~n12051 ) ;
  assign n12053 = n11932 ^ n11797 ^ x89 ;
  assign n12054 = n11984 ^ n11797 ^ 1'b0 ;
  assign n12055 = ( n11797 & n12053 ) | ( n11797 & ~n12054 ) | ( n12053 & ~n12054 ) ;
  assign n12056 = n11931 ^ n11799 ^ x88 ;
  assign n12057 = n11984 ^ n11799 ^ 1'b0 ;
  assign n12058 = ( n11799 & n12056 ) | ( n11799 & ~n12057 ) | ( n12056 & ~n12057 ) ;
  assign n12059 = n11928 ^ n11805 ^ x85 ;
  assign n12060 = n11984 ^ n11805 ^ 1'b0 ;
  assign n12061 = ( n11805 & n12059 ) | ( n11805 & ~n12060 ) | ( n12059 & ~n12060 ) ;
  assign n12062 = n11927 ^ n11807 ^ x84 ;
  assign n12063 = n11984 ^ n11807 ^ 1'b0 ;
  assign n12064 = ( n11807 & n12062 ) | ( n11807 & ~n12063 ) | ( n12062 & ~n12063 ) ;
  assign n12065 = n11926 ^ n11809 ^ x83 ;
  assign n12066 = n11984 ^ n11809 ^ 1'b0 ;
  assign n12067 = ( n11809 & n12065 ) | ( n11809 & ~n12066 ) | ( n12065 & ~n12066 ) ;
  assign n12068 = n11925 ^ n11811 ^ x82 ;
  assign n12069 = n11984 ^ n11811 ^ 1'b0 ;
  assign n12070 = ( n11811 & n12068 ) | ( n11811 & ~n12069 ) | ( n12068 & ~n12069 ) ;
  assign n12071 = n11924 ^ n11813 ^ x81 ;
  assign n12072 = n11984 ^ n11813 ^ 1'b0 ;
  assign n12073 = ( n11813 & n12071 ) | ( n11813 & ~n12072 ) | ( n12071 & ~n12072 ) ;
  assign n12074 = n11923 ^ n11815 ^ x80 ;
  assign n12075 = n11984 ^ n11815 ^ 1'b0 ;
  assign n12076 = ( n11815 & n12074 ) | ( n11815 & ~n12075 ) | ( n12074 & ~n12075 ) ;
  assign n12077 = n11922 ^ n11817 ^ x79 ;
  assign n12078 = n11984 ^ n11817 ^ 1'b0 ;
  assign n12079 = ( n11817 & n12077 ) | ( n11817 & ~n12078 ) | ( n12077 & ~n12078 ) ;
  assign n12080 = n11914 ^ n11771 ^ x71 ;
  assign n12081 = n11984 ^ n11771 ^ 1'b0 ;
  assign n12082 = ( n11771 & n12080 ) | ( n11771 & ~n12081 ) | ( n12080 & ~n12081 ) ;
  assign n12083 = n11913 ^ n11773 ^ x70 ;
  assign n12084 = n11984 ^ n11773 ^ 1'b0 ;
  assign n12085 = ( n11773 & n12083 ) | ( n11773 & ~n12084 ) | ( n12083 & ~n12084 ) ;
  assign n12086 = n11968 ^ n11898 ^ x112 ;
  assign n12087 = n11984 ^ n11898 ^ 1'b0 ;
  assign n12088 = ( n11898 & n12086 ) | ( n11898 & ~n12087 ) | ( n12086 & ~n12087 ) ;
  assign n12089 = n11967 ^ n11901 ^ x111 ;
  assign n12090 = n11984 ^ n11901 ^ 1'b0 ;
  assign n12091 = ( n11901 & n12089 ) | ( n11901 & ~n12090 ) | ( n12089 & ~n12090 ) ;
  assign n12092 = n11966 ^ n11904 ^ x110 ;
  assign n12093 = n11984 ^ n11904 ^ 1'b0 ;
  assign n12094 = ( n11904 & n12092 ) | ( n11904 & ~n12093 ) | ( n12092 & ~n12093 ) ;
  assign n12095 = n11965 ^ n11829 ^ x109 ;
  assign n12096 = n11984 ^ n11829 ^ 1'b0 ;
  assign n12097 = ( n11829 & n12095 ) | ( n11829 & ~n12096 ) | ( n12095 & ~n12096 ) ;
  assign n12098 = n11964 ^ n11832 ^ x108 ;
  assign n12099 = n11984 ^ n11832 ^ 1'b0 ;
  assign n12100 = ( n11832 & n12098 ) | ( n11832 & ~n12099 ) | ( n12098 & ~n12099 ) ;
  assign n12101 = n11963 ^ n11835 ^ x107 ;
  assign n12102 = n11984 ^ n11835 ^ 1'b0 ;
  assign n12103 = ( n11835 & n12101 ) | ( n11835 & ~n12102 ) | ( n12101 & ~n12102 ) ;
  assign n12104 = n11984 ^ n11838 ^ 1'b0 ;
  assign n12105 = n11961 ^ n11841 ^ x105 ;
  assign n12106 = n11984 ^ n11841 ^ 1'b0 ;
  assign n12107 = ( n11841 & n12105 ) | ( n11841 & ~n12106 ) | ( n12105 & ~n12106 ) ;
  assign n12108 = n11960 ^ n11844 ^ x104 ;
  assign n12109 = n11984 ^ n11844 ^ 1'b0 ;
  assign n12110 = n11962 ^ n11838 ^ x106 ;
  assign n12111 = ( n11838 & ~n12104 ) | ( n11838 & n12110 ) | ( ~n12104 & n12110 ) ;
  assign n12112 = ( n11844 & n12108 ) | ( n11844 & ~n12109 ) | ( n12108 & ~n12109 ) ;
  assign n12113 = n11947 ^ n11847 ^ x103 ;
  assign n12114 = n11984 ^ n11847 ^ 1'b0 ;
  assign n12115 = ( n11847 & n12113 ) | ( n11847 & ~n12114 ) | ( n12113 & ~n12114 ) ;
  assign n12116 = n11946 ^ n11850 ^ x102 ;
  assign n12117 = n11984 ^ n11850 ^ 1'b0 ;
  assign n12118 = ( n11850 & n12116 ) | ( n11850 & ~n12117 ) | ( n12116 & ~n12117 ) ;
  assign n12119 = n11943 ^ n11856 ^ x100 ;
  assign n12120 = n11984 ^ n11856 ^ 1'b0 ;
  assign n12121 = ( n11856 & n12119 ) | ( n11856 & ~n12120 ) | ( n12119 & ~n12120 ) ;
  assign n12122 = n11942 ^ n11859 ^ x99 ;
  assign n12123 = n11984 ^ n11859 ^ 1'b0 ;
  assign n12124 = ( n11859 & n12122 ) | ( n11859 & ~n12123 ) | ( n12122 & ~n12123 ) ;
  assign n12125 = n11940 ^ n11865 ^ x97 ;
  assign n12126 = n11984 ^ n11865 ^ 1'b0 ;
  assign n12127 = ( n11865 & n12125 ) | ( n11865 & ~n12126 ) | ( n12125 & ~n12126 ) ;
  assign n12128 = n11939 ^ n11783 ^ x96 ;
  assign n12129 = n11984 ^ n11783 ^ 1'b0 ;
  assign n12130 = ( n11783 & n12128 ) | ( n11783 & ~n12129 ) | ( n12128 & ~n12129 ) ;
  assign n12131 = n11938 ^ n11785 ^ x95 ;
  assign n12132 = n11984 ^ n11785 ^ 1'b0 ;
  assign n12133 = ( n11785 & n12131 ) | ( n11785 & ~n12132 ) | ( n12131 & ~n12132 ) ;
  assign n12134 = n11978 ^ n11868 ^ x122 ;
  assign n12135 = n11984 ^ n11868 ^ 1'b0 ;
  assign n12136 = ( n11868 & n12134 ) | ( n11868 & ~n12135 ) | ( n12134 & ~n12135 ) ;
  assign n12137 = n11944 ^ n11853 ^ x101 ;
  assign n12138 = n11984 ^ n11853 ^ 1'b0 ;
  assign n12139 = ( n11853 & n12137 ) | ( n11853 & ~n12138 ) | ( n12137 & ~n12138 ) ;
  assign n12140 = n11941 ^ n11862 ^ x98 ;
  assign n12141 = n11984 ^ n11862 ^ 1'b0 ;
  assign n12142 = ( n11862 & n12140 ) | ( n11862 & ~n12141 ) | ( n12140 & ~n12141 ) ;
  assign n12143 = n11930 ^ n11801 ^ x87 ;
  assign n12144 = n11984 ^ n11801 ^ 1'b0 ;
  assign n12145 = n11929 ^ n11803 ^ x86 ;
  assign n12146 = n11984 ^ n11803 ^ 1'b0 ;
  assign n12147 = ( n11803 & n12145 ) | ( n11803 & ~n12146 ) | ( n12145 & ~n12146 ) ;
  assign n12148 = n11915 ^ n11769 ^ x72 ;
  assign n12149 = n11984 ^ n11769 ^ 1'b0 ;
  assign n12150 = ( n11769 & n12148 ) | ( n11769 & ~n12149 ) | ( n12148 & ~n12149 ) ;
  assign n12151 = n11910 ^ n11821 ^ x67 ;
  assign n12152 = n11984 ^ n11821 ^ 1'b0 ;
  assign n12153 = ( n11821 & n12151 ) | ( n11821 & ~n12152 ) | ( n12151 & ~n12152 ) ;
  assign n12154 = ( n11801 & n12143 ) | ( n11801 & ~n12144 ) | ( n12143 & ~n12144 ) ;
  assign n12155 = x64 & n11984 ;
  assign n12156 = n12155 ^ x64 ^ x2 ;
  assign n12157 = n12156 ^ n9313 ^ x65 ;
  assign n12158 = ( x65 & n9313 ) | ( x65 & n12157 ) | ( n9313 & n12157 ) ;
  assign n12159 = n12158 ^ n12027 ^ x66 ;
  assign n12160 = ( x66 & n12158 ) | ( x66 & n12159 ) | ( n12158 & n12159 ) ;
  assign n12161 = ( x67 & ~n12025 ) | ( x67 & n12160 ) | ( ~n12025 & n12160 ) ;
  assign n12162 = ( x68 & ~n12153 ) | ( x68 & n12161 ) | ( ~n12153 & n12161 ) ;
  assign n12163 = ( x69 & ~n12023 ) | ( x69 & n12162 ) | ( ~n12023 & n12162 ) ;
  assign n12164 = ( x70 & ~n12021 ) | ( x70 & n12163 ) | ( ~n12021 & n12163 ) ;
  assign n12165 = n322 | n12028 ;
  assign n12166 = n147 & n12165 ;
  assign n12167 = ( x127 & n147 ) | ( x127 & ~n12028 ) | ( n147 & ~n12028 ) ;
  assign n12168 = x126 & n12165 ;
  assign n12169 = ( n12165 & n12167 ) | ( n12165 & ~n12168 ) | ( n12167 & ~n12168 ) ;
  assign n12170 = n12162 ^ n12023 ^ x69 ;
  assign n12171 = n12161 ^ n12153 ^ x68 ;
  assign n12172 = n12160 ^ n12025 ^ x67 ;
  assign n12173 = ( x71 & ~n12085 ) | ( x71 & n12164 ) | ( ~n12085 & n12164 ) ;
  assign n12174 = ( x72 & ~n12082 ) | ( x72 & n12173 ) | ( ~n12082 & n12173 ) ;
  assign n12175 = ( x73 & ~n12150 ) | ( x73 & n12174 ) | ( ~n12150 & n12174 ) ;
  assign n12176 = ( x74 & ~n12019 ) | ( x74 & n12175 ) | ( ~n12019 & n12175 ) ;
  assign n12177 = ( x75 & ~n12017 ) | ( x75 & n12176 ) | ( ~n12017 & n12176 ) ;
  assign n12178 = ( x76 & ~n12015 ) | ( x76 & n12177 ) | ( ~n12015 & n12177 ) ;
  assign n12179 = ( x77 & ~n12013 ) | ( x77 & n12178 ) | ( ~n12013 & n12178 ) ;
  assign n12180 = ( x78 & ~n12011 ) | ( x78 & n12179 ) | ( ~n12011 & n12179 ) ;
  assign n12181 = ( x79 & ~n12007 ) | ( x79 & n12180 ) | ( ~n12007 & n12180 ) ;
  assign n12182 = ( x80 & ~n12079 ) | ( x80 & n12181 ) | ( ~n12079 & n12181 ) ;
  assign n12183 = ( x81 & ~n12076 ) | ( x81 & n12182 ) | ( ~n12076 & n12182 ) ;
  assign n12184 = ( x82 & ~n12073 ) | ( x82 & n12183 ) | ( ~n12073 & n12183 ) ;
  assign n12185 = ( x83 & ~n12070 ) | ( x83 & n12184 ) | ( ~n12070 & n12184 ) ;
  assign n12186 = ( x84 & ~n12067 ) | ( x84 & n12185 ) | ( ~n12067 & n12185 ) ;
  assign n12187 = ( x85 & ~n12064 ) | ( x85 & n12186 ) | ( ~n12064 & n12186 ) ;
  assign n12188 = ( x86 & ~n12061 ) | ( x86 & n12187 ) | ( ~n12061 & n12187 ) ;
  assign n12189 = ( x87 & ~n12147 ) | ( x87 & n12188 ) | ( ~n12147 & n12188 ) ;
  assign n12190 = ( x88 & ~n12154 ) | ( x88 & n12189 ) | ( ~n12154 & n12189 ) ;
  assign n12191 = ( x89 & ~n12058 ) | ( x89 & n12190 ) | ( ~n12058 & n12190 ) ;
  assign n12192 = ( x90 & ~n12055 ) | ( x90 & n12191 ) | ( ~n12055 & n12191 ) ;
  assign n12193 = ( x91 & ~n12052 ) | ( x91 & n12192 ) | ( ~n12052 & n12192 ) ;
  assign n12194 = ( x92 & ~n12049 ) | ( x92 & n12193 ) | ( ~n12049 & n12193 ) ;
  assign n12195 = ( x93 & ~n12046 ) | ( x93 & n12194 ) | ( ~n12046 & n12194 ) ;
  assign n12196 = ( x94 & ~n12043 ) | ( x94 & n12195 ) | ( ~n12043 & n12195 ) ;
  assign n12197 = ( x95 & ~n12040 ) | ( x95 & n12196 ) | ( ~n12040 & n12196 ) ;
  assign n12198 = ( x96 & ~n12133 ) | ( x96 & n12197 ) | ( ~n12133 & n12197 ) ;
  assign n12199 = ( x97 & ~n12130 ) | ( x97 & n12198 ) | ( ~n12130 & n12198 ) ;
  assign n12200 = ( x98 & ~n12127 ) | ( x98 & n12199 ) | ( ~n12127 & n12199 ) ;
  assign n12201 = ( x99 & ~n12142 ) | ( x99 & n12200 ) | ( ~n12142 & n12200 ) ;
  assign n12202 = ( x100 & ~n12124 ) | ( x100 & n12201 ) | ( ~n12124 & n12201 ) ;
  assign n12203 = ( x101 & ~n12121 ) | ( x101 & n12202 ) | ( ~n12121 & n12202 ) ;
  assign n12204 = ( x102 & ~n12139 ) | ( x102 & n12203 ) | ( ~n12139 & n12203 ) ;
  assign n12205 = n12174 ^ n12150 ^ x73 ;
  assign n12206 = n12173 ^ n12082 ^ x72 ;
  assign n12207 = ( x103 & ~n12118 ) | ( x103 & n12204 ) | ( ~n12118 & n12204 ) ;
  assign n12208 = ( x104 & ~n12115 ) | ( x104 & n12207 ) | ( ~n12115 & n12207 ) ;
  assign n12209 = ( x105 & ~n12112 ) | ( x105 & n12208 ) | ( ~n12112 & n12208 ) ;
  assign n12210 = ( x106 & ~n12107 ) | ( x106 & n12209 ) | ( ~n12107 & n12209 ) ;
  assign n12211 = n12164 ^ n12085 ^ x71 ;
  assign n12212 = n12208 ^ n12112 ^ x105 ;
  assign n12213 = n12163 ^ n12021 ^ x70 ;
  assign n12214 = n12207 ^ n12115 ^ x104 ;
  assign n12215 = n12209 ^ n12107 ^ x106 ;
  assign n12216 = ( x107 & ~n12111 ) | ( x107 & n12210 ) | ( ~n12111 & n12210 ) ;
  assign n12217 = n12216 ^ n12103 ^ x108 ;
  assign n12218 = n12210 ^ n12111 ^ x107 ;
  assign n12219 = n12204 ^ n12118 ^ x103 ;
  assign n12220 = ( x108 & ~n12103 ) | ( x108 & n12216 ) | ( ~n12103 & n12216 ) ;
  assign n12221 = ( x109 & ~n12100 ) | ( x109 & n12220 ) | ( ~n12100 & n12220 ) ;
  assign n12222 = ( x110 & ~n12097 ) | ( x110 & n12221 ) | ( ~n12097 & n12221 ) ;
  assign n12223 = ( x111 & ~n12094 ) | ( x111 & n12222 ) | ( ~n12094 & n12222 ) ;
  assign n12224 = ( x112 & ~n12091 ) | ( x112 & n12223 ) | ( ~n12091 & n12223 ) ;
  assign n12225 = ( x113 & ~n12088 ) | ( x113 & n12224 ) | ( ~n12088 & n12224 ) ;
  assign n12226 = ( x114 & ~n12037 ) | ( x114 & n12225 ) | ( ~n12037 & n12225 ) ;
  assign n12227 = ( x115 & ~n12034 ) | ( x115 & n12226 ) | ( ~n12034 & n12226 ) ;
  assign n12228 = ( x116 & ~n12031 ) | ( x116 & n12227 ) | ( ~n12031 & n12227 ) ;
  assign n12229 = ( x117 & ~n12010 ) | ( x117 & n12228 ) | ( ~n12010 & n12228 ) ;
  assign n12230 = ( x118 & ~n12004 ) | ( x118 & n12229 ) | ( ~n12004 & n12229 ) ;
  assign n12231 = ( x119 & ~n12001 ) | ( x119 & n12230 ) | ( ~n12001 & n12230 ) ;
  assign n12232 = ( x120 & ~n11998 ) | ( x120 & n12231 ) | ( ~n11998 & n12231 ) ;
  assign n12233 = ( x121 & ~n11995 ) | ( x121 & n12232 ) | ( ~n11995 & n12232 ) ;
  assign n12234 = ( x122 & ~n11992 ) | ( x122 & n12233 ) | ( ~n11992 & n12233 ) ;
  assign n12235 = ( x123 & ~n12136 ) | ( x123 & n12234 ) | ( ~n12136 & n12234 ) ;
  assign n12236 = ( x124 & ~n11989 ) | ( x124 & n12235 ) | ( ~n11989 & n12235 ) ;
  assign n12237 = ( x125 & ~n11986 ) | ( x125 & n12236 ) | ( ~n11986 & n12236 ) ;
  assign n12238 = n12169 | n12237 ;
  assign n12239 = ( ~n12165 & n12166 ) | ( ~n12165 & n12238 ) | ( n12166 & n12238 ) ;
  assign n12240 = n12239 ^ n12118 ^ 1'b0 ;
  assign n12241 = ( n12118 & n12219 ) | ( n12118 & ~n12240 ) | ( n12219 & ~n12240 ) ;
  assign n12242 = n12239 ^ n12150 ^ 1'b0 ;
  assign n12243 = n12239 ^ n12111 ^ 1'b0 ;
  assign n12244 = n12235 ^ n11989 ^ x124 ;
  assign n12245 = ( n12111 & n12218 ) | ( n12111 & ~n12243 ) | ( n12218 & ~n12243 ) ;
  assign n12246 = n12239 ^ n12115 ^ 1'b0 ;
  assign n12247 = n12239 ^ n12082 ^ 1'b0 ;
  assign n12248 = ( n12150 & n12205 ) | ( n12150 & ~n12242 ) | ( n12205 & ~n12242 ) ;
  assign n12249 = n12239 ^ n12107 ^ 1'b0 ;
  assign n12250 = n12239 ^ n12021 ^ 1'b0 ;
  assign n12251 = ( n12107 & n12215 ) | ( n12107 & ~n12249 ) | ( n12215 & ~n12249 ) ;
  assign n12252 = n12239 ^ n12025 ^ 1'b0 ;
  assign n12253 = ( n12025 & n12172 ) | ( n12025 & ~n12252 ) | ( n12172 & ~n12252 ) ;
  assign n12254 = n12239 ^ n12159 ^ 1'b0 ;
  assign n12255 = n12239 ^ n12112 ^ 1'b0 ;
  assign n12256 = n12239 ^ n12157 ^ 1'b0 ;
  assign n12257 = ~n12166 & n12238 ;
  assign n12258 = ( n12027 & n12159 ) | ( n12027 & n12254 ) | ( n12159 & n12254 ) ;
  assign n12259 = ( n12082 & n12206 ) | ( n12082 & ~n12247 ) | ( n12206 & ~n12247 ) ;
  assign n12260 = ( n12112 & n12212 ) | ( n12112 & ~n12255 ) | ( n12212 & ~n12255 ) ;
  assign n12261 = n12239 ^ n12153 ^ 1'b0 ;
  assign n12262 = ( n12153 & n12171 ) | ( n12153 & ~n12261 ) | ( n12171 & ~n12261 ) ;
  assign n12263 = n12239 ^ n12023 ^ 1'b0 ;
  assign n12264 = n12239 ^ n12085 ^ 1'b0 ;
  assign n12265 = ( n12156 & n12157 ) | ( n12156 & n12256 ) | ( n12157 & n12256 ) ;
  assign n12266 = ( n322 & n12238 ) | ( n322 & ~n12257 ) | ( n12238 & ~n12257 ) ;
  assign n12267 = ( n12085 & n12211 ) | ( n12085 & ~n12264 ) | ( n12211 & ~n12264 ) ;
  assign n12268 = ( n12115 & n12214 ) | ( n12115 & ~n12246 ) | ( n12214 & ~n12246 ) ;
  assign n12269 = n12239 ^ n11989 ^ 1'b0 ;
  assign n12270 = ( n12021 & n12213 ) | ( n12021 & ~n12250 ) | ( n12213 & ~n12250 ) ;
  assign n12271 = ( n12023 & n12170 ) | ( n12023 & ~n12263 ) | ( n12170 & ~n12263 ) ;
  assign n12272 = ( n11989 & n12244 ) | ( n11989 & ~n12269 ) | ( n12244 & ~n12269 ) ;
  assign n12273 = n12239 ^ n12103 ^ 1'b0 ;
  assign n12274 = ( n12103 & n12217 ) | ( n12103 & ~n12273 ) | ( n12217 & ~n12273 ) ;
  assign n12275 = n12236 ^ n11986 ^ x125 ;
  assign n12276 = n12239 ^ n11986 ^ 1'b0 ;
  assign n12277 = ( n11986 & n12275 ) | ( n11986 & ~n12276 ) | ( n12275 & ~n12276 ) ;
  assign n12278 = n12234 ^ n12136 ^ x123 ;
  assign n12279 = n12239 ^ n12136 ^ 1'b0 ;
  assign n12280 = ( n12136 & n12278 ) | ( n12136 & ~n12279 ) | ( n12278 & ~n12279 ) ;
  assign n12281 = n12233 ^ n11992 ^ x122 ;
  assign n12282 = n12239 ^ n11992 ^ 1'b0 ;
  assign n12283 = ( n11992 & n12281 ) | ( n11992 & ~n12282 ) | ( n12281 & ~n12282 ) ;
  assign n12284 = n12232 ^ n11995 ^ x121 ;
  assign n12285 = n12239 ^ n11995 ^ 1'b0 ;
  assign n12286 = ( n11995 & n12284 ) | ( n11995 & ~n12285 ) | ( n12284 & ~n12285 ) ;
  assign n12287 = n12231 ^ n11998 ^ x120 ;
  assign n12288 = n12239 ^ n11998 ^ 1'b0 ;
  assign n12289 = ( n11998 & n12287 ) | ( n11998 & ~n12288 ) | ( n12287 & ~n12288 ) ;
  assign n12290 = n12230 ^ n12001 ^ x119 ;
  assign n12291 = n12239 ^ n12001 ^ 1'b0 ;
  assign n12292 = ( n12001 & n12290 ) | ( n12001 & ~n12291 ) | ( n12290 & ~n12291 ) ;
  assign n12293 = n12229 ^ n12004 ^ x118 ;
  assign n12294 = n12239 ^ n12004 ^ 1'b0 ;
  assign n12295 = ( n12004 & n12293 ) | ( n12004 & ~n12294 ) | ( n12293 & ~n12294 ) ;
  assign n12296 = n12228 ^ n12010 ^ x117 ;
  assign n12297 = n12239 ^ n12010 ^ 1'b0 ;
  assign n12298 = ( n12010 & n12296 ) | ( n12010 & ~n12297 ) | ( n12296 & ~n12297 ) ;
  assign n12299 = n12227 ^ n12031 ^ x116 ;
  assign n12300 = n12239 ^ n12031 ^ 1'b0 ;
  assign n12301 = ( n12031 & n12299 ) | ( n12031 & ~n12300 ) | ( n12299 & ~n12300 ) ;
  assign n12302 = n12226 ^ n12034 ^ x115 ;
  assign n12303 = n12239 ^ n12034 ^ 1'b0 ;
  assign n12304 = ( n12034 & n12302 ) | ( n12034 & ~n12303 ) | ( n12302 & ~n12303 ) ;
  assign n12305 = n12225 ^ n12037 ^ x114 ;
  assign n12306 = n12239 ^ n12037 ^ 1'b0 ;
  assign n12307 = ( n12037 & n12305 ) | ( n12037 & ~n12306 ) | ( n12305 & ~n12306 ) ;
  assign n12308 = n12224 ^ n12088 ^ x113 ;
  assign n12309 = n12239 ^ n12088 ^ 1'b0 ;
  assign n12310 = ( n12088 & n12308 ) | ( n12088 & ~n12309 ) | ( n12308 & ~n12309 ) ;
  assign n12311 = n12223 ^ n12091 ^ x112 ;
  assign n12312 = n12239 ^ n12091 ^ 1'b0 ;
  assign n12313 = ( n12091 & n12311 ) | ( n12091 & ~n12312 ) | ( n12311 & ~n12312 ) ;
  assign n12314 = n12222 ^ n12094 ^ x111 ;
  assign n12315 = n12239 ^ n12094 ^ 1'b0 ;
  assign n12316 = ( n12094 & n12314 ) | ( n12094 & ~n12315 ) | ( n12314 & ~n12315 ) ;
  assign n12317 = n12221 ^ n12097 ^ x110 ;
  assign n12318 = n12239 ^ n12097 ^ 1'b0 ;
  assign n12319 = ( n12097 & n12317 ) | ( n12097 & ~n12318 ) | ( n12317 & ~n12318 ) ;
  assign n12320 = n12220 ^ n12100 ^ x109 ;
  assign n12321 = n12239 ^ n12100 ^ 1'b0 ;
  assign n12322 = ( n12100 & n12320 ) | ( n12100 & ~n12321 ) | ( n12320 & ~n12321 ) ;
  assign n12323 = n12203 ^ n12139 ^ x102 ;
  assign n12324 = n12239 ^ n12139 ^ 1'b0 ;
  assign n12325 = ( n12139 & n12323 ) | ( n12139 & ~n12324 ) | ( n12323 & ~n12324 ) ;
  assign n12326 = n12202 ^ n12121 ^ x101 ;
  assign n12327 = n12239 ^ n12121 ^ 1'b0 ;
  assign n12328 = ( n12121 & n12326 ) | ( n12121 & ~n12327 ) | ( n12326 & ~n12327 ) ;
  assign n12329 = n12187 ^ n12061 ^ x86 ;
  assign n12330 = n12239 ^ n12061 ^ 1'b0 ;
  assign n12331 = ( n12061 & n12329 ) | ( n12061 & ~n12330 ) | ( n12329 & ~n12330 ) ;
  assign n12332 = n12186 ^ n12064 ^ x85 ;
  assign n12333 = n12239 ^ n12064 ^ 1'b0 ;
  assign n12334 = ( n12064 & n12332 ) | ( n12064 & ~n12333 ) | ( n12332 & ~n12333 ) ;
  assign n12335 = n12185 ^ n12067 ^ x84 ;
  assign n12336 = n12239 ^ n12067 ^ 1'b0 ;
  assign n12337 = ( n12067 & n12335 ) | ( n12067 & ~n12336 ) | ( n12335 & ~n12336 ) ;
  assign n12338 = n12184 ^ n12070 ^ x83 ;
  assign n12339 = n12239 ^ n12070 ^ 1'b0 ;
  assign n12340 = ( n12070 & n12338 ) | ( n12070 & ~n12339 ) | ( n12338 & ~n12339 ) ;
  assign n12341 = n12183 ^ n12073 ^ x82 ;
  assign n12342 = n12239 ^ n12073 ^ 1'b0 ;
  assign n12343 = ( n12073 & n12341 ) | ( n12073 & ~n12342 ) | ( n12341 & ~n12342 ) ;
  assign n12344 = n12182 ^ n12076 ^ x81 ;
  assign n12345 = n12239 ^ n12076 ^ 1'b0 ;
  assign n12346 = ( n12076 & n12344 ) | ( n12076 & ~n12345 ) | ( n12344 & ~n12345 ) ;
  assign n12347 = n12181 ^ n12079 ^ x80 ;
  assign n12348 = n12239 ^ n12079 ^ 1'b0 ;
  assign n12349 = ( n12079 & n12347 ) | ( n12079 & ~n12348 ) | ( n12347 & ~n12348 ) ;
  assign n12350 = n12180 ^ n12007 ^ x79 ;
  assign n12351 = n12239 ^ n12007 ^ 1'b0 ;
  assign n12352 = ( n12007 & n12350 ) | ( n12007 & ~n12351 ) | ( n12350 & ~n12351 ) ;
  assign n12353 = n12179 ^ n12011 ^ x78 ;
  assign n12354 = n12239 ^ n12011 ^ 1'b0 ;
  assign n12355 = ( n12011 & n12353 ) | ( n12011 & ~n12354 ) | ( n12353 & ~n12354 ) ;
  assign n12356 = n12178 ^ n12013 ^ x77 ;
  assign n12357 = n12239 ^ n12013 ^ 1'b0 ;
  assign n12358 = ( n12013 & n12356 ) | ( n12013 & ~n12357 ) | ( n12356 & ~n12357 ) ;
  assign n12359 = n12177 ^ n12015 ^ x76 ;
  assign n12360 = n12239 ^ n12015 ^ 1'b0 ;
  assign n12361 = ( n12015 & n12359 ) | ( n12015 & ~n12360 ) | ( n12359 & ~n12360 ) ;
  assign n12362 = n12176 ^ n12017 ^ x75 ;
  assign n12363 = n12239 ^ n12017 ^ 1'b0 ;
  assign n12364 = ( n12017 & n12362 ) | ( n12017 & ~n12363 ) | ( n12362 & ~n12363 ) ;
  assign n12365 = n12175 ^ n12019 ^ x74 ;
  assign n12366 = n12239 ^ n12019 ^ 1'b0 ;
  assign n12367 = ( n12019 & n12365 ) | ( n12019 & ~n12366 ) | ( n12365 & ~n12366 ) ;
  assign n12368 = n12201 ^ n12124 ^ x100 ;
  assign n12369 = n12239 ^ n12124 ^ 1'b0 ;
  assign n12370 = ( n12124 & n12368 ) | ( n12124 & ~n12369 ) | ( n12368 & ~n12369 ) ;
  assign n12371 = n12200 ^ n12142 ^ x99 ;
  assign n12372 = n12239 ^ n12142 ^ 1'b0 ;
  assign n12373 = ( n12142 & n12371 ) | ( n12142 & ~n12372 ) | ( n12371 & ~n12372 ) ;
  assign n12374 = n12198 ^ n12130 ^ x97 ;
  assign n12375 = n12239 ^ n12130 ^ 1'b0 ;
  assign n12376 = ( n12130 & n12374 ) | ( n12130 & ~n12375 ) | ( n12374 & ~n12375 ) ;
  assign n12377 = n12197 ^ n12133 ^ x96 ;
  assign n12378 = n12239 ^ n12133 ^ 1'b0 ;
  assign n12379 = ( n12133 & n12377 ) | ( n12133 & ~n12378 ) | ( n12377 & ~n12378 ) ;
  assign n12380 = n12196 ^ n12040 ^ x95 ;
  assign n12381 = n12239 ^ n12040 ^ 1'b0 ;
  assign n12382 = ( n12040 & n12380 ) | ( n12040 & ~n12381 ) | ( n12380 & ~n12381 ) ;
  assign n12383 = n12195 ^ n12043 ^ x94 ;
  assign n12384 = n12239 ^ n12043 ^ 1'b0 ;
  assign n12385 = ( n12043 & n12383 ) | ( n12043 & ~n12384 ) | ( n12383 & ~n12384 ) ;
  assign n12386 = n12194 ^ n12046 ^ x93 ;
  assign n12387 = n12239 ^ n12046 ^ 1'b0 ;
  assign n12388 = ( n12046 & n12386 ) | ( n12046 & ~n12387 ) | ( n12386 & ~n12387 ) ;
  assign n12389 = n12193 ^ n12049 ^ x92 ;
  assign n12390 = n12239 ^ n12049 ^ 1'b0 ;
  assign n12391 = ( n12049 & n12389 ) | ( n12049 & ~n12390 ) | ( n12389 & ~n12390 ) ;
  assign n12392 = n12192 ^ n12052 ^ x91 ;
  assign n12393 = n12239 ^ n12052 ^ 1'b0 ;
  assign n12394 = ( n12052 & n12392 ) | ( n12052 & ~n12393 ) | ( n12392 & ~n12393 ) ;
  assign n12395 = n12191 ^ n12055 ^ x90 ;
  assign n12396 = n12239 ^ n12055 ^ 1'b0 ;
  assign n12397 = ( n12055 & n12395 ) | ( n12055 & ~n12396 ) | ( n12395 & ~n12396 ) ;
  assign n12398 = n12190 ^ n12058 ^ x89 ;
  assign n12399 = n12239 ^ n12058 ^ 1'b0 ;
  assign n12400 = ( n12058 & n12398 ) | ( n12058 & ~n12399 ) | ( n12398 & ~n12399 ) ;
  assign n12401 = n12189 ^ n12154 ^ x88 ;
  assign n12402 = n12239 ^ n12154 ^ 1'b0 ;
  assign n12403 = ( n12154 & n12401 ) | ( n12154 & ~n12402 ) | ( n12401 & ~n12402 ) ;
  assign n12404 = n12188 ^ n12147 ^ x87 ;
  assign n12405 = n12239 ^ n12147 ^ 1'b0 ;
  assign n12406 = ( n12147 & n12404 ) | ( n12147 & ~n12405 ) | ( n12404 & ~n12405 ) ;
  assign n12407 = x64 & n12239 ;
  assign n12408 = n12407 ^ x64 ^ x1 ;
  assign n12409 = n12408 ^ n9440 ^ x65 ;
  assign n12410 = ( x65 & n9440 ) | ( x65 & n12409 ) | ( n9440 & n12409 ) ;
  assign n12411 = n12410 ^ n12265 ^ x66 ;
  assign n12412 = ( x66 & n12410 ) | ( x66 & n12411 ) | ( n12410 & n12411 ) ;
  assign n12413 = ( x67 & ~n12258 ) | ( x67 & n12412 ) | ( ~n12258 & n12412 ) ;
  assign n12414 = ( x68 & ~n12253 ) | ( x68 & n12413 ) | ( ~n12253 & n12413 ) ;
  assign n12415 = ( x69 & ~n12262 ) | ( x69 & n12414 ) | ( ~n12262 & n12414 ) ;
  assign n12416 = ( x70 & ~n12271 ) | ( x70 & n12415 ) | ( ~n12271 & n12415 ) ;
  assign n12417 = n12199 ^ n12127 ^ x98 ;
  assign n12418 = n12239 ^ n12127 ^ 1'b0 ;
  assign n12419 = ( x71 & ~n12270 ) | ( x71 & n12416 ) | ( ~n12270 & n12416 ) ;
  assign n12420 = ( x72 & ~n12267 ) | ( x72 & n12419 ) | ( ~n12267 & n12419 ) ;
  assign n12421 = ( x73 & ~n12259 ) | ( x73 & n12420 ) | ( ~n12259 & n12420 ) ;
  assign n12422 = ( x74 & ~n12248 ) | ( x74 & n12421 ) | ( ~n12248 & n12421 ) ;
  assign n12423 = ( x75 & ~n12367 ) | ( x75 & n12422 ) | ( ~n12367 & n12422 ) ;
  assign n12424 = ( x76 & ~n12364 ) | ( x76 & n12423 ) | ( ~n12364 & n12423 ) ;
  assign n12425 = ( x77 & ~n12361 ) | ( x77 & n12424 ) | ( ~n12361 & n12424 ) ;
  assign n12426 = ( x78 & ~n12358 ) | ( x78 & n12425 ) | ( ~n12358 & n12425 ) ;
  assign n12427 = ( x79 & ~n12355 ) | ( x79 & n12426 ) | ( ~n12355 & n12426 ) ;
  assign n12428 = ( x80 & ~n12352 ) | ( x80 & n12427 ) | ( ~n12352 & n12427 ) ;
  assign n12429 = ( x81 & ~n12349 ) | ( x81 & n12428 ) | ( ~n12349 & n12428 ) ;
  assign n12430 = ( x82 & ~n12346 ) | ( x82 & n12429 ) | ( ~n12346 & n12429 ) ;
  assign n12431 = ( x83 & ~n12343 ) | ( x83 & n12430 ) | ( ~n12343 & n12430 ) ;
  assign n12432 = ( x84 & ~n12340 ) | ( x84 & n12431 ) | ( ~n12340 & n12431 ) ;
  assign n12433 = ( x85 & ~n12337 ) | ( x85 & n12432 ) | ( ~n12337 & n12432 ) ;
  assign n12434 = ( x86 & ~n12334 ) | ( x86 & n12433 ) | ( ~n12334 & n12433 ) ;
  assign n12435 = ( x87 & ~n12331 ) | ( x87 & n12434 ) | ( ~n12331 & n12434 ) ;
  assign n12436 = ( x88 & ~n12406 ) | ( x88 & n12435 ) | ( ~n12406 & n12435 ) ;
  assign n12437 = ( x89 & ~n12403 ) | ( x89 & n12436 ) | ( ~n12403 & n12436 ) ;
  assign n12438 = ( x90 & ~n12400 ) | ( x90 & n12437 ) | ( ~n12400 & n12437 ) ;
  assign n12439 = ( x91 & ~n12397 ) | ( x91 & n12438 ) | ( ~n12397 & n12438 ) ;
  assign n12440 = ( x92 & ~n12394 ) | ( x92 & n12439 ) | ( ~n12394 & n12439 ) ;
  assign n12441 = ( x93 & ~n12391 ) | ( x93 & n12440 ) | ( ~n12391 & n12440 ) ;
  assign n12442 = ( x94 & ~n12388 ) | ( x94 & n12441 ) | ( ~n12388 & n12441 ) ;
  assign n12443 = n12442 ^ n12385 ^ x95 ;
  assign n12444 = n12424 ^ n12361 ^ x77 ;
  assign n12445 = n12423 ^ n12364 ^ x76 ;
  assign n12446 = n12422 ^ n12367 ^ x75 ;
  assign n12447 = n12421 ^ n12248 ^ x74 ;
  assign n12448 = n12431 ^ n12340 ^ x84 ;
  assign n12449 = n12420 ^ n12259 ^ x73 ;
  assign n12450 = n12419 ^ n12267 ^ x72 ;
  assign n12451 = n12416 ^ n12270 ^ x71 ;
  assign n12452 = n12415 ^ n12271 ^ x70 ;
  assign n12453 = n12414 ^ n12262 ^ x69 ;
  assign n12454 = n12413 ^ n12253 ^ x68 ;
  assign n12455 = n12412 ^ n12258 ^ x67 ;
  assign n12456 = n12425 ^ n12358 ^ x78 ;
  assign n12457 = n12426 ^ n12355 ^ x79 ;
  assign n12458 = n12427 ^ n12352 ^ x80 ;
  assign n12459 = n12428 ^ n12349 ^ x81 ;
  assign n12460 = n12429 ^ n12346 ^ x82 ;
  assign n12461 = n12430 ^ n12343 ^ x83 ;
  assign n12462 = ( n12127 & n12417 ) | ( n12127 & ~n12418 ) | ( n12417 & ~n12418 ) ;
  assign n12463 = n12432 ^ n12337 ^ x85 ;
  assign n12464 = n12433 ^ n12334 ^ x86 ;
  assign n12465 = n12441 ^ n12388 ^ x94 ;
  assign n12466 = n12435 ^ n12406 ^ x88 ;
  assign n12467 = n12436 ^ n12403 ^ x89 ;
  assign n12468 = n12437 ^ n12400 ^ x90 ;
  assign n12469 = n12438 ^ n12397 ^ x91 ;
  assign n12470 = n12439 ^ n12394 ^ x92 ;
  assign n12471 = n12440 ^ n12391 ^ x93 ;
  assign n12472 = ( x95 & ~n12385 ) | ( x95 & n12442 ) | ( ~n12385 & n12442 ) ;
  assign n12473 = ( x96 & ~n12382 ) | ( x96 & n12472 ) | ( ~n12382 & n12472 ) ;
  assign n12474 = n12472 ^ n12382 ^ x96 ;
  assign n12475 = ( x97 & ~n12379 ) | ( x97 & n12473 ) | ( ~n12379 & n12473 ) ;
  assign n12476 = n12434 ^ n12331 ^ x87 ;
  assign n12477 = ( x98 & ~n12376 ) | ( x98 & n12475 ) | ( ~n12376 & n12475 ) ;
  assign n12478 = ( x99 & ~n12462 ) | ( x99 & n12477 ) | ( ~n12462 & n12477 ) ;
  assign n12479 = ( x100 & ~n12373 ) | ( x100 & n12478 ) | ( ~n12373 & n12478 ) ;
  assign n12480 = ( x101 & ~n12370 ) | ( x101 & n12479 ) | ( ~n12370 & n12479 ) ;
  assign n12481 = ( x102 & ~n12328 ) | ( x102 & n12480 ) | ( ~n12328 & n12480 ) ;
  assign n12482 = ( x103 & ~n12325 ) | ( x103 & n12481 ) | ( ~n12325 & n12481 ) ;
  assign n12483 = ( x104 & ~n12241 ) | ( x104 & n12482 ) | ( ~n12241 & n12482 ) ;
  assign n12484 = ( x105 & ~n12268 ) | ( x105 & n12483 ) | ( ~n12268 & n12483 ) ;
  assign n12485 = ( x106 & ~n12260 ) | ( x106 & n12484 ) | ( ~n12260 & n12484 ) ;
  assign n12486 = ( x107 & ~n12251 ) | ( x107 & n12485 ) | ( ~n12251 & n12485 ) ;
  assign n12487 = ( x108 & ~n12245 ) | ( x108 & n12486 ) | ( ~n12245 & n12486 ) ;
  assign n12488 = ( x109 & ~n12274 ) | ( x109 & n12487 ) | ( ~n12274 & n12487 ) ;
  assign n12489 = ( x110 & ~n12322 ) | ( x110 & n12488 ) | ( ~n12322 & n12488 ) ;
  assign n12490 = ( x111 & ~n12319 ) | ( x111 & n12489 ) | ( ~n12319 & n12489 ) ;
  assign n12491 = ( x112 & ~n12316 ) | ( x112 & n12490 ) | ( ~n12316 & n12490 ) ;
  assign n12492 = ( x113 & ~n12313 ) | ( x113 & n12491 ) | ( ~n12313 & n12491 ) ;
  assign n12493 = ( x114 & ~n12310 ) | ( x114 & n12492 ) | ( ~n12310 & n12492 ) ;
  assign n12494 = ( x115 & ~n12307 ) | ( x115 & n12493 ) | ( ~n12307 & n12493 ) ;
  assign n12495 = ( x116 & ~n12304 ) | ( x116 & n12494 ) | ( ~n12304 & n12494 ) ;
  assign n12496 = ( x117 & ~n12301 ) | ( x117 & n12495 ) | ( ~n12301 & n12495 ) ;
  assign n12497 = ( x118 & ~n12298 ) | ( x118 & n12496 ) | ( ~n12298 & n12496 ) ;
  assign n12498 = ( x119 & ~n12295 ) | ( x119 & n12497 ) | ( ~n12295 & n12497 ) ;
  assign n12499 = ( x120 & ~n12292 ) | ( x120 & n12498 ) | ( ~n12292 & n12498 ) ;
  assign n12500 = ( x121 & ~n12289 ) | ( x121 & n12499 ) | ( ~n12289 & n12499 ) ;
  assign n12501 = ( x122 & ~n12286 ) | ( x122 & n12500 ) | ( ~n12286 & n12500 ) ;
  assign n12502 = ( x123 & ~n12283 ) | ( x123 & n12501 ) | ( ~n12283 & n12501 ) ;
  assign n12503 = ( x124 & ~n12280 ) | ( x124 & n12502 ) | ( ~n12280 & n12502 ) ;
  assign n12504 = ( x125 & ~n12272 ) | ( x125 & n12503 ) | ( ~n12272 & n12503 ) ;
  assign n12505 = ( x126 & ~n12277 ) | ( x126 & n12504 ) | ( ~n12277 & n12504 ) ;
  assign n12506 = ( x127 & ~n12266 ) | ( x127 & n12505 ) | ( ~n12266 & n12505 ) ;
  assign n12507 = ~n12266 & n12506 ;
  assign n12508 = ( n322 & n12506 ) | ( n322 & ~n12507 ) | ( n12506 & ~n12507 ) ;
  assign n12509 = n12506 ^ n12474 ^ 1'b0 ;
  assign n12510 = ( n12382 & n12474 ) | ( n12382 & n12509 ) | ( n12474 & n12509 ) ;
  assign n12511 = n12506 ^ n12443 ^ 1'b0 ;
  assign n12512 = n12506 ^ n12465 ^ 1'b0 ;
  assign n12513 = ( n12388 & n12465 ) | ( n12388 & n12512 ) | ( n12465 & n12512 ) ;
  assign n12514 = n12506 ^ n12469 ^ 1'b0 ;
  assign n12515 = ( n12397 & n12469 ) | ( n12397 & n12514 ) | ( n12469 & n12514 ) ;
  assign n12516 = n12506 ^ n12470 ^ 1'b0 ;
  assign n12517 = n12506 ^ n12467 ^ 1'b0 ;
  assign n12518 = ( n12403 & n12467 ) | ( n12403 & n12517 ) | ( n12467 & n12517 ) ;
  assign n12519 = n12506 ^ n12468 ^ 1'b0 ;
  assign n12520 = n12506 ^ n12455 ^ 1'b0 ;
  assign n12521 = ( n12385 & n12443 ) | ( n12385 & n12511 ) | ( n12443 & n12511 ) ;
  assign n12522 = n12506 ^ n12454 ^ 1'b0 ;
  assign n12523 = ( n12253 & n12454 ) | ( n12253 & n12522 ) | ( n12454 & n12522 ) ;
  assign n12524 = n12506 ^ n12471 ^ 1'b0 ;
  assign n12525 = n12506 ^ n12409 ^ 1'b0 ;
  assign n12526 = n12506 ^ n12411 ^ 1'b0 ;
  assign n12527 = ( n12400 & n12468 ) | ( n12400 & n12519 ) | ( n12468 & n12519 ) ;
  assign n12528 = ( n12265 & n12411 ) | ( n12265 & n12526 ) | ( n12411 & n12526 ) ;
  assign n12529 = ( n12391 & n12471 ) | ( n12391 & n12524 ) | ( n12471 & n12524 ) ;
  assign n12530 = ( n12408 & n12409 ) | ( n12408 & n12525 ) | ( n12409 & n12525 ) ;
  assign n12531 = ( n12258 & n12455 ) | ( n12258 & n12520 ) | ( n12455 & n12520 ) ;
  assign n12532 = ( n12394 & n12470 ) | ( n12394 & n12516 ) | ( n12470 & n12516 ) ;
  assign n12533 = n12506 ^ n12453 ^ 1'b0 ;
  assign n12534 = ( n12262 & n12453 ) | ( n12262 & n12533 ) | ( n12453 & n12533 ) ;
  assign n12535 = n12506 ^ n12452 ^ 1'b0 ;
  assign n12536 = ( n12271 & n12452 ) | ( n12271 & n12535 ) | ( n12452 & n12535 ) ;
  assign n12537 = n12506 ^ n12451 ^ 1'b0 ;
  assign n12538 = ( n12270 & n12451 ) | ( n12270 & n12537 ) | ( n12451 & n12537 ) ;
  assign n12539 = n12506 ^ n12450 ^ 1'b0 ;
  assign n12540 = ( n12267 & n12450 ) | ( n12267 & n12539 ) | ( n12450 & n12539 ) ;
  assign n12541 = n12506 ^ n12449 ^ 1'b0 ;
  assign n12542 = ( n12259 & n12449 ) | ( n12259 & n12541 ) | ( n12449 & n12541 ) ;
  assign n12543 = n12506 ^ n12447 ^ 1'b0 ;
  assign n12544 = ( n12248 & n12447 ) | ( n12248 & n12543 ) | ( n12447 & n12543 ) ;
  assign n12545 = n12506 ^ n12446 ^ 1'b0 ;
  assign n12546 = ( n12367 & n12446 ) | ( n12367 & n12545 ) | ( n12446 & n12545 ) ;
  assign n12547 = n12506 ^ n12445 ^ 1'b0 ;
  assign n12548 = ( n12364 & n12445 ) | ( n12364 & n12547 ) | ( n12445 & n12547 ) ;
  assign n12549 = n12506 ^ n12456 ^ 1'b0 ;
  assign n12550 = ( n12358 & n12456 ) | ( n12358 & n12549 ) | ( n12456 & n12549 ) ;
  assign n12551 = n12506 ^ n12457 ^ 1'b0 ;
  assign n12552 = ( n12355 & n12457 ) | ( n12355 & n12551 ) | ( n12457 & n12551 ) ;
  assign n12553 = n12506 ^ n12458 ^ 1'b0 ;
  assign n12554 = ( n12352 & n12458 ) | ( n12352 & n12553 ) | ( n12458 & n12553 ) ;
  assign n12555 = n12506 ^ n12459 ^ 1'b0 ;
  assign n12556 = ( n12349 & n12459 ) | ( n12349 & n12555 ) | ( n12459 & n12555 ) ;
  assign n12557 = n12506 ^ n12460 ^ 1'b0 ;
  assign n12558 = ( n12346 & n12460 ) | ( n12346 & n12557 ) | ( n12460 & n12557 ) ;
  assign n12559 = n12506 ^ n12461 ^ 1'b0 ;
  assign n12560 = ( n12343 & n12461 ) | ( n12343 & n12559 ) | ( n12461 & n12559 ) ;
  assign n12561 = n12506 ^ n12448 ^ 1'b0 ;
  assign n12562 = n12506 ^ n12444 ^ 1'b0 ;
  assign n12563 = ( n12361 & n12444 ) | ( n12361 & n12562 ) | ( n12444 & n12562 ) ;
  assign n12564 = ( n12340 & n12448 ) | ( n12340 & n12561 ) | ( n12448 & n12561 ) ;
  assign n12565 = n12506 ^ n12463 ^ 1'b0 ;
  assign n12566 = ( n12337 & n12463 ) | ( n12337 & n12565 ) | ( n12463 & n12565 ) ;
  assign n12567 = n12506 ^ n12464 ^ 1'b0 ;
  assign n12568 = ( n12334 & n12464 ) | ( n12334 & n12567 ) | ( n12464 & n12567 ) ;
  assign n12569 = n12506 ^ n12476 ^ 1'b0 ;
  assign n12570 = ( n12331 & n12476 ) | ( n12331 & n12569 ) | ( n12476 & n12569 ) ;
  assign n12571 = n12506 ^ n12466 ^ 1'b0 ;
  assign n12572 = ( n12406 & n12466 ) | ( n12406 & n12571 ) | ( n12466 & n12571 ) ;
  assign n12573 = n12503 ^ n12272 ^ x125 ;
  assign n12574 = n12573 ^ n12506 ^ 1'b0 ;
  assign n12575 = ( n12272 & n12573 ) | ( n12272 & n12574 ) | ( n12573 & n12574 ) ;
  assign n12576 = n12504 ^ n12277 ^ x126 ;
  assign n12577 = n12576 ^ n12506 ^ 1'b0 ;
  assign n12578 = ( n12277 & n12576 ) | ( n12277 & n12577 ) | ( n12576 & n12577 ) ;
  assign n12579 = n12488 ^ n12322 ^ x110 ;
  assign n12580 = n12579 ^ n12506 ^ 1'b0 ;
  assign n12581 = ( n12322 & n12579 ) | ( n12322 & n12580 ) | ( n12579 & n12580 ) ;
  assign n12582 = n12489 ^ n12319 ^ x111 ;
  assign n12583 = n12582 ^ n12506 ^ 1'b0 ;
  assign n12584 = n12490 ^ n12316 ^ x112 ;
  assign n12585 = n12584 ^ n12506 ^ 1'b0 ;
  assign n12586 = ( n12316 & n12584 ) | ( n12316 & n12585 ) | ( n12584 & n12585 ) ;
  assign n12587 = n12491 ^ n12313 ^ x113 ;
  assign n12588 = n12587 ^ n12506 ^ 1'b0 ;
  assign n12589 = ( n12313 & n12587 ) | ( n12313 & n12588 ) | ( n12587 & n12588 ) ;
  assign n12590 = n12492 ^ n12310 ^ x114 ;
  assign n12591 = n12590 ^ n12506 ^ 1'b0 ;
  assign n12592 = ( n12310 & n12590 ) | ( n12310 & n12591 ) | ( n12590 & n12591 ) ;
  assign n12593 = n12493 ^ n12307 ^ x115 ;
  assign n12594 = n12593 ^ n12506 ^ 1'b0 ;
  assign n12595 = ( n12307 & n12593 ) | ( n12307 & n12594 ) | ( n12593 & n12594 ) ;
  assign n12596 = n12494 ^ n12304 ^ x116 ;
  assign n12597 = n12596 ^ n12506 ^ 1'b0 ;
  assign n12598 = ( n12304 & n12596 ) | ( n12304 & n12597 ) | ( n12596 & n12597 ) ;
  assign n12599 = n12495 ^ n12301 ^ x117 ;
  assign n12600 = n12599 ^ n12506 ^ 1'b0 ;
  assign n12601 = ( n12301 & n12599 ) | ( n12301 & n12600 ) | ( n12599 & n12600 ) ;
  assign n12602 = n12496 ^ n12298 ^ x118 ;
  assign n12603 = n12602 ^ n12506 ^ 1'b0 ;
  assign n12604 = ( n12298 & n12602 ) | ( n12298 & n12603 ) | ( n12602 & n12603 ) ;
  assign n12605 = n12497 ^ n12295 ^ x119 ;
  assign n12606 = n12605 ^ n12506 ^ 1'b0 ;
  assign n12607 = ( n12295 & n12605 ) | ( n12295 & n12606 ) | ( n12605 & n12606 ) ;
  assign n12608 = n12498 ^ n12292 ^ x120 ;
  assign n12609 = n12608 ^ n12506 ^ 1'b0 ;
  assign n12610 = ( n12292 & n12608 ) | ( n12292 & n12609 ) | ( n12608 & n12609 ) ;
  assign n12611 = n12499 ^ n12289 ^ x121 ;
  assign n12612 = n12611 ^ n12506 ^ 1'b0 ;
  assign n12613 = ( n12289 & n12611 ) | ( n12289 & n12612 ) | ( n12611 & n12612 ) ;
  assign n12614 = n12500 ^ n12286 ^ x122 ;
  assign n12615 = n12614 ^ n12506 ^ 1'b0 ;
  assign n12616 = ( n12286 & n12614 ) | ( n12286 & n12615 ) | ( n12614 & n12615 ) ;
  assign n12617 = n12501 ^ n12283 ^ x123 ;
  assign n12618 = n12617 ^ n12506 ^ 1'b0 ;
  assign n12619 = ( n12283 & n12617 ) | ( n12283 & n12618 ) | ( n12617 & n12618 ) ;
  assign n12620 = n12502 ^ n12280 ^ x124 ;
  assign n12621 = ( n12319 & n12582 ) | ( n12319 & n12583 ) | ( n12582 & n12583 ) ;
  assign n12622 = n12620 ^ n12506 ^ 1'b0 ;
  assign n12623 = ( n12280 & n12620 ) | ( n12280 & n12622 ) | ( n12620 & n12622 ) ;
  assign n12624 = n12481 ^ n12325 ^ x103 ;
  assign n12625 = n12487 ^ n12274 ^ x109 ;
  assign n12626 = n12473 ^ n12379 ^ x97 ;
  assign n12627 = n12626 ^ n12506 ^ 1'b0 ;
  assign n12628 = ( n12379 & n12626 ) | ( n12379 & n12627 ) | ( n12626 & n12627 ) ;
  assign n12629 = n12624 ^ n12506 ^ 1'b0 ;
  assign n12630 = n12485 ^ n12251 ^ x107 ;
  assign n12631 = n12482 ^ n12241 ^ x104 ;
  assign n12632 = n12475 ^ n12376 ^ x98 ;
  assign n12633 = n12625 ^ n12506 ^ 1'b0 ;
  assign n12634 = n12480 ^ n12328 ^ x102 ;
  assign n12635 = ( n12325 & n12624 ) | ( n12325 & n12629 ) | ( n12624 & n12629 ) ;
  assign n12636 = n12632 ^ n12506 ^ 1'b0 ;
  assign n12637 = ( n12376 & n12632 ) | ( n12376 & n12636 ) | ( n12632 & n12636 ) ;
  assign n12638 = n12634 ^ n12506 ^ 1'b0 ;
  assign n12639 = n12483 ^ n12268 ^ x105 ;
  assign n12640 = n12631 ^ n12506 ^ 1'b0 ;
  assign n12641 = n12630 ^ n12506 ^ 1'b0 ;
  assign n12642 = n12479 ^ n12370 ^ x101 ;
  assign n12643 = ( n12251 & n12630 ) | ( n12251 & n12641 ) | ( n12630 & n12641 ) ;
  assign n12644 = x64 & n12506 ;
  assign n12645 = n12477 ^ n12462 ^ x99 ;
  assign n12646 = n12486 ^ n12245 ^ x108 ;
  assign n12647 = n12642 ^ n12506 ^ 1'b0 ;
  assign n12648 = n12484 ^ n12260 ^ x106 ;
  assign n12649 = ( n12370 & n12642 ) | ( n12370 & n12647 ) | ( n12642 & n12647 ) ;
  assign n12650 = n12646 ^ n12506 ^ 1'b0 ;
  assign n12651 = n12648 ^ n12506 ^ 1'b0 ;
  assign n12652 = ( n12260 & n12648 ) | ( n12260 & n12651 ) | ( n12648 & n12651 ) ;
  assign n12653 = n12645 ^ n12506 ^ 1'b0 ;
  assign n12654 = n12639 ^ n12506 ^ 1'b0 ;
  assign n12655 = n12478 ^ n12373 ^ x100 ;
  assign n12656 = n12655 ^ n12506 ^ 1'b0 ;
  assign n12657 = ( n12274 & n12625 ) | ( n12274 & n12633 ) | ( n12625 & n12633 ) ;
  assign n12658 = ( n12328 & n12634 ) | ( n12328 & n12638 ) | ( n12634 & n12638 ) ;
  assign n12659 = ( n12373 & n12655 ) | ( n12373 & n12656 ) | ( n12655 & n12656 ) ;
  assign n12660 = ( n12245 & n12646 ) | ( n12245 & n12650 ) | ( n12646 & n12650 ) ;
  assign n12661 = ( n12462 & n12645 ) | ( n12462 & n12653 ) | ( n12645 & n12653 ) ;
  assign n12662 = n12644 ^ x64 ^ x0 ;
  assign n12663 = ( n12241 & n12631 ) | ( n12241 & n12640 ) | ( n12631 & n12640 ) ;
  assign n12664 = ( n12268 & n12639 ) | ( n12268 & n12654 ) | ( n12639 & n12654 ) ;
  assign y0 = ~n9628 ;
  assign y1 = ~n9396 ;
  assign y2 = ~n9135 ;
  assign y3 = ~n8900 ;
  assign y4 = ~n8653 ;
  assign y5 = ~n8410 ;
  assign y6 = ~n8172 ;
  assign y7 = ~n7944 ;
  assign y8 = ~n7723 ;
  assign y9 = ~n7480 ;
  assign y10 = ~n7258 ;
  assign y11 = ~n7044 ;
  assign y12 = ~n6829 ;
  assign y13 = ~n6621 ;
  assign y14 = ~n6212 ;
  assign y15 = ~n6006 ;
  assign y16 = ~n5410 ;
  assign y17 = ~n4950 ;
  assign y18 = ~n4733 ;
  assign y19 = ~n4540 ;
  assign y20 = ~n4360 ;
  assign y21 = ~n4180 ;
  assign y22 = ~n4012 ;
  assign y23 = ~n3837 ;
  assign y24 = ~n3662 ;
  assign y25 = ~n3506 ;
  assign y26 = ~n3340 ;
  assign y27 = ~n3182 ;
  assign y28 = ~n3051 ;
  assign y29 = ~n2900 ;
  assign y30 = ~n2746 ;
  assign y31 = ~n2623 ;
  assign y32 = ~n2482 ;
  assign y33 = ~n2345 ;
  assign y34 = ~n2237 ;
  assign y35 = ~n2106 ;
  assign y36 = ~n1985 ;
  assign y37 = ~n1885 ;
  assign y38 = ~n1765 ;
  assign y39 = ~n1653 ;
  assign y40 = ~n1554 ;
  assign y41 = ~n1449 ;
  assign y42 = ~n1359 ;
  assign y43 = ~n1266 ;
  assign y44 = ~n1175 ;
  assign y45 = ~n1095 ;
  assign y46 = ~n1021 ;
  assign y47 = ~n942 ;
  assign y48 = ~n872 ;
  assign y49 = ~n817 ;
  assign y50 = ~n744 ;
  assign y51 = ~n686 ;
  assign y52 = ~n635 ;
  assign y53 = ~n585 ;
  assign y54 = ~n539 ;
  assign y55 = ~n497 ;
  assign y56 = ~n452 ;
  assign y57 = ~n422 ;
  assign y58 = ~n396 ;
  assign y59 = ~n353 ;
  assign y60 = ~n314 ;
  assign y61 = ~n282 ;
  assign y62 = ~n279 ;
  assign y63 = ~n305 ;
  assign y64 = n12662 ;
  assign y65 = n12530 ;
  assign y66 = n12528 ;
  assign y67 = n12531 ;
  assign y68 = n12523 ;
  assign y69 = n12534 ;
  assign y70 = n12536 ;
  assign y71 = n12538 ;
  assign y72 = n12540 ;
  assign y73 = n12542 ;
  assign y74 = n12544 ;
  assign y75 = n12546 ;
  assign y76 = n12548 ;
  assign y77 = n12563 ;
  assign y78 = n12550 ;
  assign y79 = n12552 ;
  assign y80 = n12554 ;
  assign y81 = n12556 ;
  assign y82 = n12558 ;
  assign y83 = n12560 ;
  assign y84 = n12564 ;
  assign y85 = n12566 ;
  assign y86 = n12568 ;
  assign y87 = n12570 ;
  assign y88 = n12572 ;
  assign y89 = n12518 ;
  assign y90 = n12527 ;
  assign y91 = n12515 ;
  assign y92 = n12532 ;
  assign y93 = n12529 ;
  assign y94 = n12513 ;
  assign y95 = n12521 ;
  assign y96 = n12510 ;
  assign y97 = n12628 ;
  assign y98 = n12637 ;
  assign y99 = n12661 ;
  assign y100 = n12659 ;
  assign y101 = n12649 ;
  assign y102 = n12658 ;
  assign y103 = n12635 ;
  assign y104 = n12663 ;
  assign y105 = n12664 ;
  assign y106 = n12652 ;
  assign y107 = n12643 ;
  assign y108 = n12660 ;
  assign y109 = n12657 ;
  assign y110 = n12581 ;
  assign y111 = n12621 ;
  assign y112 = n12586 ;
  assign y113 = n12589 ;
  assign y114 = n12592 ;
  assign y115 = n12595 ;
  assign y116 = n12598 ;
  assign y117 = n12601 ;
  assign y118 = n12604 ;
  assign y119 = n12607 ;
  assign y120 = n12610 ;
  assign y121 = n12613 ;
  assign y122 = n12616 ;
  assign y123 = n12619 ;
  assign y124 = n12623 ;
  assign y125 = n12575 ;
  assign y126 = n12578 ;
  assign y127 = n12508 ;
endmodule
