module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 ;
  assign n33 = x23 & ~x26 ;
  assign n34 = ~x29 & x30 ;
  assign n35 = x27 & x28 ;
  assign n36 = x29 & x30 ;
  assign n37 = x29 & ~x30 ;
  assign n38 = x24 & ~x25 ;
  assign n39 = ~x27 & x28 ;
  assign n40 = x24 | x25 ;
  assign n41 = x27 | x28 ;
  assign n42 = x23 | x26 ;
  assign n43 = x24 & x25 ;
  assign n44 = ~x23 & x26 ;
  assign n45 = n33 & n43 ;
  assign n46 = n34 & ~n41 ;
  assign n47 = n40 | n42 ;
  assign n48 = x29 | x30 ;
  assign n49 = n35 & n37 ;
  assign n50 = ~x24 & x25 ;
  assign n51 = n39 & ~n48 ;
  assign n52 = n35 & ~n48 ;
  assign n53 = ~n42 & n50 ;
  assign n54 = x23 & x26 ;
  assign n55 = ~n40 & n54 ;
  assign n56 = n35 & n36 ;
  assign n57 = n43 & n54 ;
  assign n58 = n33 & n50 ;
  assign n59 = n37 & ~n41 ;
  assign n60 = n38 & n44 ;
  assign n61 = n36 & n39 ;
  assign n62 = n33 & n38 ;
  assign n63 = ~n42 & n43 ;
  assign n64 = n38 & n54 ;
  assign n65 = n37 & n39 ;
  assign n66 = n33 & ~n40 ;
  assign n67 = n41 | n48 ;
  assign n68 = x27 & ~x28 ;
  assign n69 = n38 & ~n42 ;
  assign n70 = n34 & n39 ;
  assign n71 = n36 & ~n41 ;
  assign n72 = n50 & n54 ;
  assign n73 = n44 & n50 ;
  assign n74 = n34 & n35 ;
  assign n75 = ~n48 & n68 ;
  assign n76 = ~n40 & n44 ;
  assign n77 = n34 & n68 ;
  assign n78 = n37 & n68 ;
  assign n79 = n36 & n68 ;
  assign n80 = n43 & n44 ;
  assign n81 = n58 & n70 ;
  assign n82 = n64 & n70 ;
  assign n83 = n66 & n74 ;
  assign n84 = n63 & n70 ;
  assign n85 = n82 | n84 ;
  assign n86 = n53 & n70 ;
  assign n87 = n58 & n65 ;
  assign n88 = ~n47 & n51 ;
  assign n89 = n63 & n78 ;
  assign n90 = n51 & n73 ;
  assign n91 = n62 & n70 ;
  assign n92 = n60 & n70 ;
  assign n93 = n70 & n76 ;
  assign n94 = n45 & n77 ;
  assign n95 = n46 & n53 ;
  assign n96 = n60 & n61 ;
  assign n97 = n55 & n70 ;
  assign n98 = n70 & n80 ;
  assign n99 = n86 | n95 ;
  assign n100 = n57 & ~n67 ;
  assign n101 = n61 & n64 ;
  assign n102 = ~n67 & n76 ;
  assign n103 = n79 & n80 ;
  assign n104 = n93 | n98 ;
  assign n105 = n46 & n64 ;
  assign n106 = n93 | n105 ;
  assign n107 = n49 & n63 ;
  assign n108 = n92 | n97 ;
  assign n109 = n70 & n72 ;
  assign n110 = n81 | n109 ;
  assign n111 = ~n67 & n73 ;
  assign n112 = n102 | n107 ;
  assign n113 = n85 | n110 ;
  assign n114 = n104 | n113 ;
  assign n115 = n83 | n114 ;
  assign n116 = n64 & n79 ;
  assign n117 = n112 | n116 ;
  assign n118 = n99 | n117 ;
  assign n119 = n101 | n111 ;
  assign n120 = ( ~n106 & n118 ) | ( ~n106 & n119 ) | ( n118 & n119 ) ;
  assign n121 = n106 | n120 ;
  assign n122 = n62 & n78 ;
  assign n123 = n88 | n121 ;
  assign n124 = n75 & n80 ;
  assign n125 = n55 & n77 ;
  assign n126 = n124 | n125 ;
  assign n127 = n84 | n103 ;
  assign n128 = n45 & n71 ;
  assign n129 = n94 | n100 ;
  assign n130 = n108 | n129 ;
  assign n131 = n94 | n128 ;
  assign n132 = n117 | n126 ;
  assign n133 = n74 & n80 ;
  assign n134 = n127 | n132 ;
  assign n135 = n91 | n133 ;
  assign n136 = n131 | n135 ;
  assign n137 = n90 | n96 ;
  assign n138 = n136 | n137 ;
  assign n139 = n52 & n62 ;
  assign n140 = ( ~n89 & n134 ) | ( ~n89 & n139 ) | ( n134 & n139 ) ;
  assign n141 = n89 | n140 ;
  assign n142 = ( ~n87 & n122 ) | ( ~n87 & n138 ) | ( n122 & n138 ) ;
  assign n143 = n87 | n142 ;
  assign n144 = n46 & n80 ;
  assign n145 = n55 & n56 ;
  assign n146 = n60 & n65 ;
  assign n147 = n56 & n63 ;
  assign n148 = ~n67 & n72 ;
  assign n149 = n57 & n79 ;
  assign n150 = n73 & n74 ;
  assign n151 = n93 | n146 ;
  assign n152 = n97 | n150 ;
  assign n153 = n46 & n76 ;
  assign n154 = n72 & n74 ;
  assign n155 = n144 | n153 ;
  assign n156 = n149 | n155 ;
  assign n157 = n98 | n154 ;
  assign n158 = n156 | n157 ;
  assign n159 = n96 | n152 ;
  assign n160 = n158 | n159 ;
  assign n161 = n57 & n77 ;
  assign n162 = n66 & n75 ;
  assign n163 = n161 | n162 ;
  assign n164 = n66 & ~n67 ;
  assign n165 = n63 & n77 ;
  assign n166 = n152 | n163 ;
  assign n167 = n53 & n75 ;
  assign n168 = n73 & n75 ;
  assign n169 = n56 & n69 ;
  assign n170 = n165 | n169 ;
  assign n171 = n130 | n170 ;
  assign n172 = n72 & n75 ;
  assign n173 = n58 & n71 ;
  assign n174 = n172 | n173 ;
  assign n175 = n51 & n55 ;
  assign n176 = n124 | n168 ;
  assign n177 = n45 & n78 ;
  assign n178 = ( ~n164 & n171 ) | ( ~n164 & n177 ) | ( n171 & n177 ) ;
  assign n179 = n101 | n177 ;
  assign n180 = n145 | n175 ;
  assign n181 = n164 | n178 ;
  assign n182 = n73 & n78 ;
  assign n183 = n53 & n61 ;
  assign n184 = n53 & n56 ;
  assign n185 = ( ~n147 & n160 ) | ( ~n147 & n184 ) | ( n160 & n184 ) ;
  assign n186 = n147 | n185 ;
  assign n187 = n59 & n66 ;
  assign n188 = n78 & n80 ;
  assign n189 = ( n148 & ~n168 ) | ( n148 & n186 ) | ( ~n168 & n186 ) ;
  assign n190 = n168 | n189 ;
  assign n191 = n162 | n179 ;
  assign n192 = n174 | n191 ;
  assign n193 = n180 | n183 ;
  assign n194 = n192 | n193 ;
  assign n195 = n175 | n187 ;
  assign n196 = n176 | n195 ;
  assign n197 = ~n47 & n52 ;
  assign n198 = ( ~n182 & n188 ) | ( ~n182 & n190 ) | ( n188 & n190 ) ;
  assign n199 = n191 | n196 ;
  assign n200 = ( n167 & n194 ) | ( n167 & ~n197 ) | ( n194 & ~n197 ) ;
  assign n201 = n182 | n198 ;
  assign n202 = n151 | n166 ;
  assign n203 = n59 & n63 ;
  assign n204 = n181 | n203 ;
  assign n205 = n197 | n200 ;
  assign n206 = n49 & n64 ;
  assign n207 = n66 & n77 ;
  assign n208 = n91 | n206 ;
  assign n209 = n51 & n62 ;
  assign n210 = n51 & n60 ;
  assign n211 = n72 & n77 ;
  assign n212 = n69 & n74 ;
  assign n213 = n100 | n167 ;
  assign n214 = n61 & n72 ;
  assign n215 = n197 | n214 ;
  assign n216 = n211 | n213 ;
  assign n217 = n207 | n210 ;
  assign n218 = n91 | n212 ;
  assign n219 = n65 & n73 ;
  assign n220 = n61 & n62 ;
  assign n221 = n53 & n71 ;
  assign n222 = n52 & n73 ;
  assign n223 = n214 | n219 ;
  assign n224 = n64 & n74 ;
  assign n225 = n64 & n77 ;
  assign n226 = n83 | n224 ;
  assign n227 = n133 | n225 ;
  assign n228 = ~n47 & n77 ;
  assign n229 = n63 & n74 ;
  assign n230 = n223 | n226 ;
  assign n231 = ~n47 & n49 ;
  assign n232 = n52 & n80 ;
  assign n233 = n211 | n228 ;
  assign n234 = n46 & n72 ;
  assign n235 = n45 & n51 ;
  assign n236 = n168 | n217 ;
  assign n237 = n229 | n231 ;
  assign n238 = n209 | n235 ;
  assign n239 = n208 | n238 ;
  assign n240 = n234 | n239 ;
  assign n241 = n63 & n71 ;
  assign n242 = n215 | n241 ;
  assign n243 = n227 | n242 ;
  assign n244 = n236 | n243 ;
  assign n245 = n49 & n73 ;
  assign n246 = n60 & n77 ;
  assign n247 = n52 & n76 ;
  assign n248 = n56 & n62 ;
  assign n249 = n201 | n245 ;
  assign n250 = n58 & n61 ;
  assign n251 = n211 | n246 ;
  assign n252 = ( n222 & ~n232 ) | ( n222 & n244 ) | ( ~n232 & n244 ) ;
  assign n253 = n233 | n240 ;
  assign n254 = n232 | n252 ;
  assign n255 = n58 & n77 ;
  assign n256 = n237 | n255 ;
  assign n257 = n242 | n256 ;
  assign n258 = n45 & n46 ;
  assign n259 = n216 | n245 ;
  assign n260 = n218 | n259 ;
  assign n261 = n250 | n258 ;
  assign n262 = n230 | n261 ;
  assign n263 = ( ~n167 & n221 ) | ( ~n167 & n262 ) | ( n221 & n262 ) ;
  assign n264 = n167 | n263 ;
  assign n265 = n253 | n257 ;
  assign n266 = ( n103 & ~n220 ) | ( n103 & n265 ) | ( ~n220 & n265 ) ;
  assign n267 = n220 | n266 ;
  assign n268 = ( n247 & ~n248 ) | ( n247 & n267 ) | ( ~n248 & n267 ) ;
  assign n269 = n248 | n268 ;
  assign n270 = n187 | n269 ;
  assign n271 = n49 & n72 ;
  assign n272 = n103 | n271 ;
  assign n273 = n251 | n258 ;
  assign n274 = n272 | n273 ;
  assign n275 = n148 | n264 ;
  assign n276 = n51 & n57 ;
  assign n277 = ( n87 & n254 ) | ( n87 & ~n276 ) | ( n254 & ~n276 ) ;
  assign n278 = n276 | n277 ;
  assign n279 = n55 & ~n67 ;
  assign n280 = n133 | n279 ;
  assign n281 = n45 & n70 ;
  assign n282 = n57 & n70 ;
  assign n283 = n62 & n74 ;
  assign n284 = n165 | n255 ;
  assign n285 = n97 | n207 ;
  assign n286 = n70 & n73 ;
  assign n287 = n45 & n74 ;
  assign n288 = n62 & n77 ;
  assign n289 = n66 & n70 ;
  assign n290 = n55 & n74 ;
  assign n291 = n225 | n289 ;
  assign n292 = n100 | n169 ;
  assign n293 = n76 & n77 ;
  assign n294 = n53 & n77 ;
  assign n295 = n73 & n77 ;
  assign n296 = ~n47 & n70 ;
  assign n297 = n211 | n288 ;
  assign n298 = n294 | n297 ;
  assign n299 = ~n55 & n77 ;
  assign n300 = n58 & n74 ;
  assign n301 = n161 | n295 ;
  assign n302 = ~n47 & n74 ;
  assign n303 = n60 & n74 ;
  assign n304 = n77 & n80 ;
  assign n305 = n229 | n300 ;
  assign n306 = n74 & n76 ;
  assign n307 = n94 | n296 ;
  assign n308 = n293 | n301 ;
  assign n309 = n280 | n298 ;
  assign n310 = n285 | n302 ;
  assign n311 = n307 | n308 ;
  assign n312 = n290 | n306 ;
  assign n313 = n69 & n70 ;
  assign n314 = n305 | n312 ;
  assign n315 = n291 | n311 ;
  assign n316 = n284 | n298 ;
  assign n317 = n315 | n316 ;
  assign n318 = n69 & n77 ;
  assign n319 = ( n246 & n304 ) | ( n246 & ~n317 ) | ( n304 & ~n317 ) ;
  assign n320 = n317 | n319 ;
  assign n321 = ( n77 & ~n299 ) | ( n77 & n320 ) | ( ~n299 & n320 ) ;
  assign n322 = n91 | n313 ;
  assign n323 = n92 | n282 ;
  assign n324 = n310 | n314 ;
  assign n325 = n280 | n292 ;
  assign n326 = n322 | n324 ;
  assign n327 = n286 | n323 ;
  assign n328 = n115 | n327 ;
  assign n329 = n321 | n328 ;
  assign n330 = n326 | n329 ;
  assign n331 = ( ~n86 & n281 ) | ( ~n86 & n330 ) | ( n281 & n330 ) ;
  assign n332 = n53 & n74 ;
  assign n333 = n86 | n331 ;
  assign n334 = ( ~n303 & n332 ) | ( ~n303 & n333 ) | ( n332 & n333 ) ;
  assign n335 = n303 | n334 ;
  assign n336 = n57 & n74 ;
  assign n337 = ( ~n212 & n283 ) | ( ~n212 & n335 ) | ( n283 & n335 ) ;
  assign n338 = n212 | n337 ;
  assign n339 = ( n287 & ~n318 ) | ( n287 & n338 ) | ( ~n318 & n338 ) ;
  assign n340 = n318 | n339 ;
  assign n341 = n61 & n66 ;
  assign n342 = n46 & n58 ;
  assign n343 = n55 & n59 ;
  assign n344 = n145 | n343 ;
  assign n345 = n52 & n63 ;
  assign n346 = n161 | n345 ;
  assign n347 = n83 | n168 ;
  assign n348 = n72 & n79 ;
  assign n349 = n66 & n71 ;
  assign n350 = n341 | n342 ;
  assign n351 = n51 & n76 ;
  assign n352 = ~n47 & n61 ;
  assign n353 = n348 | n349 ;
  assign n354 = n184 | n350 ;
  assign n355 = n295 | n306 ;
  assign n356 = n102 | n250 ;
  assign n357 = n51 & n63 ;
  assign n358 = n51 & n64 ;
  assign n359 = n212 | n356 ;
  assign n360 = n51 & n53 ;
  assign n361 = n357 | n360 ;
  assign n362 = n52 & n72 ;
  assign n363 = n344 | n361 ;
  assign n364 = n346 | n353 ;
  assign n365 = n363 | n364 ;
  assign n366 = n147 | n352 ;
  assign n367 = n51 & n80 ;
  assign n368 = ( ~n362 & n365 ) | ( ~n362 & n367 ) | ( n365 & n367 ) ;
  assign n369 = n153 | n172 ;
  assign n370 = n246 | n342 ;
  assign n371 = n53 & ~n67 ;
  assign n372 = n49 & n53 ;
  assign n373 = n46 & n66 ;
  assign n374 = n372 | n373 ;
  assign n375 = n56 & n64 ;
  assign n376 = n351 | n375 ;
  assign n377 = n358 | n376 ;
  assign n378 = n63 & n65 ;
  assign n379 = n88 | n281 ;
  assign n380 = n370 | n379 ;
  assign n381 = n49 & n69 ;
  assign n382 = n362 | n368 ;
  assign n383 = n214 | n381 ;
  assign n384 = n128 | n372 ;
  assign n385 = n371 | n383 ;
  assign n386 = n283 | n384 ;
  assign n387 = n347 | n386 ;
  assign n388 = n361 | n386 ;
  assign n389 = n369 | n381 ;
  assign n390 = n248 | n366 ;
  assign n391 = n308 | n390 ;
  assign n392 = n374 | n389 ;
  assign n393 = n312 | n385 ;
  assign n394 = n354 | n388 ;
  assign n395 = n86 | n98 ;
  assign n396 = n391 | n394 ;
  assign n397 = ~n47 & n75 ;
  assign n398 = n355 | n385 ;
  assign n399 = n395 | n398 ;
  assign n400 = n49 & n76 ;
  assign n401 = n332 | n344 ;
  assign n402 = n359 | n377 ;
  assign n403 = n401 | n402 ;
  assign n404 = ( n103 & ~n362 ) | ( n103 & n403 ) | ( ~n362 & n403 ) ;
  assign n405 = n362 | n404 ;
  assign n406 = ( ~n100 & n378 ) | ( ~n100 & n405 ) | ( n378 & n405 ) ;
  assign n407 = n100 | n406 ;
  assign n408 = ( n345 & ~n397 ) | ( n345 & n399 ) | ( ~n397 & n399 ) ;
  assign n409 = n397 | n408 ;
  assign n410 = n59 & n73 ;
  assign n411 = ( ~n400 & n407 ) | ( ~n400 & n410 ) | ( n407 & n410 ) ;
  assign n412 = n400 | n411 ;
  assign n413 = n206 | n412 ;
  assign n414 = n65 & n66 ;
  assign n415 = n62 & n71 ;
  assign n416 = n62 & ~n67 ;
  assign n417 = ~n47 & n56 ;
  assign n418 = n283 | n360 ;
  assign n419 = n212 | n294 ;
  assign n420 = n56 & n76 ;
  assign n421 = n294 | n420 ;
  assign n422 = n57 & n61 ;
  assign n423 = n66 & n79 ;
  assign n424 = n83 | n422 ;
  assign n425 = n65 & n76 ;
  assign n426 = n45 & n65 ;
  assign n427 = n57 & n59 ;
  assign n428 = n423 | n427 ;
  assign n429 = n109 | n241 ;
  assign n430 = n92 | n283 ;
  assign n431 = n349 | n424 ;
  assign n432 = n429 | n431 ;
  assign n433 = n75 & n76 ;
  assign n434 = n65 & n72 ;
  assign n435 = n281 | n434 ;
  assign n436 = n362 | n435 ;
  assign n437 = n46 & n73 ;
  assign n438 = n290 | n397 ;
  assign n439 = n87 | n437 ;
  assign n440 = n84 | n439 ;
  assign n441 = n221 | n422 ;
  assign n442 = n64 & n75 ;
  assign n443 = n415 | n423 ;
  assign n444 = n45 & n49 ;
  assign n445 = n207 | n437 ;
  assign n446 = n443 | n445 ;
  assign n447 = ~n47 & n79 ;
  assign n448 = n63 & n75 ;
  assign n449 = n414 | n448 ;
  assign n450 = n419 | n447 ;
  assign n451 = n441 | n449 ;
  assign n452 = n421 | n446 ;
  assign n453 = ( n167 & ~n232 ) | ( n167 & n452 ) | ( ~n232 & n452 ) ;
  assign n454 = n232 | n453 ;
  assign n455 = n444 | n447 ;
  assign n456 = n279 | n454 ;
  assign n457 = n418 | n428 ;
  assign n458 = n184 | n433 ;
  assign n459 = n457 | n458 ;
  assign n460 = n450 | n459 ;
  assign n461 = n55 & n71 ;
  assign n462 = n442 | n460 ;
  assign n463 = n438 | n451 ;
  assign n464 = n462 | n463 ;
  assign n465 = n440 | n464 ;
  assign n466 = n88 | n461 ;
  assign n467 = n387 | n455 ;
  assign n468 = n57 & n78 ;
  assign n469 = n392 | n436 ;
  assign n470 = n465 | n469 ;
  assign n471 = ( n103 & ~n296 ) | ( n103 & n470 ) | ( ~n296 & n470 ) ;
  assign n472 = n296 | n471 ;
  assign n473 = n434 | n447 ;
  assign n474 = n430 | n473 ;
  assign n475 = n466 | n474 ;
  assign n476 = n51 & n72 ;
  assign n477 = ( n209 & ~n468 ) | ( n209 & n475 ) | ( ~n468 & n475 ) ;
  assign n478 = n468 | n477 ;
  assign n479 = ( ~n414 & n425 ) | ( ~n414 & n478 ) | ( n425 & n478 ) ;
  assign n480 = n414 | n479 ;
  assign n481 = ( n417 & ~n420 ) | ( n417 & n472 ) | ( ~n420 & n472 ) ;
  assign n482 = n420 | n481 ;
  assign n483 = ( n416 & ~n476 ) | ( n416 & n482 ) | ( ~n476 & n482 ) ;
  assign n484 = n476 | n483 ;
  assign n485 = ( n426 & ~n468 ) | ( n426 & n484 ) | ( ~n468 & n484 ) ;
  assign n486 = n468 | n485 ;
  assign n487 = n203 | n486 ;
  assign n488 = n239 | n487 ;
  assign n489 = n59 & n76 ;
  assign n490 = n46 & n62 ;
  assign n491 = n332 | n490 ;
  assign n492 = n213 | n416 ;
  assign n493 = n341 | n447 ;
  assign n494 = n255 | n447 ;
  assign n495 = n101 | n491 ;
  assign n496 = n107 | n489 ;
  assign n497 = n45 & n52 ;
  assign n498 = n281 | n494 ;
  assign n499 = n61 & n76 ;
  assign n500 = n497 | n499 ;
  assign n501 = n53 & n59 ;
  assign n502 = n69 & n71 ;
  assign n503 = n53 & n79 ;
  assign n504 = n154 | n502 ;
  assign n505 = n493 | n504 ;
  assign n506 = n351 | n503 ;
  assign n507 = n492 | n498 ;
  assign n508 = n449 | n500 ;
  assign n509 = n505 | n508 ;
  assign n510 = n60 & n79 ;
  assign n511 = ( n167 & ~n420 ) | ( n167 & n509 ) | ( ~n420 & n509 ) ;
  assign n512 = n506 | n510 ;
  assign n513 = n495 | n507 ;
  assign n514 = n358 | n423 ;
  assign n515 = ( ~n276 & n358 ) | ( ~n276 & n513 ) | ( n358 & n513 ) ;
  assign n516 = n276 | n515 ;
  assign n517 = n496 | n514 ;
  assign n518 = n498 | n512 ;
  assign n519 = n432 | n518 ;
  assign n520 = n76 & n79 ;
  assign n521 = n420 | n511 ;
  assign n522 = n55 & n75 ;
  assign n523 = ( n248 & n519 ) | ( n248 & ~n520 ) | ( n519 & ~n520 ) ;
  assign n524 = n520 | n523 ;
  assign n525 = ( ~n427 & n501 ) | ( ~n427 & n524 ) | ( n501 & n524 ) ;
  assign n526 = ( n124 & n521 ) | ( n124 & ~n522 ) | ( n521 & ~n522 ) ;
  assign n527 = n480 | n512 ;
  assign n528 = n427 | n525 ;
  assign n529 = n522 | n526 ;
  assign n530 = n49 & n60 ;
  assign n531 = n139 | n530 ;
  assign n532 = n61 & n73 ;
  assign n533 = n231 | n532 ;
  assign n534 = n71 & n76 ;
  assign n535 = n286 | n332 ;
  assign n536 = n313 | n410 ;
  assign n537 = n224 | n358 ;
  assign n538 = n188 | n224 ;
  assign n539 = n182 | n289 ;
  assign n540 = n536 | n537 ;
  assign n541 = n535 | n540 ;
  assign n542 = n439 | n539 ;
  assign n543 = n541 | n542 ;
  assign n544 = n531 | n539 ;
  assign n545 = n533 | n544 ;
  assign n546 = n61 & n80 ;
  assign n547 = n69 & n79 ;
  assign n548 = n222 | n546 ;
  assign n549 = n547 | n548 ;
  assign n550 = n241 | n420 ;
  assign n551 = n196 | n550 ;
  assign n552 = n52 & n58 ;
  assign n553 = n219 | n425 ;
  assign n554 = n549 | n551 ;
  assign n555 = n58 & n59 ;
  assign n556 = n545 | n554 ;
  assign n557 = n423 | n552 ;
  assign n558 = ( ~n209 & n534 ) | ( ~n209 & n543 ) | ( n534 & n543 ) ;
  assign n559 = n76 & n78 ;
  assign n560 = n336 | n559 ;
  assign n561 = n109 | n144 ;
  assign n562 = ( ~n184 & n271 ) | ( ~n184 & n556 ) | ( n271 & n556 ) ;
  assign n563 = n209 | n558 ;
  assign n564 = n538 | n560 ;
  assign n565 = n203 | n522 ;
  assign n566 = n396 | n562 ;
  assign n567 = n184 | n562 ;
  assign n568 = ( n557 & ~n565 ) | ( n557 & n566 ) | ( ~n565 & n566 ) ;
  assign n569 = n565 | n568 ;
  assign n570 = ( ~n553 & n561 ) | ( ~n553 & n569 ) | ( n561 & n569 ) ;
  assign n571 = n553 | n570 ;
  assign n572 = ( ~n302 & n502 ) | ( ~n302 & n571 ) | ( n502 & n571 ) ;
  assign n573 = n302 | n572 ;
  assign n574 = ( n169 & ~n197 ) | ( n169 & n573 ) | ( ~n197 & n573 ) ;
  assign n575 = n197 | n574 ;
  assign n576 = n555 | n575 ;
  assign n577 = n463 | n576 ;
  assign n578 = n66 & n78 ;
  assign n579 = n98 | n578 ;
  assign n580 = ~n47 & n59 ;
  assign n581 = n539 | n579 ;
  assign n582 = n303 | n580 ;
  assign n583 = n47 | n67 ;
  assign n584 = ~n246 & n583 ;
  assign n585 = n55 & n61 ;
  assign n586 = n183 | n585 ;
  assign n587 = n229 | n345 ;
  assign n588 = n352 | n499 ;
  assign n589 = ~n47 & n78 ;
  assign n590 = n149 | n220 ;
  assign n591 = n56 & n72 ;
  assign n592 = n60 & n71 ;
  assign n593 = n61 & n63 ;
  assign n594 = n90 | n351 ;
  assign n595 = n349 | n547 ;
  assign n596 = n593 | n595 ;
  assign n597 = n103 | n587 ;
  assign n598 = n584 & ~n597 ;
  assign n599 = ~n293 & n598 ;
  assign n600 = n60 & n78 ;
  assign n601 = n49 & n55 ;
  assign n602 = n45 & n61 ;
  assign n603 = ~n581 & n599 ;
  assign n604 = n591 | n592 ;
  assign n605 = n56 & n80 ;
  assign n606 = ~n409 & n583 ;
  assign n607 = n46 & ~n47 ;
  assign n608 = n57 & n65 ;
  assign n609 = ( n516 & n589 ) | ( n516 & ~n600 ) | ( n589 & ~n600 ) ;
  assign n610 = n586 | n588 ;
  assign n611 = n309 | n604 ;
  assign n612 = n45 & n75 ;
  assign n613 = n582 | n586 ;
  assign n614 = n603 & ~n613 ;
  assign n615 = n600 | n609 ;
  assign n616 = n281 | n489 ;
  assign n617 = n590 | n610 ;
  assign n618 = n290 | n607 ;
  assign n619 = n94 | n618 ;
  assign n620 = n596 | n619 ;
  assign n621 = n546 | n605 ;
  assign n622 = ( ~n219 & n601 ) | ( ~n219 & n615 ) | ( n601 & n615 ) ;
  assign n623 = n612 | n616 ;
  assign n624 = n594 | n623 ;
  assign n625 = n532 | n591 ;
  assign n626 = n145 | n625 ;
  assign n627 = n621 | n626 ;
  assign n628 = n58 & n78 ;
  assign n629 = n219 | n622 ;
  assign n630 = ( ~n375 & n608 ) | ( ~n375 & n620 ) | ( n608 & n620 ) ;
  assign n631 = n61 & n69 ;
  assign n632 = n375 | n630 ;
  assign n633 = ( n382 & ~n578 ) | ( n382 & n628 ) | ( ~n578 & n628 ) ;
  assign n634 = n601 | n632 ;
  assign n635 = ( n358 & ~n426 ) | ( n358 & n614 ) | ( ~n426 & n614 ) ;
  assign n636 = ~n358 & n635 ;
  assign n637 = n578 | n633 ;
  assign n638 = ~n501 & n636 ;
  assign n639 = n602 | n607 ;
  assign n640 = n154 | n276 ;
  assign n641 = n612 | n631 ;
  assign n642 = n224 | n532 ;
  assign n643 = n56 & n57 ;
  assign n644 = n63 & n79 ;
  assign n645 = n59 & n62 ;
  assign n646 = n169 | n182 ;
  assign n647 = n58 & ~n67 ;
  assign n648 = n144 | n212 ;
  assign n649 = n64 & n71 ;
  assign n650 = n52 & n69 ;
  assign n651 = n49 & n62 ;
  assign n652 = n606 & ~n651 ;
  assign n653 = n52 & n55 ;
  assign n654 = n304 | n653 ;
  assign n655 = n49 & n66 ;
  assign n656 = n591 | n655 ;
  assign n657 = n499 | n648 ;
  assign n658 = n60 & n75 ;
  assign n659 = n64 & n78 ;
  assign n660 = ~n67 & n80 ;
  assign n661 = n164 | n490 ;
  assign n662 = n116 | n644 ;
  assign n663 = n652 & ~n662 ;
  assign n664 = n640 | n641 ;
  assign n665 = n219 | n534 ;
  assign n666 = n660 | n661 ;
  assign n667 = n642 | n666 ;
  assign n668 = n439 | n665 ;
  assign n669 = n667 | n668 ;
  assign n670 = n360 | n647 ;
  assign n671 = n105 | n150 ;
  assign n672 = n654 | n671 ;
  assign n673 = n643 | n653 ;
  assign n674 = n664 | n673 ;
  assign n675 = n670 | n674 ;
  assign n676 = n650 | n658 ;
  assign n677 = n94 | n676 ;
  assign n678 = n318 | n639 ;
  assign n679 = n656 | n657 ;
  assign n680 = n646 | n679 ;
  assign n681 = n666 | n678 ;
  assign n682 = n663 & ~n680 ;
  assign n683 = ~n47 & n71 ;
  assign n684 = ~n681 & n682 ;
  assign n685 = n677 | n679 ;
  assign n686 = n537 | n587 ;
  assign n687 = ( ~n649 & n669 ) | ( ~n649 & n683 ) | ( n669 & n683 ) ;
  assign n688 = n649 | n687 ;
  assign n689 = ( n520 & ~n605 ) | ( n520 & n688 ) | ( ~n605 & n688 ) ;
  assign n690 = n685 | n686 ;
  assign n691 = n107 | n530 ;
  assign n692 = n527 | n690 ;
  assign n693 = n46 & n63 ;
  assign n694 = ~n47 & n65 ;
  assign n695 = n605 | n689 ;
  assign n696 = ( n177 & ~n645 ) | ( n177 & n675 ) | ( ~n645 & n675 ) ;
  assign n697 = n645 | n696 ;
  assign n698 = n684 & ~n697 ;
  assign n699 = n659 | n676 ;
  assign n700 = n691 | n699 ;
  assign n701 = n69 & n78 ;
  assign n702 = n63 & ~n67 ;
  assign n703 = ( ~n522 & n643 ) | ( ~n522 & n695 ) | ( n643 & n695 ) ;
  assign n704 = n522 | n703 ;
  assign n705 = ( n148 & ~n702 ) | ( n148 & n704 ) | ( ~n702 & n704 ) ;
  assign n706 = ~n281 & n698 ;
  assign n707 = ( n373 & ~n502 ) | ( n373 & n706 ) | ( ~n502 & n706 ) ;
  assign n708 = ~n373 & n707 ;
  assign n709 = ( n168 & ~n197 ) | ( n168 & n708 ) | ( ~n197 & n708 ) ;
  assign n710 = ~n168 & n709 ;
  assign n711 = ( ~n468 & n701 ) | ( ~n468 & n710 ) | ( n701 & n710 ) ;
  assign n712 = ~n701 & n711 ;
  assign n713 = n64 & ~n67 ;
  assign n714 = n56 & n60 ;
  assign n715 = ~n67 & n69 ;
  assign n716 = n293 | n713 ;
  assign n717 = n59 & n69 ;
  assign n718 = n175 | n716 ;
  assign n719 = n60 & ~n67 ;
  assign n720 = n608 | n719 ;
  assign n721 = n53 & n65 ;
  assign n722 = ( n712 & n717 ) | ( n712 & ~n721 ) | ( n717 & ~n721 ) ;
  assign n723 = n56 & n73 ;
  assign n724 = n714 | n723 ;
  assign n725 = n221 | n246 ;
  assign n726 = n279 | n720 ;
  assign n727 = n651 | n714 ;
  assign n728 = ~n717 & n722 ;
  assign n729 = n296 | n715 ;
  assign n730 = n434 | n729 ;
  assign n731 = n46 & n69 ;
  assign n732 = n286 | n607 ;
  assign n733 = n86 | n182 ;
  assign n734 = n422 | n476 ;
  assign n735 = n52 & n57 ;
  assign n736 = n148 | n735 ;
  assign n737 = n727 | n734 ;
  assign n738 = n726 | n736 ;
  assign n739 = n111 | n713 ;
  assign n740 = n314 | n739 ;
  assign n741 = n738 | n740 ;
  assign n742 = n503 | n659 ;
  assign n743 = ( n231 & ~n580 ) | ( n231 & n741 ) | ( ~n580 & n741 ) ;
  assign n744 = n45 & ~n67 ;
  assign n745 = n286 | n723 ;
  assign n746 = n214 | n727 ;
  assign n747 = n62 & n75 ;
  assign n748 = n650 | n747 ;
  assign n749 = n742 | n748 ;
  assign n750 = n220 | n731 ;
  assign n751 = n153 | n747 ;
  assign n752 = n750 | n751 ;
  assign n753 = n745 | n752 ;
  assign n754 = n52 & n66 ;
  assign n755 = n598 & ~n754 ;
  assign n756 = n53 & n78 ;
  assign n757 = n72 & n78 ;
  assign n758 = n295 | n757 ;
  assign n759 = n55 & n78 ;
  assign n760 = ( n692 & ~n724 ) | ( n692 & n758 ) | ( ~n724 & n758 ) ;
  assign n761 = n724 | n760 ;
  assign n762 = ( n246 & ~n313 ) | ( n246 & n761 ) | ( ~n313 & n761 ) ;
  assign n763 = n718 | n725 ;
  assign n764 = n313 | n762 ;
  assign n765 = n522 | n744 ;
  assign n766 = n724 | n765 ;
  assign n767 = ( ~n420 & n713 ) | ( ~n420 & n764 ) | ( n713 & n764 ) ;
  assign n768 = n420 | n767 ;
  assign n769 = n733 | n766 ;
  assign n770 = n552 | n732 ;
  assign n771 = n732 | n737 ;
  assign n772 = n763 | n771 ;
  assign n773 = ( ~n372 & n434 ) | ( ~n372 & n772 ) | ( n434 & n772 ) ;
  assign n774 = n89 | n232 ;
  assign n775 = n473 | n737 ;
  assign n776 = n730 | n774 ;
  assign n777 = n580 | n743 ;
  assign n778 = n51 & n66 ;
  assign n779 = n52 & n53 ;
  assign n780 = ( n753 & ~n757 ) | ( n753 & n778 ) | ( ~n757 & n778 ) ;
  assign n781 = ( ~n187 & n719 ) | ( ~n187 & n768 ) | ( n719 & n768 ) ;
  assign n782 = n757 | n780 ;
  assign n783 = n372 | n773 ;
  assign n784 = n694 | n782 ;
  assign n785 = n187 | n781 ;
  assign n786 = n56 & n66 ;
  assign n787 = n231 | n783 ;
  assign n788 = n52 & n64 ;
  assign n789 = n647 | n788 ;
  assign n790 = n46 & n57 ;
  assign n791 = n235 | n790 ;
  assign n792 = n461 | n582 ;
  assign n793 = n789 | n791 ;
  assign n794 = n95 | n97 ;
  assign n795 = n173 | n794 ;
  assign n796 = n96 | n631 ;
  assign n797 = n145 | n754 ;
  assign n798 = n90 | n520 ;
  assign n799 = n154 | n717 ;
  assign n800 = n443 | n798 ;
  assign n801 = n791 | n796 ;
  assign n802 = n795 | n797 ;
  assign n803 = n792 | n799 ;
  assign n804 = n564 | n801 ;
  assign n805 = n793 | n803 ;
  assign n806 = n96 | n362 ;
  assign n807 = n759 | n798 ;
  assign n808 = n187 | n601 ;
  assign n809 = n800 | n802 ;
  assign n810 = n52 & n60 ;
  assign n811 = ( ~n343 & n425 ) | ( ~n343 & n804 ) | ( n425 & n804 ) ;
  assign n812 = n116 | n300 ;
  assign n813 = n343 | n811 ;
  assign n814 = n807 | n812 ;
  assign n815 = n806 | n808 ;
  assign n816 = n183 | n557 ;
  assign n817 = n814 | n816 ;
  assign n818 = ( n448 & ~n788 ) | ( n448 & n817 ) | ( ~n788 & n817 ) ;
  assign n819 = n788 | n818 ;
  assign n820 = ( n111 & ~n468 ) | ( n111 & n809 ) | ( ~n468 & n809 ) ;
  assign n821 = ( ~n372 & n694 ) | ( ~n372 & n819 ) | ( n694 & n819 ) ;
  assign n822 = n468 | n820 ;
  assign n823 = n46 & n55 ;
  assign n824 = n372 | n821 ;
  assign n825 = n46 & n60 ;
  assign n826 = n377 | n823 ;
  assign n827 = n59 & n60 ;
  assign n828 = n595 | n827 ;
  assign n829 = n71 & n80 ;
  assign n830 = n442 | n829 ;
  assign n831 = n358 | n830 ;
  assign n832 = n55 & n65 ;
  assign n833 = n65 & n69 ;
  assign n834 = n69 & n75 ;
  assign n835 = n779 | n834 ;
  assign n836 = n89 | n833 ;
  assign n837 = n831 | n832 ;
  assign n838 = ~n427 & n583 ;
  assign n839 = n290 | n313 ;
  assign n840 = n749 | n837 ;
  assign n841 = n51 & n69 ;
  assign n842 = n447 | n841 ;
  assign n843 = n296 | n754 ;
  assign n844 = n842 | n843 ;
  assign n845 = n380 | n844 ;
  assign n846 = n55 & n79 ;
  assign n847 = n829 | n846 ;
  assign n848 = n660 | n836 ;
  assign n849 = n59 & n64 ;
  assign n850 = n410 | n849 ;
  assign n851 = n839 | n848 ;
  assign n852 = n220 | n491 ;
  assign n853 = n826 | n851 ;
  assign n854 = n360 | n850 ;
  assign n855 = n831 | n854 ;
  assign n856 = ~n834 & n838 ;
  assign n857 = n212 | n221 ;
  assign n858 = n847 | n857 ;
  assign n859 = n756 | n841 ;
  assign n860 = n855 | n859 ;
  assign n861 = n302 | n502 ;
  assign n862 = n51 & n58 ;
  assign n863 = ( ~n580 & n628 ) | ( ~n580 & n845 ) | ( n628 & n845 ) ;
  assign n864 = n856 & ~n861 ;
  assign n865 = n835 | n852 ;
  assign n866 = n580 | n863 ;
  assign n867 = n169 | n605 ;
  assign n868 = n487 | n867 ;
  assign n869 = n503 | n779 ;
  assign n870 = ~n770 & n864 ;
  assign n871 = n426 | n433 ;
  assign n872 = n64 & n65 ;
  assign n873 = n869 | n871 ;
  assign n874 = n539 | n867 ;
  assign n875 = n858 | n874 ;
  assign n876 = ( n209 & ~n414 ) | ( n209 & n875 ) | ( ~n414 & n875 ) ;
  assign n877 = n414 | n876 ;
  assign n878 = n503 | n649 ;
  assign n879 = n92 | n381 ;
  assign n880 = n520 | n658 ;
  assign n881 = n352 | n607 ;
  assign n882 = n720 | n881 ;
  assign n883 = n98 | n600 ;
  assign n884 = n57 & n71 ;
  assign n885 = n313 | n439 ;
  assign n886 = n231 | n416 ;
  assign n887 = n45 & n79 ;
  assign n888 = n547 | n829 ;
  assign n889 = n302 | n887 ;
  assign n890 = n883 | n886 ;
  assign n891 = n71 & n72 ;
  assign n892 = n842 | n888 ;
  assign n893 = n164 | n655 ;
  assign n894 = n93 | n893 ;
  assign n895 = n846 | n880 ;
  assign n896 = n894 | n895 ;
  assign n897 = n892 | n896 ;
  assign n898 = ( n442 & n510 ) | ( n442 & ~n897 ) | ( n510 & ~n897 ) ;
  assign n899 = n295 | n553 ;
  assign n900 = n73 & n79 ;
  assign n901 = n153 | n891 ;
  assign n902 = n879 | n901 ;
  assign n903 = n885 | n902 ;
  assign n904 = n878 | n888 ;
  assign n905 = n882 | n903 ;
  assign n906 = ( ~n591 & n900 ) | ( ~n591 & n905 ) | ( n900 & n905 ) ;
  assign n907 = n591 | n906 ;
  assign n908 = ( n100 & ~n723 ) | ( n100 & n907 ) | ( ~n723 & n907 ) ;
  assign n909 = n897 | n898 ;
  assign n910 = n341 | n900 ;
  assign n911 = n592 | n884 ;
  assign n912 = n662 | n911 ;
  assign n913 = n662 | n889 ;
  assign n914 = n899 | n913 ;
  assign n915 = n904 | n912 ;
  assign n916 = n101 | n103 ;
  assign n917 = n796 | n910 ;
  assign n918 = n250 | n593 ;
  assign n919 = n602 | n916 ;
  assign n920 = n917 | n919 ;
  assign n921 = n617 | n918 ;
  assign n922 = n920 | n921 ;
  assign n923 = n71 & n73 ;
  assign n924 = ( n410 & n833 ) | ( n410 & ~n909 ) | ( n833 & ~n909 ) ;
  assign n925 = n909 | n924 ;
  assign n926 = n723 | n908 ;
  assign n927 = n168 | n602 ;
  assign n928 = n92 | n255 ;
  assign n929 = n890 | n928 ;
  assign n930 = n362 | n829 ;
  assign n931 = n147 | n279 ;
  assign n932 = n927 | n931 ;
  assign n933 = n930 | n932 ;
  assign n934 = n57 & ~n59 ;
  assign n935 = ( n57 & n925 ) | ( n57 & ~n934 ) | ( n925 & ~n934 ) ;
  assign n936 = ( n57 & n933 ) | ( n57 & ~n934 ) | ( n933 & ~n934 ) ;
  assign n937 = ~n72 & n79 ;
  assign n938 = ( n79 & n922 ) | ( n79 & ~n937 ) | ( n922 & ~n937 ) ;
  assign n939 = n716 | n918 ;
  assign n940 = n929 | n939 ;
  assign n941 = n58 & n79 ;
  assign n942 = n59 & n72 ;
  assign n943 = n62 & n79 ;
  assign n944 = ( n846 & n915 ) | ( n846 & ~n941 ) | ( n915 & ~n941 ) ;
  assign n945 = n62 & n65 ;
  assign n946 = ( n294 & ~n829 ) | ( n294 & n940 ) | ( ~n829 & n940 ) ;
  assign n947 = n829 | n946 ;
  assign n948 = n941 | n944 ;
  assign n949 = n789 | n881 ;
  assign n950 = n583 & ~n926 ;
  assign n951 = ( n122 & ~n644 ) | ( n122 & n947 ) | ( ~n644 & n947 ) ;
  assign n952 = n644 | n951 ;
  assign n953 = n65 & n80 ;
  assign n954 = n235 | n378 ;
  assign n955 = n57 & n75 ;
  assign n956 = n210 | n283 ;
  assign n957 = n90 | n530 ;
  assign n958 = n638 & ~n957 ;
  assign n959 = n672 | n954 ;
  assign n960 = n58 & n75 ;
  assign n961 = n49 & n80 ;
  assign n962 = n209 | n349 ;
  assign n963 = n59 & n80 ;
  assign n964 = n701 | n962 ;
  assign n965 = n45 & n56 ;
  assign n966 = n952 | n963 ;
  assign n967 = n49 & n58 ;
  assign n968 = n891 | n955 ;
  assign n969 = n49 & n57 ;
  assign n970 = n461 | n862 ;
  assign n971 = n958 & ~n959 ;
  assign n972 = n84 | n891 ;
  assign n973 = n45 & n59 ;
  assign n974 = ~n533 & n638 ;
  assign n975 = n833 | n973 ;
  assign n976 = n258 | n975 ;
  assign n977 = n965 | n972 ;
  assign n978 = n348 | n956 ;
  assign n979 = n968 | n978 ;
  assign n980 = n970 | n979 ;
  assign n981 = n336 | n658 ;
  assign n982 = n976 | n981 ;
  assign n983 = ( n219 & ~n849 ) | ( n219 & n980 ) | ( ~n849 & n980 ) ;
  assign n984 = n849 | n983 ;
  assign n985 = n964 | n977 ;
  assign n986 = n971 & ~n985 ;
  assign n987 = n416 | n715 ;
  assign n988 = ( n173 & n986 ) | ( n173 & ~n987 ) | ( n986 & ~n987 ) ;
  assign n989 = ~n173 & n988 ;
  assign n990 = ( n164 & ~n810 ) | ( n164 & n989 ) | ( ~n810 & n989 ) ;
  assign n991 = ~n164 & n990 ;
  assign n992 = ( n148 & ~n841 ) | ( n148 & n991 ) | ( ~n841 & n991 ) ;
  assign n993 = ~n148 & n992 ;
  assign n994 = ( n400 & ~n414 ) | ( n400 & n993 ) | ( ~n414 & n993 ) ;
  assign n995 = ~n400 & n994 ;
  assign n996 = ~n961 & n995 ;
  assign n997 = n187 | n757 ;
  assign n998 = n258 | n294 ;
  assign n999 = n872 | n941 ;
  assign n1000 = n437 | n960 ;
  assign n1001 = n417 | n612 ;
  assign n1002 = n547 | n1001 ;
  assign n1003 = n228 | n790 ;
  assign n1004 = n260 | n999 ;
  assign n1005 = n974 & ~n1004 ;
  assign n1006 = n211 | n318 ;
  assign n1007 = n235 | n306 ;
  assign n1008 = n998 | n1002 ;
  assign n1009 = n225 | n701 ;
  assign n1010 = n146 | n1000 ;
  assign n1011 = n500 | n1003 ;
  assign n1012 = n1009 | n1010 ;
  assign n1013 = n90 | n786 ;
  assign n1014 = n865 | n1008 ;
  assign n1015 = n393 | n1011 ;
  assign n1016 = n1005 & ~n1014 ;
  assign n1017 = ~n815 & n1016 ;
  assign n1018 = n161 | n1006 ;
  assign n1019 = n153 | n721 ;
  assign n1020 = n87 | n694 ;
  assign n1021 = n1000 | n1019 ;
  assign n1022 = n1007 | n1021 ;
  assign n1023 = n1013 | n1022 ;
  assign n1024 = n756 | n961 ;
  assign n1025 = ~n307 & n1017 ;
  assign n1026 = n1020 | n1024 ;
  assign n1027 = n825 | n997 ;
  assign n1028 = n1023 | n1027 ;
  assign n1029 = ( n628 & ~n778 ) | ( n628 & n1028 ) | ( ~n778 & n1028 ) ;
  assign n1030 = n778 | n1029 ;
  assign n1031 = ( ~n414 & n827 ) | ( ~n414 & n1030 ) | ( n827 & n1030 ) ;
  assign n1032 = n414 | n1031 ;
  assign n1033 = n1018 | n1026 ;
  assign n1034 = n1015 | n1033 ;
  assign n1035 = n302 | n645 ;
  assign n1036 = ( ~n553 & n1025 ) | ( ~n553 & n1035 ) | ( n1025 & n1035 ) ;
  assign n1037 = ~n1035 & n1036 ;
  assign n1038 = ( ~n879 & n1019 ) | ( ~n879 & n1037 ) | ( n1019 & n1037 ) ;
  assign n1039 = ~n1019 & n1038 ;
  assign n1040 = ( ~n109 & n290 ) | ( ~n109 & n1039 ) | ( n290 & n1039 ) ;
  assign n1041 = ~n290 & n1040 ;
  assign n1042 = ( n555 & ~n790 ) | ( n555 & n1041 ) | ( ~n790 & n1041 ) ;
  assign n1043 = ~n555 & n1042 ;
  assign n1044 = ~n410 & n1043 ;
  assign n1045 = n300 | n786 ;
  assign n1046 = n107 | n177 ;
  assign n1047 = n116 | n829 ;
  assign n1048 = n448 | n715 ;
  assign n1049 = n183 | n1045 ;
  assign n1050 = n289 | n862 ;
  assign n1051 = n89 | n659 ;
  assign n1052 = n427 | n846 ;
  assign n1053 = n282 | n1051 ;
  assign n1054 = n150 | n1050 ;
  assign n1055 = n310 | n1048 ;
  assign n1056 = n245 | n961 ;
  assign n1057 = n410 | n1056 ;
  assign n1058 = n1046 | n1057 ;
  assign n1059 = n510 | n900 ;
  assign n1060 = n1049 | n1053 ;
  assign n1061 = n357 | n1059 ;
  assign n1062 = n1055 | n1061 ;
  assign n1063 = ( ~n357 & n589 ) | ( ~n357 & n1060 ) | ( n589 & n1060 ) ;
  assign n1064 = n624 | n1058 ;
  assign n1065 = n1062 | n1064 ;
  assign n1066 = n1047 | n1054 ;
  assign n1067 = n744 | n1052 ;
  assign n1068 = n1063 | n1065 ;
  assign n1069 = n660 | n1067 ;
  assign n1070 = n1066 | n1069 ;
  assign n1071 = n357 | n1063 ;
  assign n1072 = n846 | n965 ;
  assign n1073 = n295 | n502 ;
  assign n1074 = n1072 | n1073 ;
  assign n1075 = ( ~n87 & n1068 ) | ( ~n87 & n1070 ) | ( n1068 & n1070 ) ;
  assign n1076 = n87 | n1070 ;
  assign n1077 = n87 | n1075 ;
  assign n1078 = ( ~n553 & n998 ) | ( ~n553 & n1077 ) | ( n998 & n1077 ) ;
  assign n1079 = n553 | n1078 ;
  assign n1080 = ( n348 & ~n643 ) | ( n348 & n1079 ) | ( ~n643 & n1079 ) ;
  assign n1081 = n643 | n1080 ;
  assign n1082 = ( n271 & ~n400 ) | ( n271 & n1081 ) | ( ~n400 & n1081 ) ;
  assign n1083 = n400 | n1082 ;
  assign n1084 = n1056 | n1074 ;
  assign n1085 = n873 | n1084 ;
  assign n1086 = n209 | n644 ;
  assign n1087 = n101 | n1051 ;
  assign n1088 = n224 | n923 ;
  assign n1089 = n650 | n731 ;
  assign n1090 = n1087 | n1088 ;
  assign n1091 = n552 | n714 ;
  assign n1092 = n843 | n998 ;
  assign n1093 = n336 | n1048 ;
  assign n1094 = n1086 | n1093 ;
  assign n1095 = n827 | n862 ;
  assign n1096 = ( n1034 & ~n1089 ) | ( n1034 & n1094 ) | ( ~n1089 & n1094 ) ;
  assign n1097 = n260 | n1091 ;
  assign n1098 = n278 | n1095 ;
  assign n1099 = n1090 | n1098 ;
  assign n1100 = n1097 | n1099 ;
  assign n1101 = ( n95 & ~n318 ) | ( n95 & n1100 ) | ( ~n318 & n1100 ) ;
  assign n1102 = n318 | n1101 ;
  assign n1103 = ( n295 & ~n592 ) | ( n295 & n1102 ) | ( ~n592 & n1102 ) ;
  assign n1104 = n592 | n1103 ;
  assign n1105 = ( n116 & ~n534 ) | ( n116 & n1104 ) | ( ~n534 & n1104 ) ;
  assign n1106 = n534 | n1105 ;
  assign n1107 = n172 | n1051 ;
  assign n1108 = n714 | n1056 ;
  assign n1109 = n286 | n788 ;
  assign n1110 = n371 | n426 ;
  assign n1111 = n133 | n221 ;
  assign n1112 = n1108 | n1109 ;
  assign n1113 = ( n139 & ~n721 ) | ( n139 & n1112 ) | ( ~n721 & n1112 ) ;
  assign n1114 = n1107 | n1110 ;
  assign n1115 = ( n247 & ~n650 ) | ( n247 & n1106 ) | ( ~n650 & n1106 ) ;
  assign n1116 = n223 | n1048 ;
  assign n1117 = n232 | n426 ;
  assign n1118 = n1111 | n1117 ;
  assign n1119 = n1089 | n1096 ;
  assign n1120 = n1092 | n1114 ;
  assign n1121 = n473 | n1045 ;
  assign n1122 = n1118 | n1121 ;
  assign n1123 = n650 | n1115 ;
  assign n1124 = n1116 | n1122 ;
  assign n1125 = n410 | n827 ;
  assign n1126 = ( n1111 & n1119 ) | ( n1111 & ~n1125 ) | ( n1119 & ~n1125 ) ;
  assign n1127 = n1125 | n1126 ;
  assign n1128 = ( n805 & ~n966 ) | ( n805 & n1124 ) | ( ~n966 & n1124 ) ;
  assign n1129 = ( n719 & ~n747 ) | ( n719 & n1127 ) | ( ~n747 & n1127 ) ;
  assign n1130 = n747 | n1129 ;
  assign n1131 = ( n90 & ~n360 ) | ( n90 & n1130 ) | ( ~n360 & n1130 ) ;
  assign n1132 = n360 | n1131 ;
  assign n1133 = n966 | n1128 ;
  assign n1134 = n489 | n1132 ;
  assign n1135 = n655 | n744 ;
  assign n1136 = n427 | n973 ;
  assign n1137 = n605 | n1136 ;
  assign n1138 = n332 | n941 ;
  assign n1139 = n823 | n825 ;
  assign n1140 = n1137 | n1139 ;
  assign n1141 = n87 | n180 ;
  assign n1142 = n494 | n1138 ;
  assign n1143 = n665 | n1135 ;
  assign n1144 = n342 | n887 ;
  assign n1145 = n358 | n602 ;
  assign n1146 = n276 | n747 ;
  assign n1147 = n585 | n900 ;
  assign n1148 = n1140 | n1142 ;
  assign n1149 = ( ~n600 & n714 ) | ( ~n600 & n1148 ) | ( n714 & n1148 ) ;
  assign n1150 = n425 | n645 ;
  assign n1151 = n600 | n1149 ;
  assign n1152 = n1143 | n1151 ;
  assign n1153 = n1048 | n1145 ;
  assign n1154 = n1152 | n1153 ;
  assign n1155 = ( n637 & ~n945 ) | ( n637 & n1154 ) | ( ~n945 & n1154 ) ;
  assign n1156 = n128 | n884 ;
  assign n1157 = n945 | n1155 ;
  assign n1158 = ( ~n1144 & n1146 ) | ( ~n1144 & n1157 ) | ( n1146 & n1157 ) ;
  assign n1159 = n287 | n833 ;
  assign n1160 = n1144 | n1158 ;
  assign n1161 = ( ~n97 & n879 ) | ( ~n97 & n1160 ) | ( n879 & n1160 ) ;
  assign n1162 = n97 | n1161 ;
  assign n1163 = ( ~n128 & n144 ) | ( ~n128 & n1162 ) | ( n144 & n1162 ) ;
  assign n1164 = n128 | n1163 ;
  assign n1165 = n832 | n1141 ;
  assign n1166 = n1159 | n1165 ;
  assign n1167 = n624 | n1165 ;
  assign n1168 = n95 | n282 ;
  assign n1169 = n162 | n371 ;
  assign n1170 = ( ~n754 & n1147 ) | ( ~n754 & n1166 ) | ( n1147 & n1166 ) ;
  assign n1171 = n823 | n1169 ;
  assign n1172 = n1168 | n1171 ;
  assign n1173 = n1146 | n1156 ;
  assign n1174 = n637 | n945 ;
  assign n1175 = n1172 | n1173 ;
  assign n1176 = ( n288 & ~n891 ) | ( n288 & n1175 ) | ( ~n891 & n1175 ) ;
  assign n1177 = n891 | n1176 ;
  assign n1178 = ( ~n100 & n701 ) | ( ~n100 & n1177 ) | ( n701 & n1177 ) ;
  assign n1179 = n352 | n862 ;
  assign n1180 = ( ~n177 & n1164 ) | ( ~n177 & n1179 ) | ( n1164 & n1179 ) ;
  assign n1181 = n177 | n1180 ;
  assign n1182 = n100 | n1178 ;
  assign n1183 = n1150 | n1179 ;
  assign n1184 = n381 | n1182 ;
  assign n1185 = n279 | n378 ;
  assign n1186 = n447 | n1159 ;
  assign n1187 = n125 | n643 ;
  assign n1188 = n823 | n1187 ;
  assign n1189 = n444 | n1188 ;
  assign n1190 = n84 | n559 ;
  assign n1191 = n148 | n1190 ;
  assign n1192 = n489 | n872 ;
  assign n1193 = n168 | n357 ;
  assign n1194 = n184 | n955 ;
  assign n1195 = n207 | n318 ;
  assign n1196 = n122 | n522 ;
  assign n1197 = n490 | n1192 ;
  assign n1198 = n918 | n1195 ;
  assign n1199 = n1191 | n1196 ;
  assign n1200 = n1193 | n1199 ;
  assign n1201 = n1189 | n1197 ;
  assign n1202 = n1185 | n1200 ;
  assign n1203 = n1198 | n1201 ;
  assign n1204 = n83 | n649 ;
  assign n1205 = n1186 | n1204 ;
  assign n1206 = n224 | n447 ;
  assign n1207 = n1202 | n1205 ;
  assign n1208 = ( n795 & ~n798 ) | ( n795 & n1207 ) | ( ~n798 & n1207 ) ;
  assign n1209 = n1194 | n1206 ;
  assign n1210 = n846 | n1194 ;
  assign n1211 = n798 | n1208 ;
  assign n1212 = ~n164 & n583 ;
  assign n1213 = n517 | n1199 ;
  assign n1214 = ( n220 & ~n884 ) | ( n220 & n1203 ) | ( ~n884 & n1203 ) ;
  assign n1215 = n884 | n1214 ;
  assign n1216 = ( ~n397 & n786 ) | ( ~n397 & n1215 ) | ( n786 & n1215 ) ;
  assign n1217 = n397 | n1216 ;
  assign n1218 = ~n207 & n1212 ;
  assign n1219 = ~n517 & n1218 ;
  assign n1220 = n165 | n235 ;
  assign n1221 = n1209 | n1220 ;
  assign n1222 = n250 | n719 ;
  assign n1223 = n961 | n1222 ;
  assign n1224 = n577 | n1223 ;
  assign n1225 = n1221 | n1223 ;
  assign n1226 = n274 | n1221 ;
  assign n1227 = ~n987 & n1212 ;
  assign n1228 = ( ~n757 & n1211 ) | ( ~n757 & n1217 ) | ( n1211 & n1217 ) ;
  assign n1229 = ~n1210 & n1219 ;
  assign n1230 = n400 | n602 ;
  assign n1231 = n757 | n1228 ;
  assign n1232 = ( ~n312 & n886 ) | ( ~n312 & n1231 ) | ( n886 & n1231 ) ;
  assign n1233 = n312 | n1232 ;
  assign n1234 = ( ~n414 & n833 ) | ( ~n414 & n1229 ) | ( n833 & n1229 ) ;
  assign n1235 = ~n833 & n1234 ;
  assign n1236 = ( ~n1001 & n1230 ) | ( ~n1001 & n1233 ) | ( n1230 & n1233 ) ;
  assign n1237 = n1001 | n1236 ;
  assign n1238 = ( n165 & ~n228 ) | ( n165 & n1237 ) | ( ~n228 & n1237 ) ;
  assign n1239 = n228 | n1238 ;
  assign n1240 = ( n349 & ~n834 ) | ( n349 & n1239 ) | ( ~n834 & n1239 ) ;
  assign n1241 = n834 | n1240 ;
  assign n1242 = ( n345 & ~n756 ) | ( n345 & n1241 ) | ( ~n756 & n1241 ) ;
  assign n1243 = n756 | n1242 ;
  assign n1244 = n426 | n849 ;
  assign n1245 = n197 | n425 ;
  assign n1246 = n375 | n643 ;
  assign n1247 = n1125 | n1244 ;
  assign n1248 = n313 | n367 ;
  assign n1249 = n701 | n788 ;
  assign n1250 = n501 | n872 ;
  assign n1251 = n86 | n433 ;
  assign n1252 = n1248 | n1250 ;
  assign n1253 = n1245 | n1251 ;
  assign n1254 = n1247 | n1252 ;
  assign n1255 = n1253 | n1254 ;
  assign n1256 = n724 | n1246 ;
  assign n1257 = n583 & ~n786 ;
  assign n1258 = n520 | n693 ;
  assign n1259 = ( ~n212 & n302 ) | ( ~n212 & n1255 ) | ( n302 & n1255 ) ;
  assign n1260 = n212 | n1259 ;
  assign n1261 = ( n448 & ~n605 ) | ( n448 & n1260 ) | ( ~n605 & n1260 ) ;
  assign n1262 = n605 | n1261 ;
  assign n1263 = n1248 | n1258 ;
  assign n1264 = n1257 & ~n1263 ;
  assign n1265 = ( n210 & ~n276 ) | ( n210 & n1262 ) | ( ~n276 & n1262 ) ;
  assign n1266 = n328 | n1256 ;
  assign n1267 = n436 | n1244 ;
  assign n1268 = n1264 & ~n1267 ;
  assign n1269 = n91 | n203 ;
  assign n1270 = n658 | n754 ;
  assign n1271 = ( ~n177 & n206 ) | ( ~n177 & n1268 ) | ( n206 & n1268 ) ;
  assign n1272 = n721 | n953 ;
  assign n1273 = n555 | n973 ;
  assign n1274 = n1269 | n1273 ;
  assign n1275 = n1270 | n1274 ;
  assign n1276 = n276 | n1265 ;
  assign n1277 = ( ~n434 & n945 ) | ( ~n434 & n1276 ) | ( n945 & n1276 ) ;
  assign n1278 = n434 | n1277 ;
  assign n1279 = ( ~n343 & n378 ) | ( ~n343 & n1278 ) | ( n378 & n1278 ) ;
  assign n1280 = n343 | n1272 ;
  assign n1281 = n1266 | n1280 ;
  assign n1282 = n1249 | n1273 ;
  assign n1283 = n1167 | n1281 ;
  assign n1284 = n300 | n497 ;
  assign n1285 = n1282 | n1284 ;
  assign n1286 = n206 | n1249 ;
  assign n1287 = n246 | n943 ;
  assign n1288 = n1273 | n1287 ;
  assign n1289 = n1279 | n1283 ;
  assign n1290 = ( ~n97 & n1275 ) | ( ~n97 & n1289 ) | ( n1275 & n1289 ) ;
  assign n1291 = n97 | n1290 ;
  assign n1292 = ( ~n522 & n591 ) | ( ~n522 & n1291 ) | ( n591 & n1291 ) ;
  assign n1293 = n522 | n1292 ;
  assign n1294 = ( n358 & ~n476 ) | ( n358 & n1293 ) | ( ~n476 & n1293 ) ;
  assign n1295 = n476 | n1294 ;
  assign n1296 = ( n146 & n219 ) | ( n146 & ~n1295 ) | ( n219 & ~n1295 ) ;
  assign n1297 = n1295 | n1296 ;
  assign n1298 = ( n645 & n717 ) | ( n645 & ~n1297 ) | ( n717 & ~n1297 ) ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = n282 | n649 ;
  assign n1301 = n1286 | n1300 ;
  assign n1302 = n927 | n1286 ;
  assign n1303 = n343 | n1279 ;
  assign n1304 = n716 | n927 ;
  assign n1305 = ~n206 & n1271 ;
  assign n1306 = n105 | n271 ;
  assign n1307 = n188 | n601 ;
  assign n1308 = n88 | n378 ;
  assign n1309 = n499 | n1306 ;
  assign n1310 = n289 | n591 ;
  assign n1311 = n90 | n349 ;
  assign n1312 = n84 | n723 ;
  assign n1313 = n1059 | n1312 ;
  assign n1314 = n246 | n653 ;
  assign n1315 = n578 | n608 ;
  assign n1316 = n713 | n1309 ;
  assign n1317 = n1169 | n1315 ;
  assign n1318 = n371 | n660 ;
  assign n1319 = n1308 | n1318 ;
  assign n1320 = n1316 | n1319 ;
  assign n1321 = n1311 | n1314 ;
  assign n1322 = n1301 | n1313 ;
  assign n1323 = n683 | n973 ;
  assign n1324 = n94 | n779 ;
  assign n1325 = n1310 | n1323 ;
  assign n1326 = n425 | n557 ;
  assign n1327 = n1324 | n1325 ;
  assign n1328 = n1321 | n1327 ;
  assign n1329 = n1074 | n1326 ;
  assign n1330 = n203 | n248 ;
  assign n1331 = n276 | n415 ;
  assign n1332 = n1317 | n1329 ;
  assign n1333 = n56 & n58 ;
  assign n1334 = n1302 | n1332 ;
  assign n1335 = n660 | n1330 ;
  assign n1336 = n1321 | n1335 ;
  assign n1337 = n1251 | n1335 ;
  assign n1338 = n162 | n1333 ;
  assign n1339 = n1307 | n1331 ;
  assign n1340 = n56 & ~n58 ;
  assign n1341 = n731 | n1306 ;
  assign n1342 = n1326 | n1339 ;
  assign n1343 = n862 | n1326 ;
  assign n1344 = n1328 | n1342 ;
  assign n1345 = n169 | n214 ;
  assign n1346 = ( n461 & ~n887 ) | ( n461 & n1322 ) | ( ~n887 & n1322 ) ;
  assign n1347 = ( n678 & ~n1320 ) | ( n678 & n1344 ) | ( ~n1320 & n1344 ) ;
  assign n1348 = n1320 | n1347 ;
  assign n1349 = n177 | n628 ;
  assign n1350 = n1338 | n1349 ;
  assign n1351 = n665 | n1320 ;
  assign n1352 = n323 | n1345 ;
  assign n1353 = n1350 | n1352 ;
  assign n1354 = n81 | n107 ;
  assign n1355 = ( ~n536 & n1348 ) | ( ~n536 & n1354 ) | ( n1348 & n1354 ) ;
  assign n1356 = n1336 | n1353 ;
  assign n1357 = n536 | n1355 ;
  assign n1358 = ( ~n221 & n1192 ) | ( ~n221 & n1357 ) | ( n1192 & n1357 ) ;
  assign n1359 = n375 | n1318 ;
  assign n1360 = n221 | n1358 ;
  assign n1361 = n576 | n1359 ;
  assign n1362 = n943 | n1360 ;
  assign n1363 = n199 | n1362 ;
  assign n1364 = n105 | n234 ;
  assign n1365 = n828 | n1364 ;
  assign n1366 = n1225 | n1363 ;
  assign n1367 = n607 | n694 ;
  assign n1368 = n1325 | n1367 ;
  assign n1369 = n998 | n1341 ;
  assign n1370 = n1364 | n1368 ;
  assign n1371 = n887 | n1346 ;
  assign n1372 = ( ~n150 & n1356 ) | ( ~n150 & n1367 ) | ( n1356 & n1367 ) ;
  assign n1373 = n150 | n1372 ;
  assign n1374 = ( n437 & ~n503 ) | ( n437 & n1373 ) | ( ~n503 & n1373 ) ;
  assign n1375 = n503 | n1374 ;
  assign n1376 = ( n497 & ~n612 ) | ( n497 & n1375 ) | ( ~n612 & n1375 ) ;
  assign n1377 = n612 | n1376 ;
  assign n1378 = ( n647 & ~n832 ) | ( n647 & n1377 ) | ( ~n832 & n1377 ) ;
  assign n1379 = n832 | n1378 ;
  assign n1380 = n651 | n778 ;
  assign n1381 = n212 | n810 ;
  assign n1382 = n373 | n693 ;
  assign n1383 = n1381 | n1382 ;
  assign n1384 = n100 | n476 ;
  assign n1385 = n1380 | n1383 ;
  assign n1386 = n84 | n713 ;
  assign n1387 = n788 | n1384 ;
  assign n1388 = n124 | n653 ;
  assign n1389 = n997 | n1385 ;
  assign n1390 = n414 | n694 ;
  assign n1391 = n372 | n605 ;
  assign n1392 = n1003 | n1390 ;
  assign n1393 = n1067 | n1392 ;
  assign n1394 = n1003 | n1391 ;
  assign n1395 = n139 | n177 ;
  assign n1396 = n853 | n1395 ;
  assign n1397 = n258 | n1387 ;
  assign n1398 = n282 | n967 ;
  assign n1399 = n1385 | n1397 ;
  assign n1400 = n209 | n702 ;
  assign n1401 = n323 | n887 ;
  assign n1402 = n1394 | n1401 ;
  assign n1403 = n161 | n592 ;
  assign n1404 = n206 | n425 ;
  assign n1405 = n1386 | n1404 ;
  assign n1406 = n1398 | n1403 ;
  assign n1407 = n147 | n357 ;
  assign n1408 = n1396 | n1406 ;
  assign n1409 = n754 | n756 ;
  assign n1410 = n1400 | n1407 ;
  assign n1411 = n1405 | n1410 ;
  assign n1412 = n1408 | n1411 ;
  assign n1413 = ( n805 & ~n1388 ) | ( n805 & n1412 ) | ( ~n1388 & n1412 ) ;
  assign n1414 = n1388 | n1413 ;
  assign n1415 = n300 | n1409 ;
  assign n1416 = n246 | n823 ;
  assign n1417 = n343 | n503 ;
  assign n1418 = n1393 | n1399 ;
  assign n1419 = n1381 | n1417 ;
  assign n1420 = ( ~n318 & n415 ) | ( ~n318 & n1414 ) | ( n415 & n1414 ) ;
  assign n1421 = ( ~n943 & n1360 ) | ( ~n943 & n1418 ) | ( n1360 & n1418 ) ;
  assign n1422 = n1402 | n1419 ;
  assign n1423 = n1389 | n1405 ;
  assign n1424 = n660 | n1417 ;
  assign n1425 = n532 | n841 ;
  assign n1426 = n1424 | n1425 ;
  assign n1427 = n210 | n358 ;
  assign n1428 = n702 | n1427 ;
  assign n1429 = n1415 | n1428 ;
  assign n1430 = n659 | n778 ;
  assign n1431 = n1416 | n1430 ;
  assign n1432 = n318 | n1420 ;
  assign n1433 = ( ~n397 & n841 ) | ( ~n397 & n1432 ) | ( n841 & n1432 ) ;
  assign n1434 = n1204 | n1397 ;
  assign n1435 = n1247 | n1431 ;
  assign n1436 = n1426 | n1435 ;
  assign n1437 = n1185 | n1390 ;
  assign n1438 = n1429 | n1437 ;
  assign n1439 = ( n145 & n420 ) | ( n145 & ~n1422 ) | ( n420 & ~n1422 ) ;
  assign n1440 = n1422 | n1439 ;
  assign n1441 = ~n580 & n583 ;
  assign n1442 = ~n1440 & n1441 ;
  assign n1443 = n397 | n1433 ;
  assign n1444 = n520 | n628 ;
  assign n1445 = n943 | n1421 ;
  assign n1446 = n600 | n1436 ;
  assign n1447 = n1416 | n1444 ;
  assign n1448 = n522 | n900 ;
  assign n1449 = n150 | n1448 ;
  assign n1450 = n274 | n1449 ;
  assign n1451 = n1032 | n1449 ;
  assign n1452 = ( ~n209 & n559 ) | ( ~n209 & n1438 ) | ( n559 & n1438 ) ;
  assign n1453 = n209 | n1452 ;
  assign n1454 = n468 | n1443 ;
  assign n1455 = ( n146 & ~n400 ) | ( n146 & n1453 ) | ( ~n400 & n1453 ) ;
  assign n1456 = n400 | n1455 ;
  assign n1457 = n719 | n960 ;
  assign n1458 = n165 | n234 ;
  assign n1459 = n759 | n1457 ;
  assign n1460 = n286 | n923 ;
  assign n1461 = n222 | n600 ;
  assign n1462 = n1460 | n1461 ;
  assign n1463 = n84 | n592 ;
  assign n1464 = n211 | n715 ;
  assign n1465 = n1459 | n1464 ;
  assign n1466 = n86 | n220 ;
  assign n1467 = n332 | n757 ;
  assign n1468 = n293 | n1467 ;
  assign n1469 = n1463 | n1468 ;
  assign n1470 = n1462 | n1469 ;
  assign n1471 = n1458 | n1465 ;
  assign n1472 = n172 | n303 ;
  assign n1473 = ( ~n197 & n348 ) | ( ~n197 & n1470 ) | ( n348 & n1470 ) ;
  assign n1474 = n1185 | n1466 ;
  assign n1475 = n1472 | n1474 ;
  assign n1476 = n351 | n448 ;
  assign n1477 = n1457 | n1476 ;
  assign n1478 = n197 | n1473 ;
  assign n1479 = n1170 | n1461 ;
  assign n1480 = n755 & ~n1479 ;
  assign n1481 = n550 | n1478 ;
  assign n1482 = n1471 | n1481 ;
  assign n1483 = n467 | n1409 ;
  assign n1484 = n1482 | n1483 ;
  assign n1485 = n717 | n834 ;
  assign n1486 = ( ~n1095 & n1484 ) | ( ~n1095 & n1485 ) | ( n1484 & n1485 ) ;
  assign n1487 = n1095 | n1486 ;
  assign n1488 = ( ~n288 & n341 ) | ( ~n288 & n1487 ) | ( n341 & n1487 ) ;
  assign n1489 = n288 | n1488 ;
  assign n1490 = ( n235 & ~n702 ) | ( n235 & n1489 ) | ( ~n702 & n1489 ) ;
  assign n1491 = n702 | n1490 ;
  assign n1492 = n467 | n1145 ;
  assign n1493 = ( n177 & ~n945 ) | ( n177 & n1491 ) | ( ~n945 & n1491 ) ;
  assign n1494 = n945 | n1493 ;
  assign n1495 = ( ~n580 & n953 ) | ( ~n580 & n1494 ) | ( n953 & n1494 ) ;
  assign n1496 = n580 | n1495 ;
  assign n1497 = n534 | n644 ;
  assign n1498 = n175 | n660 ;
  assign n1499 = n887 | n1388 ;
  assign n1500 = n91 | n101 ;
  assign n1501 = n116 | n279 ;
  assign n1502 = n510 | n534 ;
  assign n1503 = n1500 | n1502 ;
  assign n1504 = n1498 | n1499 ;
  assign n1505 = n162 | n1497 ;
  assign n1506 = n1501 | n1505 ;
  assign n1507 = n867 | n1475 ;
  assign n1508 = n295 | n825 ;
  assign n1509 = n220 | n923 ;
  assign n1510 = n984 | n1508 ;
  assign n1511 = n1507 | n1510 ;
  assign n1512 = n651 | n655 ;
  assign n1513 = n1251 | n1512 ;
  assign n1514 = n146 | n945 ;
  assign n1515 = n1461 | n1514 ;
  assign n1516 = n984 | n1509 ;
  assign n1517 = n1513 | n1516 ;
  assign n1518 = n1451 | n1517 ;
  assign n1519 = n1503 | n1515 ;
  assign n1520 = n960 | n963 ;
  assign n1521 = n1504 | n1519 ;
  assign n1522 = n1511 | n1521 ;
  assign n1523 = ( n886 & ~n1417 ) | ( n886 & n1522 ) | ( ~n1417 & n1522 ) ;
  assign n1524 = n923 | n965 ;
  assign n1525 = n1417 | n1523 ;
  assign n1526 = n81 | n1524 ;
  assign n1527 = n823 | n1526 ;
  assign n1528 = n1506 | n1527 ;
  assign n1529 = n304 | n723 ;
  assign n1530 = ( ~n1520 & n1525 ) | ( ~n1520 & n1529 ) | ( n1525 & n1529 ) ;
  assign n1531 = n1520 | n1530 ;
  assign n1532 = ( n289 & ~n302 ) | ( n289 & n1531 ) | ( ~n302 & n1531 ) ;
  assign n1533 = n302 | n1532 ;
  assign n1534 = ( n417 & ~n823 ) | ( n417 & n1533 ) | ( ~n823 & n1533 ) ;
  assign n1535 = n823 | n1534 ;
  assign n1536 = ( ~n759 & n779 ) | ( ~n759 & n1535 ) | ( n779 & n1535 ) ;
  assign n1537 = n759 | n1536 ;
  assign n1538 = n400 | n1537 ;
  assign n1539 = n1526 | n1538 ;
  assign n1540 = n1423 | n1539 ;
  assign n1541 = ( n866 & n1134 ) | ( n866 & ~n1540 ) | ( n1134 & ~n1540 ) ;
  assign n1542 = n1540 | n1541 ;
  assign n1543 = ( n188 & n367 ) | ( n188 & ~n1528 ) | ( n367 & ~n1528 ) ;
  assign n1544 = n1528 | n1543 ;
  assign n1545 = n410 | n532 ;
  assign n1546 = n124 | n963 ;
  assign n1547 = n234 | n1546 ;
  assign n1548 = n589 | n1192 ;
  assign n1549 = n287 | n713 ;
  assign n1550 = n417 | n1549 ;
  assign n1551 = n550 | n1548 ;
  assign n1552 = n146 | n723 ;
  assign n1553 = n83 | n476 ;
  assign n1554 = n302 | n884 ;
  assign n1555 = n296 | n1554 ;
  assign n1556 = n148 | n534 ;
  assign n1557 = n258 | n1552 ;
  assign n1558 = n89 | n304 ;
  assign n1559 = n246 | n969 ;
  assign n1560 = n1547 | n1553 ;
  assign n1561 = n1345 | n1485 ;
  assign n1562 = n776 | n1561 ;
  assign n1563 = n1560 | n1562 ;
  assign n1564 = n167 | n534 ;
  assign n1565 = n1545 | n1564 ;
  assign n1566 = n1343 | n1565 ;
  assign n1567 = n221 | n643 ;
  assign n1568 = ( n283 & ~n887 ) | ( n283 & n1563 ) | ( ~n887 & n1563 ) ;
  assign n1569 = n1550 | n1556 ;
  assign n1570 = n258 | n1559 ;
  assign n1571 = n1564 | n1570 ;
  assign n1572 = n949 | n1571 ;
  assign n1573 = ( n169 & ~n747 ) | ( n169 & n1572 ) | ( ~n747 & n1572 ) ;
  assign n1574 = n747 | n1573 ;
  assign n1575 = n433 | n1567 ;
  assign n1576 = n128 | n1575 ;
  assign n1577 = n102 | n987 ;
  assign n1578 = n510 | n1558 ;
  assign n1579 = n887 | n1568 ;
  assign n1580 = n649 | n1559 ;
  assign n1581 = n502 | n1580 ;
  assign n1582 = n1576 | n1581 ;
  assign n1583 = ( n530 & ~n645 ) | ( n530 & n1582 ) | ( ~n645 & n1582 ) ;
  assign n1584 = n645 | n1583 ;
  assign n1585 = n234 | n358 ;
  assign n1586 = n1578 | n1585 ;
  assign n1587 = n883 | n1559 ;
  assign n1588 = n1557 | n1569 ;
  assign n1589 = ( ~n343 & n357 ) | ( ~n343 & n1588 ) | ( n357 & n1588 ) ;
  assign n1590 = n343 | n1589 ;
  assign n1591 = n444 | n1590 ;
  assign n1592 = ( n367 & ~n442 ) | ( n367 & n1579 ) | ( ~n442 & n1579 ) ;
  assign n1593 = n442 | n1592 ;
  assign n1594 = n775 | n1551 ;
  assign n1595 = n214 | n716 ;
  assign n1596 = n834 | n1554 ;
  assign n1597 = n1553 | n1596 ;
  assign n1598 = n144 | n1577 ;
  assign n1599 = n1595 | n1597 ;
  assign n1600 = n437 | n973 ;
  assign n1601 = n1598 | n1600 ;
  assign n1602 = n1409 | n1575 ;
  assign n1603 = n813 | n1601 ;
  assign n1604 = n1324 | n1409 ;
  assign n1605 = ( ~n872 & n945 ) | ( ~n872 & n1599 ) | ( n945 & n1599 ) ;
  assign n1606 = n1550 | n1602 ;
  assign n1607 = n967 | n1349 ;
  assign n1608 = n580 | n1607 ;
  assign n1609 = n1601 | n1608 ;
  assign n1610 = n1594 | n1609 ;
  assign n1611 = ( n275 & n1586 ) | ( n275 & ~n1610 ) | ( n1586 & ~n1610 ) ;
  assign n1612 = n1610 | n1611 ;
  assign n1613 = ( n1144 & ~n1381 ) | ( n1144 & n1612 ) | ( ~n1381 & n1612 ) ;
  assign n1614 = n1381 | n1613 ;
  assign n1615 = ( n293 & ~n693 ) | ( n293 & n1614 ) | ( ~n693 & n1614 ) ;
  assign n1616 = n693 | n1615 ;
  assign n1617 = ( n124 & ~n631 ) | ( n124 & n1616 ) | ( ~n631 & n1616 ) ;
  assign n1618 = n631 | n1617 ;
  assign n1619 = ( ~n206 & n245 ) | ( ~n206 & n1618 ) | ( n245 & n1618 ) ;
  assign n1620 = n872 | n1605 ;
  assign n1621 = n206 | n1619 ;
  assign n1622 = n92 | n188 ;
  assign n1623 = n245 | n721 ;
  assign n1624 = n850 | n1622 ;
  assign n1625 = n468 | n631 ;
  assign n1626 = n693 | n1555 ;
  assign n1627 = n97 | n1626 ;
  assign n1628 = n303 | n747 ;
  assign n1629 = n82 | n490 ;
  assign n1630 = n397 | n942 ;
  assign n1631 = n1577 | n1627 ;
  assign n1632 = n281 | n1555 ;
  assign n1633 = n258 | n1630 ;
  assign n1634 = n1625 | n1633 ;
  assign n1635 = n943 | n1629 ;
  assign n1636 = n1628 | n1635 ;
  assign n1637 = n437 | n1636 ;
  assign n1638 = n367 | n1637 ;
  assign n1639 = n1624 | n1638 ;
  assign n1640 = n1631 | n1639 ;
  assign n1641 = ( ~n424 & n565 ) | ( ~n424 & n1640 ) | ( n565 & n1640 ) ;
  assign n1642 = n1395 | n1638 ;
  assign n1643 = n424 | n1641 ;
  assign n1644 = n270 | n1623 ;
  assign n1645 = ( n1230 & ~n1584 ) | ( n1230 & n1643 ) | ( ~n1584 & n1643 ) ;
  assign n1646 = n1634 | n1644 ;
  assign n1647 = n1351 | n1646 ;
  assign n1648 = n352 | n1485 ;
  assign n1649 = n1584 | n1645 ;
  assign n1650 = n295 | n1584 ;
  assign n1651 = ( n306 & ~n1520 ) | ( n306 & n1649 ) | ( ~n1520 & n1649 ) ;
  assign n1652 = n1520 | n1651 ;
  assign n1653 = ( ~n532 & n1648 ) | ( ~n532 & n1652 ) | ( n1648 & n1652 ) ;
  assign n1654 = n532 | n1653 ;
  assign n1655 = ( n147 & ~n891 ) | ( n147 & n1654 ) | ( ~n891 & n1654 ) ;
  assign n1656 = n891 | n1655 ;
  assign n1657 = ( ~n489 & n955 ) | ( ~n489 & n1656 ) | ( n955 & n1656 ) ;
  assign n1658 = n489 | n1657 ;
  assign n1659 = ( ~n107 & n1647 ) | ( ~n107 & n1658 ) | ( n1647 & n1658 ) ;
  assign n1660 = n107 | n1658 ;
  assign n1661 = n279 | n1648 ;
  assign n1662 = n107 | n1659 ;
  assign n1663 = n164 | n279 ;
  assign n1664 = n154 | n735 ;
  assign n1665 = n418 | n1664 ;
  assign n1666 = n304 | n497 ;
  assign n1667 = n1663 | n1666 ;
  assign n1668 = n313 | n348 ;
  assign n1669 = n1665 | n1668 ;
  assign n1670 = n1667 | n1669 ;
  assign n1671 = ( ~n846 & n1333 ) | ( ~n846 & n1670 ) | ( n1333 & n1670 ) ;
  assign n1672 = n996 & ~n1458 ;
  assign n1673 = n846 | n1671 ;
  assign n1674 = ( n351 & ~n591 ) | ( n351 & n1673 ) | ( ~n591 & n1673 ) ;
  assign n1675 = n591 | n1674 ;
  assign n1676 = n90 | n341 ;
  assign n1677 = n713 | n1123 ;
  assign n1678 = n643 | n834 ;
  assign n1679 = n281 | n288 ;
  assign n1680 = n602 | n1679 ;
  assign n1681 = n1678 | n1680 ;
  assign n1682 = n93 | n658 ;
  assign n1683 = n1681 | n1682 ;
  assign n1684 = n357 | n683 ;
  assign n1685 = n1677 | n1684 ;
  assign n1686 = n426 | n1675 ;
  assign n1687 = n719 | n1683 ;
  assign n1688 = n1676 | n1686 ;
  assign n1689 = n996 & ~n1685 ;
  assign n1690 = n880 | n1685 ;
  assign n1691 = n1688 | n1690 ;
  assign n1692 = n125 | n1679 ;
  assign n1693 = n585 | n1692 ;
  assign n1694 = n392 | n1693 ;
  assign n1695 = n936 | n1693 ;
  assign n1696 = n1691 | n1694 ;
  assign n1697 = n810 | n829 ;
  assign n1698 = ( n634 & ~n1660 ) | ( n634 & n1696 ) | ( ~n1660 & n1696 ) ;
  assign n1699 = n1660 | n1698 ;
  assign n1700 = ( n1144 & ~n1388 ) | ( n1144 & n1699 ) | ( ~n1388 & n1699 ) ;
  assign n1701 = n149 | n655 ;
  assign n1702 = n1388 | n1700 ;
  assign n1703 = n997 | n1701 ;
  assign n1704 = n1458 | n1697 ;
  assign n1705 = ( n1136 & ~n1349 ) | ( n1136 & n1702 ) | ( ~n1349 & n1702 ) ;
  assign n1706 = n1349 | n1705 ;
  assign n1707 = n1703 | n1704 ;
  assign n1708 = ( ~n173 & n1159 ) | ( ~n173 & n1706 ) | ( n1159 & n1706 ) ;
  assign n1709 = n592 | n702 ;
  assign n1710 = n634 | n1709 ;
  assign n1711 = n1337 | n1710 ;
  assign n1712 = n206 | n779 ;
  assign n1713 = n810 | n1712 ;
  assign n1714 = n415 | n1630 ;
  assign n1715 = n245 | n655 ;
  assign n1716 = n557 | n645 ;
  assign n1717 = n107 | n1051 ;
  assign n1718 = n605 | n694 ;
  assign n1719 = n336 | n1716 ;
  assign n1720 = n646 | n1184 ;
  assign n1721 = n1713 | n1715 ;
  assign n1722 = n900 | n1717 ;
  assign n1723 = n744 | n884 ;
  assign n1724 = n1714 | n1721 ;
  assign n1725 = n672 | n1687 ;
  assign n1726 = n1720 | n1724 ;
  assign n1727 = n1551 | n1722 ;
  assign n1728 = n228 | n1333 ;
  assign n1729 = n1672 & ~n1719 ;
  assign n1730 = n1192 | n1728 ;
  assign n1731 = n1726 | n1727 ;
  assign n1732 = n165 | n923 ;
  assign n1733 = n1718 | n1732 ;
  assign n1734 = n1723 | n1730 ;
  assign n1735 = n1729 & ~n1734 ;
  assign n1736 = ( ~n312 & n1687 ) | ( ~n312 & n1735 ) | ( n1687 & n1735 ) ;
  assign n1737 = ~n1687 & n1736 ;
  assign n1738 = n373 | n532 ;
  assign n1739 = n1206 | n1712 ;
  assign n1740 = n172 | n367 ;
  assign n1741 = ( n1089 & n1731 ) | ( n1089 & ~n1733 ) | ( n1731 & ~n1733 ) ;
  assign n1742 = n1733 | n1741 ;
  assign n1743 = ( n278 & n1737 ) | ( n278 & ~n1740 ) | ( n1737 & ~n1740 ) ;
  assign n1744 = ~n278 & n1743 ;
  assign n1745 = n210 | n228 ;
  assign n1746 = ( ~n1388 & n1742 ) | ( ~n1388 & n1745 ) | ( n1742 & n1745 ) ;
  assign n1747 = n1388 | n1746 ;
  assign n1748 = ( ~n93 & n1738 ) | ( ~n93 & n1747 ) | ( n1738 & n1747 ) ;
  assign n1749 = n93 | n1748 ;
  assign n1750 = ( ~n522 & n825 ) | ( ~n522 & n1749 ) | ( n825 & n1749 ) ;
  assign n1751 = n522 | n1750 ;
  assign n1752 = ( n175 & ~n862 ) | ( n175 & n1751 ) | ( ~n862 & n1751 ) ;
  assign n1753 = n862 | n1752 ;
  assign n1754 = n833 | n1753 ;
  assign n1755 = n281 | n447 ;
  assign n1756 = n499 | n891 ;
  assign n1757 = n1723 | n1756 ;
  assign n1758 = n232 | n417 ;
  assign n1759 = n1745 | n1758 ;
  assign n1760 = n1755 | n1759 ;
  assign n1761 = n1757 | n1760 ;
  assign n1762 = ( ~n714 & n941 ) | ( ~n714 & n1761 ) | ( n941 & n1761 ) ;
  assign n1763 = n714 | n1762 ;
  assign n1764 = n701 | n833 ;
  assign n1765 = ( n222 & ~n591 ) | ( n222 & n1763 ) | ( ~n591 & n1763 ) ;
  assign n1766 = n109 | n1666 ;
  assign n1767 = n82 | n303 ;
  assign n1768 = n1766 | n1767 ;
  assign n1769 = n139 | n212 ;
  assign n1770 = n397 | n953 ;
  assign n1771 = n1622 | n1769 ;
  assign n1772 = n310 | n1771 ;
  assign n1773 = n591 | n1765 ;
  assign n1774 = n150 | n207 ;
  assign n1775 = n559 | n1774 ;
  assign n1776 = n1519 | n1769 ;
  assign n1777 = n296 | n967 ;
  assign n1778 = n1770 | n1777 ;
  assign n1779 = ( n148 & ~n645 ) | ( n148 & n1773 ) | ( ~n645 & n1773 ) ;
  assign n1780 = n1772 | n1778 ;
  assign n1781 = n645 | n1779 ;
  assign n1782 = n231 | n360 ;
  assign n1783 = n1764 | n1782 ;
  assign n1784 = ( ~n840 & n1032 ) | ( ~n840 & n1780 ) | ( n1032 & n1780 ) ;
  assign n1785 = n1775 | n1783 ;
  assign n1786 = n840 | n1784 ;
  assign n1787 = n1768 | n1785 ;
  assign n1788 = ( n96 & ~n302 ) | ( n96 & n1787 ) | ( ~n302 & n1787 ) ;
  assign n1789 = n302 | n1788 ;
  assign n1790 = ( n248 & ~n461 ) | ( n248 & n1789 ) | ( ~n461 & n1789 ) ;
  assign n1791 = n461 | n1790 ;
  assign n1792 = n849 | n1791 ;
  assign n1793 = ( n840 & ~n1445 ) | ( n840 & n1792 ) | ( ~n1445 & n1792 ) ;
  assign n1794 = n1445 | n1793 ;
  assign n1795 = ( n1496 & ~n1663 ) | ( n1496 & n1794 ) | ( ~n1663 & n1794 ) ;
  assign n1796 = n310 | n1781 ;
  assign n1797 = n1663 | n1795 ;
  assign n1798 = n95 | n212 ;
  assign n1799 = ( n565 & ~n1630 ) | ( n565 & n1797 ) | ( ~n1630 & n1797 ) ;
  assign n1800 = n1391 | n1798 ;
  assign n1801 = n1630 | n1799 ;
  assign n1802 = ( ~n97 & n546 ) | ( ~n97 & n1801 ) | ( n546 & n1801 ) ;
  assign n1803 = n97 | n1802 ;
  assign n1804 = n1796 | n1800 ;
  assign n1805 = n1450 | n1804 ;
  assign n1806 = n559 | n1805 ;
  assign n1807 = n168 | n203 ;
  assign n1808 = n116 | n546 ;
  assign n1809 = n747 | n1136 ;
  assign n1810 = n381 | n643 ;
  assign n1811 = n1354 | n1809 ;
  assign n1812 = n1091 | n1811 ;
  assign n1813 = n1497 | n1811 ;
  assign n1814 = n360 | n1808 ;
  assign n1815 = n1258 | n1810 ;
  assign n1816 = n1807 | n1814 ;
  assign n1817 = n1813 | n1815 ;
  assign n1818 = n105 | n832 ;
  assign n1819 = n86 | n1818 ;
  assign n1820 = n678 | n1819 ;
  assign n1821 = n98 | n644 ;
  assign n1822 = n133 | n373 ;
  assign n1823 = n1820 | n1821 ;
  assign n1824 = n434 | n1822 ;
  assign n1825 = n1812 | n1824 ;
  assign n1826 = n537 | n1820 ;
  assign n1827 = n600 | n1035 ;
  assign n1828 = n1547 | n1823 ;
  assign n1829 = n1770 | n1827 ;
  assign n1830 = n1825 | n1826 ;
  assign n1831 = ( n914 & ~n1777 ) | ( n914 & n1830 ) | ( ~n1777 & n1830 ) ;
  assign n1832 = n1817 | n1829 ;
  assign n1833 = n111 | n442 ;
  assign n1834 = n587 | n1833 ;
  assign n1835 = ( ~n1764 & n1816 ) | ( ~n1764 & n1832 ) | ( n1816 & n1832 ) ;
  assign n1836 = n1707 | n1834 ;
  assign n1837 = n884 | n969 ;
  assign n1838 = n880 | n914 ;
  assign n1839 = ( ~n883 & n1309 ) | ( ~n883 & n1836 ) | ( n1309 & n1836 ) ;
  assign n1840 = n883 | n1839 ;
  assign n1841 = n1764 | n1835 ;
  assign n1842 = n413 | n1841 ;
  assign n1843 = ( ~n539 & n1709 ) | ( ~n539 & n1842 ) | ( n1709 & n1842 ) ;
  assign n1844 = n1777 | n1831 ;
  assign n1845 = n539 | n1843 ;
  assign n1846 = n378 | n461 ;
  assign n1847 = ( ~n1056 & n1837 ) | ( ~n1056 & n1845 ) | ( n1837 & n1845 ) ;
  assign n1848 = n1056 | n1847 ;
  assign n1849 = ( n183 & ~n612 ) | ( n183 & n1848 ) | ( ~n612 & n1848 ) ;
  assign n1850 = n612 | n1849 ;
  assign n1851 = ( n175 & ~n694 ) | ( n175 & n1850 ) | ( ~n694 & n1850 ) ;
  assign n1852 = n694 | n1851 ;
  assign n1853 = n608 | n1852 ;
  assign n1854 = n357 | n1019 ;
  assign n1855 = n169 | n306 ;
  assign n1856 = n94 | n501 ;
  assign n1857 = n548 | n1856 ;
  assign n1858 = n960 | n1514 ;
  assign n1859 = n91 | n591 ;
  assign n1860 = n589 | n941 ;
  assign n1861 = n1858 | n1859 ;
  assign n1862 = n414 | n1854 ;
  assign n1863 = n1857 | n1861 ;
  assign n1864 = n1447 | n1862 ;
  assign n1865 = n1863 | n1864 ;
  assign n1866 = ( ~n957 & n1745 ) | ( ~n957 & n1865 ) | ( n1745 & n1865 ) ;
  assign n1867 = n957 | n1866 ;
  assign n1868 = ( ~n1840 & n1855 ) | ( ~n1840 & n1860 ) | ( n1855 & n1860 ) ;
  assign n1869 = ( n81 & ~n891 ) | ( n81 & n1867 ) | ( ~n891 & n1867 ) ;
  assign n1870 = n1840 | n1868 ;
  assign n1871 = n891 | n1869 ;
  assign n1872 = ( n715 & ~n841 ) | ( n715 & n1871 ) | ( ~n841 & n1871 ) ;
  assign n1873 = n841 | n1872 ;
  assign n1874 = ( n381 & ~n651 ) | ( n381 & n1873 ) | ( ~n651 & n1873 ) ;
  assign n1875 = n651 | n1874 ;
  assign n1876 = n1204 | n1875 ;
  assign n1877 = n1606 | n1876 ;
  assign n1878 = ( ~n144 & n884 ) | ( ~n144 & n1870 ) | ( n884 & n1870 ) ;
  assign n1879 = n144 | n1878 ;
  assign n1880 = n961 | n1879 ;
  assign n1881 = ( n1792 & n1877 ) | ( n1792 & ~n1880 ) | ( n1877 & ~n1880 ) ;
  assign n1882 = n161 | n552 ;
  assign n1883 = n84 | n900 ;
  assign n1884 = n501 | n1883 ;
  assign n1885 = n444 | n1045 ;
  assign n1886 = n1882 | n1884 ;
  assign n1887 = n824 | n1827 ;
  assign n1888 = n1508 | n1827 ;
  assign n1889 = n1885 | n1886 ;
  assign n1890 = ( n579 & ~n1662 ) | ( n579 & n1889 ) | ( ~n1662 & n1889 ) ;
  assign n1891 = n1662 | n1890 ;
  assign n1892 = n91 | n92 ;
  assign n1893 = n700 | n1892 ;
  assign n1894 = n1880 | n1881 ;
  assign n1895 = n1770 | n1846 ;
  assign n1896 = n1893 | n1895 ;
  assign n1897 = n824 | n1862 ;
  assign n1898 = ( n246 & ~n294 ) | ( n246 & n1896 ) | ( ~n294 & n1896 ) ;
  assign n1899 = n207 | n683 ;
  assign n1900 = n294 | n1898 ;
  assign n1901 = n807 | n1860 ;
  assign n1902 = n444 | n967 ;
  assign n1903 = n351 | n700 ;
  assign n1904 = ( ~n522 & n943 ) | ( ~n522 & n1900 ) | ( n943 & n1900 ) ;
  assign n1905 = n522 | n1904 ;
  assign n1906 = n1553 | n1902 ;
  assign n1907 = n1899 | n1906 ;
  assign n1908 = ( n1089 & ~n1733 ) | ( n1089 & n1891 ) | ( ~n1733 & n1891 ) ;
  assign n1909 = n1733 | n1908 ;
  assign n1910 = n476 | n647 ;
  assign n1911 = n502 | n592 ;
  assign n1912 = n209 | n719 ;
  assign n1913 = n107 | n1902 ;
  assign n1914 = n283 | n945 ;
  assign n1915 = n303 | n1914 ;
  assign n1916 = n1910 | n1913 ;
  assign n1917 = n1915 | n1916 ;
  assign n1918 = n683 | n827 ;
  assign n1919 = n602 | n713 ;
  assign n1920 = n102 | n497 ;
  assign n1921 = n1912 | n1919 ;
  assign n1922 = n271 | n735 ;
  assign n1923 = n105 | n342 ;
  assign n1924 = n360 | n832 ;
  assign n1925 = n83 | n555 ;
  assign n1926 = n1921 | n1924 ;
  assign n1927 = n1922 | n1925 ;
  assign n1928 = n1913 | n1923 ;
  assign n1929 = n1912 | n1920 ;
  assign n1930 = n849 | n884 ;
  assign n1931 = n880 | n1911 ;
  assign n1932 = n1195 | n1930 ;
  assign n1933 = n282 | n501 ;
  assign n1934 = n1918 | n1933 ;
  assign n1935 = n343 | n1035 ;
  assign n1936 = n1929 | n1934 ;
  assign n1937 = n600 | n1272 ;
  assign n1938 = n1315 | n1937 ;
  assign n1939 = n1928 | n1932 ;
  assign n1940 = n627 | n1938 ;
  assign n1941 = n1917 | n1940 ;
  assign n1942 = ( ~n102 & n124 ) | ( ~n102 & n1941 ) | ( n124 & n1941 ) ;
  assign n1943 = n102 | n1942 ;
  assign n1944 = n1927 | n1935 ;
  assign n1945 = n83 | n164 ;
  assign n1946 = ( n592 & n941 ) | ( n592 & ~n1939 ) | ( n941 & ~n1939 ) ;
  assign n1947 = n1939 | n1946 ;
  assign n1948 = n1725 | n1944 ;
  assign n1949 = ( n433 & n591 ) | ( n433 & ~n1947 ) | ( n591 & ~n1947 ) ;
  assign n1950 = n1947 | n1949 ;
  assign n1951 = n1091 | n1911 ;
  assign n1952 = n1604 | n1951 ;
  assign n1953 = ( ~n188 & n778 ) | ( ~n188 & n1943 ) | ( n778 & n1943 ) ;
  assign n1954 = ( n468 & n862 ) | ( n468 & ~n1950 ) | ( n862 & ~n1950 ) ;
  assign n1955 = n1950 | n1954 ;
  assign n1956 = n188 | n1953 ;
  assign n1957 = n306 | n943 ;
  assign n1958 = n372 | n1956 ;
  assign n1959 = n721 | n1957 ;
  assign n1960 = n1447 | n1958 ;
  assign n1961 = n1948 | n1960 ;
  assign n1962 = n147 | n833 ;
  assign n1963 = n183 | n1945 ;
  assign n1964 = n210 | n1962 ;
  assign n1965 = n1334 | n1920 ;
  assign n1966 = n1888 | n1964 ;
  assign n1967 = n1931 | n1963 ;
  assign n1968 = n1504 | n1922 ;
  assign n1969 = n1936 | n1963 ;
  assign n1970 = n1936 | n1959 ;
  assign n1971 = n1966 | n1970 ;
  assign n1972 = ( n231 & n963 ) | ( n231 & ~n1955 ) | ( n963 & ~n1955 ) ;
  assign n1973 = n1955 | n1972 ;
  assign n1974 = n627 | n1256 ;
  assign n1975 = n225 | n522 ;
  assign n1976 = ( ~n224 & n1971 ) | ( ~n224 & n1975 ) | ( n1971 & n1975 ) ;
  assign n1977 = n224 | n1976 ;
  assign n1978 = ( ~n713 & n1123 ) | ( ~n713 & n1961 ) | ( n1123 & n1961 ) ;
  assign n1979 = ( ~n304 & n490 ) | ( ~n304 & n1977 ) | ( n490 & n1977 ) ;
  assign n1980 = n304 | n1979 ;
  assign n1981 = ( ~n503 & n887 ) | ( ~n503 & n1980 ) | ( n887 & n1980 ) ;
  assign n1982 = n503 | n1981 ;
  assign n1983 = n713 | n1978 ;
  assign n1984 = ( n139 & ~n965 ) | ( n139 & n1982 ) | ( ~n965 & n1982 ) ;
  assign n1985 = n965 | n1984 ;
  assign n1986 = n271 | n1985 ;
  assign n1987 = n283 | n448 ;
  assign n1988 = ~n92 & n583 ;
  assign n1989 = ~n832 & n1988 ;
  assign n1990 = ~n225 & n1989 ;
  assign n1991 = ~n1856 & n1990 ;
  assign n1992 = n172 | n717 ;
  assign n1993 = ~n1987 & n1991 ;
  assign n1994 = n97 | n133 ;
  assign n1995 = ~n1349 & n1993 ;
  assign n1996 = n336 | n1663 ;
  assign n1997 = n300 | n631 ;
  assign n1998 = n1994 | n1996 ;
  assign n1999 = n197 | n1997 ;
  assign n2000 = ~n1930 & n1993 ;
  assign n2001 = n173 | n286 ;
  assign n2002 = n1992 | n2001 ;
  assign n2003 = n1998 | n2002 ;
  assign n2004 = ( ~n503 & n591 ) | ( ~n503 & n2003 ) | ( n591 & n2003 ) ;
  assign n2005 = n503 | n2004 ;
  assign n2006 = ( n778 & ~n965 ) | ( n778 & n2005 ) | ( ~n965 & n2005 ) ;
  assign n2007 = n147 | n683 ;
  assign n2008 = n1999 | n2007 ;
  assign n2009 = n965 | n2006 ;
  assign n2010 = n758 | n1191 ;
  assign n2011 = n553 | n2007 ;
  assign n2012 = n1995 & ~n2010 ;
  assign n2013 = n2008 | n2009 ;
  assign n2014 = n2012 & ~n2013 ;
  assign n2015 = ( ~n86 & n553 ) | ( ~n86 & n2014 ) | ( n553 & n2014 ) ;
  assign n2016 = ~n553 & n2015 ;
  assign n2017 = ( ~n221 & n224 ) | ( ~n221 & n2016 ) | ( n224 & n2016 ) ;
  assign n2018 = ~n224 & n2017 ;
  assign n2019 = ( ~n723 & n754 ) | ( ~n723 & n2018 ) | ( n754 & n2018 ) ;
  assign n2020 = ~n754 & n2019 ;
  assign n2021 = ( ~n468 & n497 ) | ( ~n468 & n2020 ) | ( n497 & n2020 ) ;
  assign n2022 = ~n497 & n2021 ;
  assign n2023 = n1044 & ~n1091 ;
  assign n2024 = ~n967 & n2022 ;
  assign n2025 = ~n1091 & n2024 ;
  assign n2026 = ~n1944 & n2025 ;
  assign n2027 = ~n1776 & n2026 ;
  assign n2028 = n415 | n593 ;
  assign n2029 = n271 | n313 ;
  assign n2030 = n362 | n433 ;
  assign n2031 = n552 | n943 ;
  assign n2032 = n1338 | n2029 ;
  assign n2033 = n546 | n2028 ;
  assign n2034 = n2031 | n2033 ;
  assign n2035 = n93 | n1664 ;
  assign n2036 = n224 | n502 ;
  assign n2037 = n2035 | n2036 ;
  assign n2038 = ~n217 & n728 ;
  assign n2039 = n1509 | n1591 ;
  assign n2040 = n2038 & ~n2039 ;
  assign n2041 = n234 | n969 ;
  assign n2042 = n375 | n612 ;
  assign n2043 = n434 | n653 ;
  assign n2044 = n2029 | n2042 ;
  assign n2045 = n1650 | n2044 ;
  assign n2046 = n1191 | n2042 ;
  assign n2047 = n936 | n2046 ;
  assign n2048 = n833 | n1664 ;
  assign n2049 = n1739 | n2042 ;
  assign n2050 = n2030 | n2032 ;
  assign n2051 = n2034 | n2050 ;
  assign n2052 = n1907 | n2051 ;
  assign n2053 = n276 | n2052 ;
  assign n2054 = ( ~n1542 & n1975 ) | ( ~n1542 & n2053 ) | ( n1975 & n2053 ) ;
  assign n2055 = n1542 | n2054 ;
  assign n2056 = n884 | n955 ;
  assign n2057 = n2041 | n2056 ;
  assign n2058 = n2009 | n2057 ;
  assign n2059 = ( n93 & ~n105 ) | ( n93 & n2055 ) | ( ~n105 & n2055 ) ;
  assign n2060 = n2034 | n2037 ;
  assign n2061 = n868 | n2057 ;
  assign n2062 = n580 | n999 ;
  assign n2063 = n2060 | n2062 ;
  assign n2064 = n728 & ~n1739 ;
  assign n2065 = n887 | n891 ;
  assign n2066 = n728 & ~n2065 ;
  assign n2067 = n1502 | n2065 ;
  assign n2068 = n2043 | n2065 ;
  assign n2069 = n2023 & ~n2068 ;
  assign n2070 = ~n2058 & n2069 ;
  assign n2071 = n105 | n2059 ;
  assign n2072 = n716 | n1910 ;
  assign n2073 = n555 | n957 ;
  assign n2074 = n1369 | n2073 ;
  assign n2075 = n2072 | n2074 ;
  assign n2076 = ( ~n381 & n967 ) | ( ~n381 & n2075 ) | ( n967 & n2075 ) ;
  assign n2077 = n381 | n2076 ;
  assign n2078 = n287 | n601 ;
  assign n2079 = n313 | n862 ;
  assign n2080 = n735 | n2078 ;
  assign n2081 = n422 | n534 ;
  assign n2082 = n125 | n250 ;
  assign n2083 = n592 | n943 ;
  assign n2084 = n341 | n2082 ;
  assign n2085 = n2083 | n2084 ;
  assign n2086 = n182 | n211 ;
  assign n2087 = n1529 | n2086 ;
  assign n2088 = n2081 | n2087 ;
  assign n2089 = n2078 | n2079 ;
  assign n2090 = n286 | n1382 ;
  assign n2091 = n229 | n281 ;
  assign n2092 = n2089 | n2091 ;
  assign n2093 = n2088 | n2092 ;
  assign n2094 = ( n248 & ~n963 ) | ( n248 & n2093 ) | ( ~n963 & n2093 ) ;
  assign n2095 = n248 | n499 ;
  assign n2096 = n332 | n2095 ;
  assign n2097 = n2085 | n2096 ;
  assign n2098 = n168 | n442 ;
  assign n2099 = ( n111 & ~n400 ) | ( n111 & n2097 ) | ( ~n400 & n2097 ) ;
  assign n2100 = n400 | n2099 ;
  assign n2101 = n963 | n2094 ;
  assign n2102 = n81 | n2098 ;
  assign n2103 = ( n1754 & n2027 ) | ( n1754 & ~n2100 ) | ( n2027 & ~n2100 ) ;
  assign n2104 = ~n1754 & n2103 ;
  assign n2105 = ~n2102 & n2104 ;
  assign n2106 = n96 | n731 ;
  assign n2107 = ~n2091 & n2105 ;
  assign n2108 = n744 | n759 ;
  assign n2109 = n746 | n2106 ;
  assign n2110 = n2090 | n2108 ;
  assign n2111 = n2089 | n2109 ;
  assign n2112 = n1697 | n2100 ;
  assign n2113 = n1189 | n2109 ;
  assign n2114 = n2101 | n2110 ;
  assign n2115 = n2047 | n2114 ;
  assign n2116 = ( ~n82 & n645 ) | ( ~n82 & n2115 ) | ( n645 & n2115 ) ;
  assign n2117 = n82 | n2116 ;
  assign n2118 = n187 | n900 ;
  assign n2119 = n343 | n2117 ;
  assign n2120 = n694 | n2118 ;
  assign n2121 = n1861 | n2119 ;
  assign n2122 = n2063 | n2121 ;
  assign n2123 = n2110 | n2120 ;
  assign n2124 = n1967 | n2123 ;
  assign n2125 = n124 | n348 ;
  assign n2126 = n295 | n923 ;
  assign n2127 = n276 | n778 ;
  assign n2128 = n184 | n427 ;
  assign n2129 = n281 | n360 ;
  assign n2130 = n582 | n2127 ;
  assign n2131 = n721 | n2125 ;
  assign n2132 = n501 | n778 ;
  assign n2133 = n2126 | n2132 ;
  assign n2134 = n2131 | n2133 ;
  assign n2135 = n1058 | n2130 ;
  assign n2136 = n2128 | n2129 ;
  assign n2137 = n664 | n2125 ;
  assign n2138 = n1243 | n2136 ;
  assign n2139 = n228 | n717 ;
  assign n2140 = n2135 | n2138 ;
  assign n2141 = n206 | n246 ;
  assign n2142 = n1564 | n2132 ;
  assign n2143 = n1118 | n2132 ;
  assign n2144 = n2082 | n2139 ;
  assign n2145 = n754 | n2141 ;
  assign n2146 = n1113 | n2136 ;
  assign n2147 = n2134 | n2146 ;
  assign n2148 = n351 | n415 ;
  assign n2149 = ( ~n757 & n1217 ) | ( ~n757 & n2147 ) | ( n1217 & n2147 ) ;
  assign n2150 = n1989 & ~n2148 ;
  assign n2151 = n757 | n2149 ;
  assign n2152 = n348 | n489 ;
  assign n2153 = n2037 | n2152 ;
  assign n2154 = n2150 & ~n2153 ;
  assign n2155 = n122 | n1111 ;
  assign n2156 = n2145 | n2155 ;
  assign n2157 = n2144 | n2156 ;
  assign n2158 = n449 | n2145 ;
  assign n2159 = n580 | n1087 ;
  assign n2160 = ( ~n462 & n2124 ) | ( ~n462 & n2157 ) | ( n2124 & n2157 ) ;
  assign n2161 = n462 | n2160 ;
  assign n2162 = n153 | n183 ;
  assign n2163 = n449 | n2162 ;
  assign n2164 = n2159 | n2163 ;
  assign n2165 = n342 | n1333 ;
  assign n2166 = n282 | n2165 ;
  assign n2167 = n1724 | n2166 ;
  assign n2168 = n2126 | n2166 ;
  assign n2169 = n2164 | n2168 ;
  assign n2170 = n86 | n555 ;
  assign n2171 = n217 | n2170 ;
  assign n2172 = n225 | n645 ;
  assign n2173 = n246 | n786 ;
  assign n2174 = n245 | n841 ;
  assign n2175 = n2172 | n2174 ;
  assign n2176 = n341 | n522 ;
  assign n2177 = n372 | n400 ;
  assign n2178 = n149 | n2173 ;
  assign n2179 = n2176 | n2177 ;
  assign n2180 = n2171 | n2178 ;
  assign n2181 = n1181 | n2179 ;
  assign n2182 = n2180 | n2181 ;
  assign n2183 = n177 | n209 ;
  assign n2184 = n582 | n2183 ;
  assign n2185 = n426 | n790 ;
  assign n2186 = n90 | n2185 ;
  assign n2187 = n1775 | n2170 ;
  assign n2188 = n1120 | n1853 ;
  assign n2189 = n2184 | n2188 ;
  assign n2190 = n503 | n1883 ;
  assign n2191 = n1913 | n2177 ;
  assign n2192 = n1120 | n1758 ;
  assign n2193 = n235 | n2186 ;
  assign n2194 = n1883 | n1914 ;
  assign n2195 = n644 | n2190 ;
  assign n2196 = n2193 | n2194 ;
  assign n2197 = ( ~n302 & n647 ) | ( ~n302 & n2182 ) | ( n647 & n2182 ) ;
  assign n2198 = n302 | n2197 ;
  assign n2199 = n2142 | n2196 ;
  assign n2200 = n111 | n2139 ;
  assign n2201 = ( ~n133 & n2128 ) | ( ~n133 & n2199 ) | ( n2128 & n2199 ) ;
  assign n2202 = n2193 | n2200 ;
  assign n2203 = n2175 | n2198 ;
  assign n2204 = n2202 | n2203 ;
  assign n2205 = n250 | n1622 ;
  assign n2206 = n2175 | n2205 ;
  assign n2207 = n1859 | n2183 ;
  assign n2208 = n2206 | n2207 ;
  assign n2209 = ( n502 & ~n649 ) | ( n502 & n2208 ) | ( ~n649 & n2208 ) ;
  assign n2210 = n649 | n2209 ;
  assign n2211 = ( ~n222 & n547 ) | ( ~n222 & n2210 ) | ( n547 & n2210 ) ;
  assign n2212 = n222 | n2211 ;
  assign n2213 = n592 | n834 ;
  assign n2214 = ( ~n427 & n434 ) | ( ~n427 & n2212 ) | ( n434 & n2212 ) ;
  assign n2215 = n133 | n2201 ;
  assign n2216 = ( ~n212 & n461 ) | ( ~n212 & n2215 ) | ( n461 & n2215 ) ;
  assign n2217 = n212 | n2216 ;
  assign n2218 = n427 | n2214 ;
  assign n2219 = n744 | n2183 ;
  assign n2220 = n2213 | n2219 ;
  assign n2221 = n82 | n659 ;
  assign n2222 = n702 | n1333 ;
  assign n2223 = n91 | n645 ;
  assign n2224 = n2221 | n2222 ;
  assign n2225 = n702 | n2223 ;
  assign n2226 = n214 | n1088 ;
  assign n2227 = n93 | n756 ;
  assign n2228 = n2224 | n2226 ;
  assign n2229 = n373 | n833 ;
  assign n2230 = n88 | n955 ;
  assign n2231 = n916 | n2229 ;
  assign n2232 = n173 | n942 ;
  assign n2233 = n211 | n2232 ;
  assign n2234 = n2148 | n2231 ;
  assign n2235 = n536 | n2233 ;
  assign n2236 = ~n148 & n583 ;
  assign n2237 = n2230 | n2235 ;
  assign n2238 = n1578 | n2237 ;
  assign n2239 = n2234 | n2238 ;
  assign n2240 = n650 | n834 ;
  assign n2241 = n94 | n300 ;
  assign n2242 = n2236 & ~n2241 ;
  assign n2243 = n2228 | n2240 ;
  assign n2244 = ~n1022 & n2242 ;
  assign n2245 = ~n2239 & n2244 ;
  assign n2246 = n122 | n490 ;
  assign n2247 = ~n2227 & n2245 ;
  assign n2248 = ~n2246 & n2247 ;
  assign n2249 = ( ~n303 & n1192 ) | ( ~n303 & n2248 ) | ( n1192 & n2248 ) ;
  assign n2250 = ~n1192 & n2249 ;
  assign n2251 = n2195 | n2225 ;
  assign n2252 = ( n105 & ~n884 ) | ( n105 & n2250 ) | ( ~n884 & n2250 ) ;
  assign n2253 = ~n105 & n2252 ;
  assign n2254 = ~n468 & n2253 ;
  assign n2255 = ~n2223 & n2254 ;
  assign n2256 = ~n2243 & n2255 ;
  assign n2257 = n1361 | n1758 ;
  assign n2258 = ~n1969 & n2256 ;
  assign n2259 = n1758 | n2080 ;
  assign n2260 = n888 | n1821 ;
  assign n2261 = n2259 | n2260 ;
  assign n2262 = n982 | n2228 ;
  assign n2263 = n1056 | n2148 ;
  assign n2264 = n544 | n2232 ;
  assign n2265 = ~n1181 & n2258 ;
  assign n2266 = n437 | n823 ;
  assign n2267 = n644 | n2266 ;
  assign n2268 = n1740 | n2267 ;
  assign n2269 = n1361 | n2268 ;
  assign n2270 = n867 | n2268 ;
  assign n2271 = n2262 | n2269 ;
  assign n2272 = n87 | n95 ;
  assign n2273 = n279 | n2272 ;
  assign n2274 = ( n567 & ~n1697 ) | ( n567 & n2265 ) | ( ~n1697 & n2265 ) ;
  assign n2275 = ~n567 & n2274 ;
  assign n2276 = n2254 & ~n2273 ;
  assign n2277 = n83 | n2273 ;
  assign n2278 = ~n2257 & n2276 ;
  assign n2279 = n536 | n1663 ;
  assign n2280 = n2043 | n2240 ;
  assign n2281 = n105 | n790 ;
  assign n2282 = n2279 | n2280 ;
  assign n2283 = n437 | n943 ;
  assign n2284 = n258 | n731 ;
  assign n2285 = n150 | n503 ;
  assign n2286 = n107 | n658 ;
  assign n2287 = n2281 | n2284 ;
  assign n2288 = n241 | n283 ;
  assign n2289 = n2285 | n2286 ;
  assign n2290 = n197 | n303 ;
  assign n2291 = n2284 | n2290 ;
  assign n2292 = n1701 | n2126 ;
  assign n2293 = n2289 | n2292 ;
  assign n2294 = n841 | n1050 ;
  assign n2295 = n2283 | n2288 ;
  assign n2296 = n95 | n490 ;
  assign n2297 = n2291 | n2294 ;
  assign n2298 = n1442 & ~n2240 ;
  assign n2299 = n2178 | n2297 ;
  assign n2300 = n148 | n225 ;
  assign n2301 = n1701 | n2300 ;
  assign n2302 = n2295 | n2301 ;
  assign n2303 = n155 | n2295 ;
  assign n2304 = ~n769 & n2298 ;
  assign n2305 = n155 | n2296 ;
  assign n2306 = n2287 | n2305 ;
  assign n2307 = n1475 | n2287 ;
  assign n2308 = n2261 | n2307 ;
  assign n2309 = n838 & ~n1187 ;
  assign n2310 = ~n2303 & n2309 ;
  assign n2311 = ( ~n1146 & n1338 ) | ( ~n1146 & n2308 ) | ( n1338 & n2308 ) ;
  assign n2312 = n1146 | n2311 ;
  assign n2313 = n87 | n349 ;
  assign n2314 = n89 | n2313 ;
  assign n2315 = n2297 | n2314 ;
  assign n2316 = n1887 | n2314 ;
  assign n2317 = n1382 | n2041 ;
  assign n2318 = n2306 | n2317 ;
  assign n2319 = ( ~n342 & n2266 ) | ( ~n342 & n2318 ) | ( n2266 & n2318 ) ;
  assign n2320 = n342 | n2319 ;
  assign n2321 = ( n607 & ~n825 ) | ( n607 & n2320 ) | ( ~n825 & n2320 ) ;
  assign n2322 = n825 | n2321 ;
  assign n2323 = n94 | n342 ;
  assign n2324 = n161 | n510 ;
  assign n2325 = n293 | n1630 ;
  assign n2326 = n96 | n650 ;
  assign n2327 = n1050 | n1111 ;
  assign n2328 = n843 | n2324 ;
  assign n2329 = n555 | n744 ;
  assign n2330 = n1050 | n2329 ;
  assign n2331 = n2327 | n2328 ;
  assign n2332 = n2323 | n2330 ;
  assign n2333 = n95 | n612 ;
  assign n2334 = n256 | n2185 ;
  assign n2335 = n2332 | n2334 ;
  assign n2336 = n2325 | n2333 ;
  assign n2337 = n141 | n2336 ;
  assign n2338 = n2154 & ~n2337 ;
  assign n2339 = ( ~n1514 & n2312 ) | ( ~n1514 & n2324 ) | ( n2312 & n2324 ) ;
  assign n2340 = n1514 | n2339 ;
  assign n2341 = n2001 | n2326 ;
  assign n2342 = n1552 | n2336 ;
  assign n2343 = n2331 | n2341 ;
  assign n2344 = ( n212 & ~n790 ) | ( n212 & n2343 ) | ( ~n790 & n2343 ) ;
  assign n2345 = n790 | n2344 ;
  assign n2346 = ( n415 & ~n683 ) | ( n415 & n2345 ) | ( ~n683 & n2345 ) ;
  assign n2347 = ~n1144 & n2338 ;
  assign n2348 = ~n97 & n2347 ;
  assign n2349 = n2281 | n2326 ;
  assign n2350 = n2302 | n2349 ;
  assign n2351 = n97 | n234 ;
  assign n2352 = ( ~n649 & n2340 ) | ( ~n649 & n2351 ) | ( n2340 & n2351 ) ;
  assign n2353 = n649 | n2352 ;
  assign n2354 = ( n490 & ~n644 ) | ( n490 & n2348 ) | ( ~n644 & n2348 ) ;
  assign n2355 = ( ~n442 & n497 ) | ( ~n442 & n2335 ) | ( n497 & n2335 ) ;
  assign n2356 = ~n490 & n2354 ;
  assign n2357 = ( ~n372 & n759 ) | ( ~n372 & n2356 ) | ( n759 & n2356 ) ;
  assign n2358 = ~n759 & n2357 ;
  assign n2359 = ( ~n182 & n628 ) | ( ~n182 & n2353 ) | ( n628 & n2353 ) ;
  assign n2360 = n182 | n2359 ;
  assign n2361 = ( n203 & ~n973 ) | ( n203 & n2360 ) | ( ~n973 & n2360 ) ;
  assign n2362 = n683 | n2346 ;
  assign n2363 = n973 | n2361 ;
  assign n2364 = n442 | n2355 ;
  assign n2365 = ( ~n655 & n2161 ) | ( ~n655 & n2363 ) | ( n2161 & n2363 ) ;
  assign n2366 = n434 | n2364 ;
  assign n2367 = ~n444 & n2358 ;
  assign n2368 = n655 | n2365 ;
  assign n2369 = n197 | n2362 ;
  assign n2370 = n93 | n779 ;
  assign n2371 = n2152 | n2370 ;
  assign n2372 = n235 | n290 ;
  assign n2373 = n342 | n589 ;
  assign n2374 = n304 | n1697 ;
  assign n2375 = n1910 | n2372 ;
  assign n2376 = n2371 | n2374 ;
  assign n2377 = n2375 | n2376 ;
  assign n2378 = n162 | n423 ;
  assign n2379 = n2373 | n2378 ;
  assign n2380 = n214 | n1388 ;
  assign n2381 = ( ~n422 & n2377 ) | ( ~n422 & n2380 ) | ( n2377 & n2380 ) ;
  assign n2382 = n759 | n1318 ;
  assign n2383 = n2379 | n2382 ;
  assign n2384 = n776 | n2383 ;
  assign n2385 = n422 | n2381 ;
  assign n2386 = ( ~n649 & n658 ) | ( ~n649 & n2385 ) | ( n658 & n2385 ) ;
  assign n2387 = n649 | n2386 ;
  assign n2388 = ( n721 & ~n841 ) | ( n721 & n2387 ) | ( ~n841 & n2387 ) ;
  assign n2389 = n841 | n2388 ;
  assign n2390 = n82 | n349 ;
  assign n2391 = n2326 | n2390 ;
  assign n2392 = n1853 | n2230 ;
  assign n2393 = n2391 | n2392 ;
  assign n2394 = n2384 | n2393 ;
  assign n2395 = ( ~n678 & n2389 ) | ( ~n678 & n2394 ) | ( n2389 & n2394 ) ;
  assign n2396 = n225 | n2177 ;
  assign n2397 = n843 | n2390 ;
  assign n2398 = n325 | n2397 ;
  assign n2399 = n167 | n945 ;
  assign n2400 = n332 | n2399 ;
  assign n2401 = n2157 | n2400 ;
  assign n2402 = n415 | n2380 ;
  assign n2403 = n1195 | n2402 ;
  assign n2404 = n2401 | n2403 ;
  assign n2405 = n82 | n998 ;
  assign n2406 = ( n501 & ~n827 ) | ( n501 & n2398 ) | ( ~n827 & n2398 ) ;
  assign n2407 = n678 | n2395 ;
  assign n2408 = ( ~n886 & n2024 ) | ( ~n886 & n2407 ) | ( n2024 & n2407 ) ;
  assign n2409 = ~n2407 & n2408 ;
  assign n2410 = n2396 | n2402 ;
  assign n2411 = n1324 | n2405 ;
  assign n2412 = n1608 | n2411 ;
  assign n2413 = n352 | n468 ;
  assign n2414 = n964 | n2413 ;
  assign n2415 = n1324 | n2413 ;
  assign n2416 = n2410 | n2415 ;
  assign n2417 = n2315 | n2416 ;
  assign n2418 = n173 | n547 ;
  assign n2419 = ( ~n293 & n490 ) | ( ~n293 & n2409 ) | ( n490 & n2409 ) ;
  assign n2420 = ~n1138 & n1235 ;
  assign n2421 = n2396 | n2418 ;
  assign n2422 = n2296 | n2396 ;
  assign n2423 = ~n1193 & n1235 ;
  assign n2424 = ~n2422 & n2423 ;
  assign n2425 = n2263 | n2421 ;
  assign n2426 = n103 | n644 ;
  assign n2427 = n81 | n1349 ;
  assign n2428 = n162 | n832 ;
  assign n2429 = n122 | n375 ;
  assign n2430 = n555 | n1136 ;
  assign n2431 = n476 | n2427 ;
  assign n2432 = n343 | n2430 ;
  assign n2433 = n500 | n1623 ;
  assign n2434 = n164 | n303 ;
  assign n2435 = n2426 | n2434 ;
  assign n2436 = n2433 | n2435 ;
  assign n2437 = n476 | n530 ;
  assign n2438 = n602 | n846 ;
  assign n2439 = n2383 | n2431 ;
  assign n2440 = n2043 | n2430 ;
  assign n2441 = n209 | n872 ;
  assign n2442 = n2437 | n2441 ;
  assign n2443 = n2428 | n2435 ;
  assign n2444 = n1930 | n2429 ;
  assign n2445 = n2436 | n2439 ;
  assign n2446 = n187 | n232 ;
  assign n2447 = n2440 | n2442 ;
  assign n2448 = n580 | n2446 ;
  assign n2449 = ( n381 & ~n580 ) | ( n381 & n2445 ) | ( ~n580 & n2445 ) ;
  assign n2450 = n2443 | n2444 ;
  assign n2451 = n645 | n735 ;
  assign n2452 = n2448 | n2451 ;
  assign n2453 = n779 | n1905 ;
  assign n2454 = n580 | n2449 ;
  assign n2455 = n2432 | n2452 ;
  assign n2456 = n188 | n683 ;
  assign n2457 = n247 | n2456 ;
  assign n2458 = n2187 | n2457 ;
  assign n2459 = ( ~n779 & n1905 ) | ( ~n779 & n2454 ) | ( n1905 & n2454 ) ;
  assign n2460 = n779 | n2459 ;
  assign n2461 = n552 | n961 ;
  assign n2462 = n1001 | n2461 ;
  assign n2463 = n2457 | n2462 ;
  assign n2464 = n2450 | n2463 ;
  assign n2465 = n442 | n559 ;
  assign n2466 = n2438 | n2465 ;
  assign n2467 = n281 | n891 ;
  assign n2468 = ( ~n111 & n2198 ) | ( ~n111 & n2464 ) | ( n2198 & n2464 ) ;
  assign n2469 = n534 | n1427 ;
  assign n2470 = n2467 | n2469 ;
  assign n2471 = n100 | n631 ;
  assign n2472 = n578 | n2471 ;
  assign n2473 = n2342 | n2472 ;
  assign n2474 = n2466 | n2472 ;
  assign n2475 = n2470 | n2474 ;
  assign n2476 = n723 | n2475 ;
  assign n2477 = n221 | n345 ;
  assign n2478 = n2152 | n2477 ;
  assign n2479 = n2466 | n2478 ;
  assign n2480 = n111 | n2468 ;
  assign n2481 = n241 | n683 ;
  assign n2482 = n175 | n846 ;
  assign n2483 = n694 | n2482 ;
  assign n2484 = n2139 | n2483 ;
  assign n2485 = n1088 | n2351 ;
  assign n2486 = n2481 | n2485 ;
  assign n2487 = n187 | n591 ;
  assign n2488 = n87 | n111 ;
  assign n2489 = n841 | n2488 ;
  assign n2490 = n102 | n683 ;
  assign n2491 = n1591 | n2490 ;
  assign n2492 = n2489 | n2491 ;
  assign n2493 = n286 | n693 ;
  assign n2494 = n109 | n2493 ;
  assign n2495 = n276 | n381 ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = n2406 | n2486 ;
  assign n2498 = n419 | n2487 ;
  assign n2499 = n827 | n2406 ;
  assign n2500 = n2484 | n2492 ;
  assign n2501 = n2388 | n2500 ;
  assign n2502 = n219 | n960 ;
  assign n2503 = n1169 | n2502 ;
  assign n2504 = n848 | n2486 ;
  assign n2505 = n827 | n1846 ;
  assign n2506 = n2503 | n2505 ;
  assign n2507 = n546 | n942 ;
  assign n2508 = n923 | n2501 ;
  assign n2509 = n2497 | n2506 ;
  assign n2510 = n2498 | n2507 ;
  assign n2511 = n2479 | n2510 ;
  assign n2512 = n534 | n580 ;
  assign n2513 = n2498 | n2512 ;
  assign n2514 = n1183 | n2513 ;
  assign n2515 = n2504 | n2514 ;
  assign n2516 = n910 | n2493 ;
  assign n2517 = n1365 | n2516 ;
  assign n2518 = ( n1275 & ~n2496 ) | ( n1275 & n2511 ) | ( ~n2496 & n2511 ) ;
  assign n2519 = n2496 | n2518 ;
  assign n2520 = ( ~n1345 & n1860 ) | ( ~n1345 & n2519 ) | ( n1860 & n2519 ) ;
  assign n2521 = n1466 | n1856 ;
  assign n2522 = n714 | n2493 ;
  assign n2523 = n1345 | n2520 ;
  assign n2524 = ( ~n246 & n300 ) | ( ~n246 & n2523 ) | ( n300 & n2523 ) ;
  assign n2525 = n246 | n2524 ;
  assign n2526 = ( n96 & ~n207 ) | ( n96 & n2525 ) | ( ~n207 & n2525 ) ;
  assign n2527 = n207 | n2526 ;
  assign n2528 = ( ~n241 & n279 ) | ( ~n241 & n2527 ) | ( n279 & n2527 ) ;
  assign n2529 = n241 | n2528 ;
  assign n2530 = n2521 | n2522 ;
  assign n2531 = n428 | n1312 ;
  assign n2532 = n2483 | n2531 ;
  assign n2533 = n418 | n2529 ;
  assign n2534 = n2281 | n2529 ;
  assign n2535 = n219 | n248 ;
  assign n2536 = n116 | n849 ;
  assign n2537 = n731 | n2536 ;
  assign n2538 = n307 | n2162 ;
  assign n2539 = n552 | n655 ;
  assign n2540 = n2535 | n2537 ;
  assign n2541 = n164 | n825 ;
  assign n2542 = n415 | n647 ;
  assign n2543 = n2539 | n2542 ;
  assign n2544 = n877 | n1756 ;
  assign n2545 = n2538 | n2544 ;
  assign n2546 = n2540 | n2545 ;
  assign n2547 = ( ~n2324 & n2541 ) | ( ~n2324 & n2546 ) | ( n2541 & n2546 ) ;
  assign n2548 = n2324 | n2547 ;
  assign n2549 = n362 | n589 ;
  assign n2550 = ( ~n98 & n2548 ) | ( ~n98 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2551 = n282 | n502 ;
  assign n2552 = n631 | n2551 ;
  assign n2553 = n98 | n2550 ;
  assign n2554 = ( ~n93 & n304 ) | ( ~n93 & n2553 ) | ( n304 & n2553 ) ;
  assign n2555 = n93 | n2554 ;
  assign n2556 = n2543 | n2552 ;
  assign n2557 = n1968 | n2556 ;
  assign n2558 = ( ~n591 & n1333 ) | ( ~n591 & n2555 ) | ( n1333 & n2555 ) ;
  assign n2559 = n591 | n2558 ;
  assign n2560 = ( n167 & ~n442 ) | ( n167 & n2559 ) | ( ~n442 & n2559 ) ;
  assign n2561 = ( n501 & ~n650 ) | ( n501 & n2557 ) | ( ~n650 & n2557 ) ;
  assign n2562 = n442 | n2560 ;
  assign n2563 = n650 | n2561 ;
  assign n2564 = n973 | n2562 ;
  assign n2565 = n381 | n2563 ;
  assign n2566 = ( ~n2140 & n2564 ) | ( ~n2140 & n2565 ) | ( n2564 & n2565 ) ;
  assign n2567 = n2140 | n2566 ;
  assign n2568 = ( n716 & ~n1035 ) | ( n716 & n2567 ) | ( ~n1035 & n2567 ) ;
  assign n2569 = n1035 | n2568 ;
  assign n2570 = n1770 | n2502 ;
  assign n2571 = n2488 | n2502 ;
  assign n2572 = n2543 | n2570 ;
  assign n2573 = n96 | n1529 ;
  assign n2574 = n2571 | n2573 ;
  assign n2575 = n349 | n702 ;
  assign n2576 = n2502 | n2575 ;
  assign n2577 = n2532 | n2576 ;
  assign n2578 = ( ~n1144 & n1338 ) | ( ~n1144 & n2577 ) | ( n1338 & n2577 ) ;
  assign n2579 = n1144 | n2578 ;
  assign n2580 = ( ~n998 & n2541 ) | ( ~n998 & n2579 ) | ( n2541 & n2579 ) ;
  assign n2581 = n998 | n2580 ;
  assign n2582 = ( ~n289 & n2185 ) | ( ~n289 & n2581 ) | ( n2185 & n2581 ) ;
  assign n2583 = n289 | n2582 ;
  assign n2584 = ( n415 & ~n754 ) | ( n415 & n2583 ) | ( ~n754 & n2583 ) ;
  assign n2585 = n754 | n2584 ;
  assign n2586 = ( ~n358 & n578 ) | ( ~n358 & n2585 ) | ( n578 & n2585 ) ;
  assign n2587 = n358 | n2586 ;
  assign n2588 = ( ~n580 & n601 ) | ( ~n580 & n2587 ) | ( n601 & n2587 ) ;
  assign n2589 = n580 | n2588 ;
  assign n2590 = n173 | n1111 ;
  assign n2591 = n91 | n883 ;
  assign n2592 = n150 | n336 ;
  assign n2593 = n180 | n1679 ;
  assign n2594 = n101 | n228 ;
  assign n2595 = n1630 | n2591 ;
  assign n2596 = n1390 | n2595 ;
  assign n2597 = n2590 | n2592 ;
  assign n2598 = n2230 | n2593 ;
  assign n2599 = n468 | n884 ;
  assign n2600 = n258 | n2594 ;
  assign n2601 = n1926 | n2600 ;
  assign n2602 = n2304 & ~n2596 ;
  assign n2603 = n109 | n647 ;
  assign n2604 = n2458 | n2601 ;
  assign n2605 = n286 | n2603 ;
  assign n2606 = n2592 | n2599 ;
  assign n2607 = n100 | n900 ;
  assign n2608 = n2605 | n2607 ;
  assign n2609 = n284 | n2575 ;
  assign n2610 = n2608 | n2609 ;
  assign n2611 = n153 | n400 ;
  assign n2612 = n2412 | n2598 ;
  assign n2613 = n128 | n461 ;
  assign n2614 = ( n2602 & ~n2611 ) | ( n2602 & n2613 ) | ( ~n2611 & n2613 ) ;
  assign n2615 = ~n2613 & n2614 ;
  assign n2616 = ( n82 & ~n84 ) | ( n82 & n2615 ) | ( ~n84 & n2615 ) ;
  assign n2617 = n884 | n900 ;
  assign n2618 = ~n82 & n2616 ;
  assign n2619 = ( n281 & ~n437 ) | ( n281 & n2618 ) | ( ~n437 & n2618 ) ;
  assign n2620 = ~n281 & n2619 ;
  assign n2621 = ( ~n144 & n891 ) | ( ~n144 & n2620 ) | ( n891 & n2620 ) ;
  assign n2622 = ~n891 & n2621 ;
  assign n2623 = ( n197 & ~n232 ) | ( n197 & n2622 ) | ( ~n232 & n2622 ) ;
  assign n2624 = ~n197 & n2623 ;
  assign n2625 = ( ~n102 & n360 ) | ( ~n102 & n2624 ) | ( n360 & n2624 ) ;
  assign n2626 = ~n360 & n2625 ;
  assign n2627 = ~n651 & n2626 ;
  assign n2628 = ( ~n559 & n2610 ) | ( ~n559 & n2612 ) | ( n2610 & n2612 ) ;
  assign n2629 = n1538 | n2610 ;
  assign n2630 = n559 | n2628 ;
  assign n2631 = ( n1258 & ~n2597 ) | ( n1258 & n2630 ) | ( ~n2597 & n2630 ) ;
  assign n2632 = n2597 | n2631 ;
  assign n2633 = ( n1089 & ~n2611 ) | ( n1089 & n2632 ) | ( ~n2611 & n2632 ) ;
  assign n2634 = n2611 | n2633 ;
  assign n2635 = n214 | n608 ;
  assign n2636 = ( ~n683 & n2446 ) | ( ~n683 & n2634 ) | ( n2446 & n2634 ) ;
  assign n2637 = n683 | n2636 ;
  assign n2638 = ( n579 & n2604 ) | ( n579 & ~n2635 ) | ( n2604 & ~n2635 ) ;
  assign n2639 = ( n846 & ~n941 ) | ( n846 & n2637 ) | ( ~n941 & n2637 ) ;
  assign n2640 = n941 | n2639 ;
  assign n2641 = n2635 | n2638 ;
  assign n2642 = ( ~n1417 & n1733 ) | ( ~n1417 & n2641 ) | ( n1733 & n2641 ) ;
  assign n2643 = n1417 | n2642 ;
  assign n2644 = ( ~n93 & n2266 ) | ( ~n93 & n2643 ) | ( n2266 & n2643 ) ;
  assign n2645 = n93 | n2644 ;
  assign n2646 = ( n87 & ~n510 ) | ( n87 & n2645 ) | ( ~n510 & n2645 ) ;
  assign n2647 = n510 | n2646 ;
  assign n2648 = ( n510 & ~n714 ) | ( n510 & n2640 ) | ( ~n714 & n2640 ) ;
  assign n2649 = n714 | n2648 ;
  assign n2650 = n448 | n2649 ;
  assign n2651 = n1769 | n2366 ;
  assign n2652 = n579 | n2333 ;
  assign n2653 = n313 | n683 ;
  assign n2654 = n850 | n1629 ;
  assign n2655 = n371 | n655 ;
  assign n2656 = n175 | n2086 ;
  assign n2657 = n248 | n649 ;
  assign n2658 = n2231 | n2657 ;
  assign n2659 = n2655 | n2656 ;
  assign n2660 = n209 | n778 ;
  assign n2661 = n2654 | n2660 ;
  assign n2662 = n2651 | n2658 ;
  assign n2663 = n332 | n468 ;
  assign n2664 = n832 | n955 ;
  assign n2665 = n381 | n916 ;
  assign n2666 = n2653 | n2661 ;
  assign n2667 = n1552 | n2666 ;
  assign n2668 = n2652 | n2667 ;
  assign n2669 = n497 | n605 ;
  assign n2670 = n197 | n941 ;
  assign n2671 = n2664 | n2665 ;
  assign n2672 = n1183 | n2671 ;
  assign n2673 = n2668 | n2672 ;
  assign n2674 = ( ~n2177 & n2670 ) | ( ~n2177 & n2673 ) | ( n2670 & n2673 ) ;
  assign n2675 = n2177 | n2674 ;
  assign n2676 = n838 & ~n2223 ;
  assign n2677 = ( ~n2663 & n2669 ) | ( ~n2663 & n2675 ) | ( n2669 & n2675 ) ;
  assign n2678 = n2663 | n2677 ;
  assign n2679 = n293 | n448 ;
  assign n2680 = ( ~n133 & n2657 ) | ( ~n133 & n2678 ) | ( n2657 & n2678 ) ;
  assign n2681 = n96 | n941 ;
  assign n2682 = n133 | n2680 ;
  assign n2683 = n1920 | n2681 ;
  assign n2684 = ( ~n162 & n235 ) | ( ~n162 & n2682 ) | ( n235 & n2682 ) ;
  assign n2685 = n1339 | n2659 ;
  assign n2686 = n162 | n2684 ;
  assign n2687 = n2676 & ~n2683 ;
  assign n2688 = n757 | n2686 ;
  assign n2689 = n1621 | n2688 ;
  assign n2690 = n2685 | n2689 ;
  assign n2691 = n1695 | n2690 ;
  assign n2692 = ( n1889 & ~n2453 ) | ( n1889 & n2691 ) | ( ~n2453 & n2691 ) ;
  assign n2693 = n2453 | n2692 ;
  assign n2694 = n184 | n229 ;
  assign n2695 = n221 | n352 ;
  assign n2696 = n2049 | n2694 ;
  assign n2697 = n255 | n295 ;
  assign n2698 = n2679 | n2695 ;
  assign n2699 = ~n2143 & n2687 ;
  assign n2700 = n146 | n468 ;
  assign n2701 = ( ~n306 & n2185 ) | ( ~n306 & n2693 ) | ( n2185 & n2693 ) ;
  assign n2702 = n2697 | n2700 ;
  assign n2703 = n306 | n2701 ;
  assign n2704 = n149 | n232 ;
  assign n2705 = n2696 | n2698 ;
  assign n2706 = n2296 | n2704 ;
  assign n2707 = n2702 | n2706 ;
  assign n2708 = ( ~n963 & n2705 ) | ( ~n963 & n2707 ) | ( n2705 & n2707 ) ;
  assign n2709 = n963 | n2708 ;
  assign n2710 = ( n1738 & n2635 ) | ( n1738 & ~n2709 ) | ( n2635 & ~n2709 ) ;
  assign n2711 = n2709 | n2710 ;
  assign n2712 = n510 | n2704 ;
  assign n2713 = n963 | n2707 ;
  assign n2714 = n313 | n1764 ;
  assign n2715 = ( ~n83 & n285 ) | ( ~n83 & n2711 ) | ( n285 & n2711 ) ;
  assign n2716 = n83 | n2715 ;
  assign n2717 = n950 & ~n1629 ;
  assign n2718 = n911 | n2716 ;
  assign n2719 = n999 | n1709 ;
  assign n2720 = n999 | n1094 ;
  assign n2721 = n2714 | n2719 ;
  assign n2722 = n209 | n2296 ;
  assign n2723 = n838 & ~n1623 ;
  assign n2724 = n658 | n849 ;
  assign n2725 = ~n1815 & n2723 ;
  assign n2726 = n282 | n2724 ;
  assign n2727 = n2600 | n2726 ;
  assign n2728 = n2428 | n2726 ;
  assign n2729 = n1509 | n2428 ;
  assign n2730 = n225 | n891 ;
  assign n2731 = n229 | n1333 ;
  assign n2732 = n2730 | n2731 ;
  assign n2733 = n2727 | n2732 ;
  assign n2734 = n841 | n965 ;
  assign n2735 = n612 | n2734 ;
  assign n2736 = n2251 | n2735 ;
  assign n2737 = n2662 | n2736 ;
  assign n2738 = n1920 | n2162 ;
  assign n2739 = ( n647 & ~n963 ) | ( n647 & n2733 ) | ( ~n963 & n2733 ) ;
  assign n2740 = ~n2496 & n2627 ;
  assign n2741 = n2603 | n2735 ;
  assign n2742 = n978 | n1566 ;
  assign n2743 = n2741 | n2742 ;
  assign n2744 = n187 | n965 ;
  assign n2745 = ( n563 & n608 ) | ( n563 & ~n849 ) | ( n608 & ~n849 ) ;
  assign n2746 = ~n910 & n2242 ;
  assign n2747 = n849 | n2745 ;
  assign n2748 = ( ~n651 & n2699 ) | ( ~n651 & n2747 ) | ( n2699 & n2747 ) ;
  assign n2749 = n418 | n2507 ;
  assign n2750 = n307 | n413 ;
  assign n2751 = n1133 | n1754 ;
  assign n2752 = n2728 | n2738 ;
  assign n2753 = n532 | n790 ;
  assign n2754 = n2370 | n2753 ;
  assign n2755 = n2111 | n2752 ;
  assign n2756 = n2744 | n2754 ;
  assign n2757 = n1769 | n2162 ;
  assign n2758 = n2749 | n2756 ;
  assign n2759 = n456 | n1245 ;
  assign n2760 = n827 | n1973 ;
  assign n2761 = n2746 & ~n2759 ;
  assign n2762 = n168 | n222 ;
  assign n2763 = n2760 | n2762 ;
  assign n2764 = ~n2747 & n2748 ;
  assign n2765 = n2740 & ~n2763 ;
  assign n2766 = n102 | n154 ;
  assign n2767 = ~n1434 & n2765 ;
  assign n2768 = n476 | n2766 ;
  assign n2769 = n2757 | n2768 ;
  assign n2770 = n2120 | n2768 ;
  assign n2771 = n183 | n358 ;
  assign n2772 = n92 | n559 ;
  assign n2773 = n1256 | n1958 ;
  assign n2774 = ( ~n935 & n1410 ) | ( ~n935 & n2767 ) | ( n1410 & n2767 ) ;
  assign n2775 = n2771 | n2772 ;
  assign n2776 = n1138 | n2775 ;
  assign n2777 = n2756 | n2775 ;
  assign n2778 = n2061 | n2777 ;
  assign n2779 = n150 | n211 ;
  assign n2780 = n1821 | n2660 ;
  assign n2781 = n977 | n2779 ;
  assign n2782 = n2780 | n2781 ;
  assign n2783 = n109 | n397 ;
  assign n2784 = ( ~n371 & n502 ) | ( ~n371 & n2782 ) | ( n502 & n2782 ) ;
  assign n2785 = n461 | n2783 ;
  assign n2786 = n371 | n2784 ;
  assign n2787 = n90 | n2786 ;
  assign n2788 = n2785 | n2787 ;
  assign n2789 = n284 | n2785 ;
  assign n2790 = n2721 | n2789 ;
  assign n2791 = n434 | n651 ;
  assign n2792 = n1480 & ~n2788 ;
  assign n2793 = n647 | n786 ;
  assign n2794 = ( ~n92 & n153 ) | ( ~n92 & n2790 ) | ( n153 & n2790 ) ;
  assign n2795 = n139 | n779 ;
  assign n2796 = n294 | n713 ;
  assign n2797 = n2446 | n2796 ;
  assign n2798 = n2793 | n2797 ;
  assign n2799 = n162 | n1477 ;
  assign n2800 = n963 | n2739 ;
  assign n2801 = n827 | n2800 ;
  assign n2802 = n1018 | n2801 ;
  assign n2803 = n92 | n2794 ;
  assign n2804 = ( ~n228 & n503 ) | ( ~n228 & n2803 ) | ( n503 & n2803 ) ;
  assign n2805 = n228 | n2804 ;
  assign n2806 = ( n88 & ~n756 ) | ( n88 & n2798 ) | ( ~n756 & n2798 ) ;
  assign n2807 = n756 | n2806 ;
  assign n2808 = n2462 | n2807 ;
  assign n2809 = n1711 | n2808 ;
  assign n2810 = n1045 | n2220 ;
  assign n2811 = ( ~n1574 & n2350 ) | ( ~n1574 & n2810 ) | ( n2350 & n2810 ) ;
  assign n2812 = n81 | n144 ;
  assign n2813 = n2795 | n2812 ;
  assign n2814 = n2787 | n2813 ;
  assign n2815 = n2799 | n2814 ;
  assign n2816 = n148 | n650 ;
  assign n2817 = n2137 | n2815 ;
  assign n2818 = n150 | n499 ;
  assign n2819 = n2816 | n2818 ;
  assign n2820 = n2791 | n2819 ;
  assign n2821 = n165 | n247 ;
  assign n2822 = n2813 | n2821 ;
  assign n2823 = n2820 | n2822 ;
  assign n2824 = n123 | n2820 ;
  assign n2825 = n2725 & ~n2824 ;
  assign n2826 = n2534 | n2823 ;
  assign n2827 = ( n853 & ~n1417 ) | ( n853 & n2826 ) | ( ~n1417 & n2826 ) ;
  assign n2828 = ( ~n658 & n945 ) | ( ~n658 & n2805 ) | ( n945 & n2805 ) ;
  assign n2829 = n658 | n2828 ;
  assign n2830 = n961 | n1333 ;
  assign n2831 = n2172 | n2830 ;
  assign n2832 = n288 | n2830 ;
  assign n2833 = n784 | n2041 ;
  assign n2834 = n860 | n2832 ;
  assign n2835 = n2077 | n2832 ;
  assign n2836 = n2414 | n2835 ;
  assign n2837 = n336 | n628 ;
  assign n2838 = n2761 & ~n2834 ;
  assign n2839 = n1930 | n2837 ;
  assign n2840 = n2833 | n2839 ;
  assign n2841 = n810 | n963 ;
  assign n2842 = n2832 | n2841 ;
  assign n2843 = n2840 | n2842 ;
  assign n2844 = ( ~n1384 & n2669 ) | ( ~n1384 & n2843 ) | ( n2669 & n2843 ) ;
  assign n2845 = n1384 | n2844 ;
  assign n2846 = ( ~n302 & n532 ) | ( ~n302 & n2845 ) | ( n532 & n2845 ) ;
  assign n2847 = n188 | n756 ;
  assign n2848 = n302 | n2846 ;
  assign n2849 = ( n221 & ~n923 ) | ( n221 & n2848 ) | ( ~n923 & n2848 ) ;
  assign n2850 = n754 | n1930 ;
  assign n2851 = n1514 | n2847 ;
  assign n2852 = n1938 | n2851 ;
  assign n2853 = n1315 | n2851 ;
  assign n2854 = n2850 | n2853 ;
  assign n2855 = n95 | n289 ;
  assign n2856 = n923 | n2849 ;
  assign n2857 = ( ~n90 & n172 ) | ( ~n90 & n2856 ) | ( n172 & n2856 ) ;
  assign n2858 = n300 | n2855 ;
  assign n2859 = n90 | n2857 ;
  assign n2860 = n2192 | n2858 ;
  assign n2861 = ( ~n589 & n832 ) | ( ~n589 & n2859 ) | ( n832 & n2859 ) ;
  assign n2862 = n589 | n2861 ;
  assign n2863 = n2400 | n2862 ;
  assign n2864 = n2066 & ~n2863 ;
  assign n2865 = n283 | n1230 ;
  assign n2866 = ~n1226 & n2864 ;
  assign n2867 = n721 | n2865 ;
  assign n2868 = n2747 | n2865 ;
  assign n2869 = n2717 & ~n2867 ;
  assign n2870 = n2477 | n2841 ;
  assign n2871 = n1719 | n2870 ;
  assign n2872 = n84 | n306 ;
  assign n2873 = n629 | n2865 ;
  assign n2874 = n2860 | n2873 ;
  assign n2875 = n815 | n1001 ;
  assign n2876 = n2872 | n2875 ;
  assign n2877 = n2000 & ~n2876 ;
  assign n2878 = n2858 | n2876 ;
  assign n2879 = n287 | n530 ;
  assign n2880 = n1454 | n2879 ;
  assign n2881 = n1012 | n2880 ;
  assign n2882 = n2067 | n2881 ;
  assign n2883 = ( n2825 & ~n2862 ) | ( n2825 & n2881 ) | ( ~n2862 & n2881 ) ;
  assign n2884 = ~n2881 & n2883 ;
  assign n2885 = ( ~n561 & n815 ) | ( ~n561 & n2884 ) | ( n815 & n2884 ) ;
  assign n2886 = ~n815 & n2885 ;
  assign n2887 = n293 | n973 ;
  assign n2888 = n468 | n2887 ;
  assign n2889 = n229 | n1272 ;
  assign n2890 = n342 | n846 ;
  assign n2891 = n197 | n833 ;
  assign n2892 = n827 | n2891 ;
  assign n2893 = n356 | n2892 ;
  assign n2894 = n2889 | n2890 ;
  assign n2895 = n2888 | n2892 ;
  assign n2896 = n600 | n694 ;
  assign n2897 = n2893 | n2894 ;
  assign n2898 = n213 | n591 ;
  assign n2899 = n2896 | n2898 ;
  assign n2900 = n1307 | n1381 ;
  assign n2901 = n724 | n2900 ;
  assign n2902 = ( n149 & ~n371 ) | ( n149 & n2897 ) | ( ~n371 & n2897 ) ;
  assign n2903 = n935 | n2901 ;
  assign n2904 = n371 | n2902 ;
  assign n2905 = ( ~n90 & n555 ) | ( ~n90 & n2904 ) | ( n555 & n2904 ) ;
  assign n2906 = n90 | n2905 ;
  assign n2907 = n1824 | n2888 ;
  assign n2908 = n967 | n2906 ;
  assign n2909 = n247 | n352 ;
  assign n2910 = n2899 | n2901 ;
  assign n2911 = n2271 | n2910 ;
  assign n2912 = n1544 | n2909 ;
  assign n2913 = ( ~n2324 & n2874 ) | ( ~n2324 & n2909 ) | ( n2874 & n2909 ) ;
  assign n2914 = n769 | n2908 ;
  assign n2915 = n414 | n724 ;
  assign n2916 = n2912 | n2914 ;
  assign n2917 = n209 | n650 ;
  assign n2918 = n1250 | n1272 ;
  assign n2919 = n1586 | n2917 ;
  assign n2920 = n2324 | n2913 ;
  assign n2921 = n2918 | n2919 ;
  assign n2922 = n124 | n224 ;
  assign n2923 = n150 | n2922 ;
  assign n2924 = n2899 | n2923 ;
  assign n2925 = n2916 | n2924 ;
  assign n2926 = ( n1636 & ~n2446 ) | ( n1636 & n2925 ) | ( ~n2446 & n2925 ) ;
  assign n2927 = n2446 | n2926 ;
  assign n2928 = ( ~n101 & n1860 ) | ( ~n101 & n2927 ) | ( n1860 & n2927 ) ;
  assign n2929 = n499 | n963 ;
  assign n2930 = n101 | n2928 ;
  assign n2931 = ( n786 & ~n788 ) | ( n786 & n2930 ) | ( ~n788 & n2930 ) ;
  assign n2932 = n788 | n2931 ;
  assign n2933 = ( ~n222 & n530 ) | ( ~n222 & n2932 ) | ( n530 & n2932 ) ;
  assign n2934 = n832 | n2929 ;
  assign n2935 = n2050 | n2934 ;
  assign n2936 = n2921 | n2935 ;
  assign n2937 = n222 | n2933 ;
  assign n2938 = n1627 | n2937 ;
  assign n2939 = n735 | n953 ;
  assign n2940 = ( n585 & n2920 ) | ( n585 & ~n2939 ) | ( n2920 & ~n2939 ) ;
  assign n2941 = n2939 | n2940 ;
  assign n2942 = n220 | n658 ;
  assign n2943 = n169 | n2942 ;
  assign n2944 = n1508 | n1911 ;
  assign n2945 = n2943 | n2944 ;
  assign n2946 = n2907 | n2945 ;
  assign n2947 = n122 | n660 ;
  assign n2948 = ( ~n177 & n345 ) | ( ~n177 & n2946 ) | ( n345 & n2946 ) ;
  assign n2949 = n177 | n2948 ;
  assign n2950 = n969 | n2949 ;
  assign n2951 = n2947 | n2950 ;
  assign n2952 = n2080 | n2950 ;
  assign n2953 = n1045 | n2947 ;
  assign n2954 = ( ~n422 & n713 ) | ( ~n422 & n2941 ) | ( n713 & n2941 ) ;
  assign n2955 = n422 | n2954 ;
  assign n2956 = n1689 & ~n2953 ;
  assign n2957 = n744 | n2955 ;
  assign n2958 = n2517 | n2957 ;
  assign n2959 = n2951 | n2958 ;
  assign n2960 = n228 | n1712 ;
  assign n2961 = n2917 | n2960 ;
  assign n2962 = n702 | n2917 ;
  assign n2963 = n202 | n2962 ;
  assign n2964 = n2167 | n2959 ;
  assign n2965 = ( ~n1248 & n1875 ) | ( ~n1248 & n2964 ) | ( n1875 & n2964 ) ;
  assign n2966 = n717 | n719 ;
  assign n2967 = n705 | n1856 ;
  assign n2968 = n2963 | n2967 ;
  assign n2969 = n559 | n2915 ;
  assign n2970 = n2915 | n2966 ;
  assign n2971 = n1856 | n2969 ;
  assign n2972 = n721 | n1975 ;
  assign n2973 = n2132 | n2969 ;
  assign n2974 = n1663 | n2372 ;
  assign n2975 = n961 | n2972 ;
  assign n2976 = n2974 | n2975 ;
  assign n2977 = n2971 | n2976 ;
  assign n2978 = ( n550 & ~n1248 ) | ( n550 & n2977 ) | ( ~n1248 & n2977 ) ;
  assign n2979 = n1248 | n2978 ;
  assign n2980 = ( n557 & ~n1187 ) | ( n557 & n2979 ) | ( ~n1187 & n2979 ) ;
  assign n2981 = n1187 | n2980 ;
  assign n2982 = n954 | n2679 ;
  assign n2983 = n2975 | n2982 ;
  assign n2984 = n1245 | n2086 ;
  assign n2985 = n2983 | n2984 ;
  assign n2986 = ( n2251 & ~n2942 ) | ( n2251 & n2981 ) | ( ~n2942 & n2981 ) ;
  assign n2987 = ( n283 & ~n302 ) | ( n283 & n2985 ) | ( ~n302 & n2985 ) ;
  assign n2988 = n302 | n2987 ;
  assign n2989 = ( ~n778 & n955 ) | ( ~n778 & n2988 ) | ( n955 & n2988 ) ;
  assign n2990 = n2942 | n2986 ;
  assign n2991 = n778 | n2989 ;
  assign n2992 = n447 | n943 ;
  assign n2993 = n520 | n923 ;
  assign n2994 = n154 | n442 ;
  assign n2995 = n2067 | n2992 ;
  assign n2996 = n2011 | n2994 ;
  assign n2997 = n546 | n585 ;
  assign n2998 = n2993 | n2995 ;
  assign n2999 = n500 | n2997 ;
  assign n3000 = n1477 | n2996 ;
  assign n3001 = n2999 | n3000 ;
  assign n3002 = n1477 | n1666 ;
  assign n3003 = n423 | n461 ;
  assign n3004 = n2679 | n3003 ;
  assign n3005 = n2952 | n3001 ;
  assign n3006 = n2048 | n3004 ;
  assign n3007 = n205 | n2997 ;
  assign n3008 = n948 | n3003 ;
  assign n3009 = ( ~n332 & n1187 ) | ( ~n332 & n3005 ) | ( n1187 & n3005 ) ;
  assign n3010 = n332 | n3009 ;
  assign n3011 = ( ~n165 & n607 ) | ( ~n165 & n3010 ) | ( n607 & n3010 ) ;
  assign n3012 = n651 | n2821 ;
  assign n3013 = n165 | n3011 ;
  assign n3014 = n3007 | n3012 ;
  assign n3015 = ( n94 & ~n294 ) | ( n94 & n3013 ) | ( ~n294 & n3013 ) ;
  assign n3016 = n294 | n3015 ;
  assign n3017 = n146 | n3016 ;
  assign n3018 = n954 | n3017 ;
  assign n3019 = n1442 & ~n3017 ;
  assign n3020 = n2868 | n3014 ;
  assign n3021 = n241 | n2635 ;
  assign n3022 = n1059 | n2837 ;
  assign n3023 = n3021 | n3022 ;
  assign n3024 = n1035 | n2488 ;
  assign n3025 = n2300 | n2488 ;
  assign n3026 = n3023 | n3025 ;
  assign n3027 = n2627 & ~n2695 ;
  assign n3028 = ~n3018 & n3027 ;
  assign n3029 = n357 | n963 ;
  assign n3030 = ( n426 & ~n520 ) | ( n426 & n3026 ) | ( ~n520 & n3026 ) ;
  assign n3031 = n520 | n3030 ;
  assign n3032 = ( ~n381 & n3029 ) | ( ~n381 & n3031 ) | ( n3029 & n3031 ) ;
  assign n3033 = n381 | n3032 ;
  assign n3034 = n2235 | n3033 ;
  assign n3035 = n3019 & ~n3034 ;
  assign n3036 = ~n2938 & n3035 ;
  assign n3037 = n501 | n841 ;
  assign n3038 = n169 | n422 ;
  assign n3039 = n3037 | n3038 ;
  assign n3040 = n547 | n945 ;
  assign n3041 = n444 | n3040 ;
  assign n3042 = n1227 & ~n2998 ;
  assign n3043 = ~n3008 & n3042 ;
  assign n3044 = n536 | n3041 ;
  assign n3045 = n1992 | n3041 ;
  assign n3046 = n559 | n3020 ;
  assign n3047 = n3039 | n3045 ;
  assign n3048 = n785 | n3047 ;
  assign n3049 = ( n1366 & ~n3033 ) | ( n1366 & n3047 ) | ( ~n3033 & n3047 ) ;
  assign n3050 = n3033 | n3049 ;
  assign n3051 = n2627 & ~n3050 ;
  assign n3052 = n628 | n862 ;
  assign n3053 = n139 | n248 ;
  assign n3054 = n371 | n3053 ;
  assign n3055 = n107 | n122 ;
  assign n3056 = n287 | n834 ;
  assign n3057 = n3052 | n3056 ;
  assign n3058 = n3055 | n3057 ;
  assign n3059 = n532 | n601 ;
  assign n3060 = n887 | n955 ;
  assign n3061 = n3059 | n3060 ;
  assign n3062 = n93 | n3054 ;
  assign n3063 = n977 | n3054 ;
  assign n3064 = n3061 | n3062 ;
  assign n3065 = n173 | n437 ;
  assign n3066 = n1403 | n3058 ;
  assign n3067 = n2316 | n3066 ;
  assign n3068 = n2992 | n3065 ;
  assign n3069 = n548 | n2992 ;
  assign n3070 = ( ~n2909 & n3064 ) | ( ~n2909 & n3067 ) | ( n3064 & n3067 ) ;
  assign n3071 = n2909 | n3070 ;
  assign n3072 = ( ~n86 & n258 ) | ( ~n86 & n3071 ) | ( n258 & n3071 ) ;
  assign n3073 = n86 | n3072 ;
  assign n3074 = ( n255 & ~n288 ) | ( n255 & n3073 ) | ( ~n288 & n3073 ) ;
  assign n3075 = n288 | n3074 ;
  assign n3076 = ( n829 & ~n941 ) | ( n829 & n3075 ) | ( ~n941 & n3075 ) ;
  assign n3077 = n941 | n3076 ;
  assign n3078 = n2996 | n3077 ;
  assign n3079 = n3068 | n3078 ;
  assign n3080 = n294 | n336 ;
  assign n3081 = n2750 | n3079 ;
  assign n3082 = n3056 | n3065 ;
  assign n3083 = n3044 | n3082 ;
  assign n3084 = n1083 | n2512 ;
  assign n3085 = n3069 | n3084 ;
  assign n3086 = n285 | n534 ;
  assign n3087 = n3080 | n3086 ;
  assign n3088 = n2564 | n3087 ;
  assign n3089 = n3077 | n3087 ;
  assign n3090 = n345 | n943 ;
  assign n3091 = n3048 | n3089 ;
  assign n3092 = n2879 | n3090 ;
  assign n3093 = n3088 | n3092 ;
  assign n3094 = n2770 | n3093 ;
  assign n3095 = n147 | n375 ;
  assign n3096 = n2512 | n3056 ;
  assign n3097 = n300 | n744 ;
  assign n3098 = n3052 | n3097 ;
  assign n3099 = n3065 | n3098 ;
  assign n3100 = n1903 | n3099 ;
  assign n3101 = n247 | n810 ;
  assign n3102 = n1192 | n3058 ;
  assign n3103 = n3095 | n3101 ;
  assign n3104 = n352 | n645 ;
  assign n3105 = n3096 | n3103 ;
  assign n3106 = ( n235 & n583 ) | ( n235 & ~n3105 ) | ( n583 & ~n3105 ) ;
  assign n3107 = n235 | n295 ;
  assign n3108 = n731 | n3107 ;
  assign n3109 = n3002 | n3108 ;
  assign n3110 = ~n235 & n3106 ;
  assign n3111 = n3104 | n3108 ;
  assign n3112 = n84 | n2446 ;
  assign n3113 = n3111 | n3112 ;
  assign n3114 = n2934 | n3113 ;
  assign n3115 = n3085 | n3114 ;
  assign n3116 = ( n2086 & ~n3064 ) | ( n2086 & n3115 ) | ( ~n3064 & n3115 ) ;
  assign n3117 = n3064 | n3116 ;
  assign n3118 = n555 | n2246 ;
  assign n3119 = n342 | n373 ;
  assign n3120 = n360 | n631 ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = n90 | n1798 ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = n589 | n647 ;
  assign n3125 = ( ~n2549 & n2968 ) | ( ~n2549 & n3123 ) | ( n2968 & n3123 ) ;
  assign n3126 = n2549 | n3125 ;
  assign n3127 = n358 | n422 ;
  assign n3128 = ( ~n105 & n336 ) | ( ~n105 & n3126 ) | ( n336 & n3126 ) ;
  assign n3129 = n105 | n3128 ;
  assign n3130 = ( ~n461 & n546 ) | ( ~n461 & n3129 ) | ( n546 & n3129 ) ;
  assign n3131 = n461 | n3130 ;
  assign n3132 = n149 | n417 ;
  assign n3133 = n3127 | n3132 ;
  assign n3134 = n3124 | n3133 ;
  assign n3135 = n1089 | n3118 ;
  assign n3136 = n3131 | n3132 ;
  assign n3137 = n3080 | n3135 ;
  assign n3138 = n2722 | n3134 ;
  assign n3139 = n255 | n593 ;
  assign n3140 = n651 | n3080 ;
  assign n3141 = ( n578 & ~n645 ) | ( n578 & n3136 ) | ( ~n645 & n3136 ) ;
  assign n3142 = n2831 | n3141 ;
  assign n3143 = n842 | n3142 ;
  assign n3144 = n1305 & ~n3133 ;
  assign n3145 = n2372 | n3135 ;
  assign n3146 = n2372 | n3140 ;
  assign n3147 = n2647 | n3140 ;
  assign n3148 = n3144 & ~n3147 ;
  assign n3149 = n715 | n1307 ;
  assign n3150 = n3120 | n3149 ;
  assign n3151 = n1676 | n3139 ;
  assign n3152 = n3137 | n3151 ;
  assign n3153 = n1085 | n3150 ;
  assign n3154 = n3152 | n3153 ;
  assign n3155 = ( n428 & ~n1697 ) | ( n428 & n3154 ) | ( ~n1697 & n3154 ) ;
  assign n3156 = n790 | n891 ;
  assign n3157 = n1697 | n3155 ;
  assign n3158 = n111 | n220 ;
  assign n3159 = n3156 | n3158 ;
  assign n3160 = ( n306 & ~n2939 ) | ( n306 & n3157 ) | ( ~n2939 & n3157 ) ;
  assign n3161 = n870 & ~n1059 ;
  assign n3162 = ~n3143 & n3161 ;
  assign n3163 = n1305 & ~n1622 ;
  assign n3164 = ( n555 & ~n757 ) | ( n555 & n3138 ) | ( ~n757 & n3138 ) ;
  assign n3165 = n2671 | n3159 ;
  assign n3166 = n2939 | n3160 ;
  assign n3167 = n3162 & ~n3165 ;
  assign n3168 = ( ~n105 & n825 ) | ( ~n105 & n3166 ) | ( n825 & n3166 ) ;
  assign n3169 = n105 | n3168 ;
  assign n3170 = n164 | n849 ;
  assign n3171 = n605 | n3159 ;
  assign n3172 = n3170 | n3171 ;
  assign n3173 = n1244 | n2841 ;
  assign n3174 = ( ~n559 & n969 ) | ( ~n559 & n3169 ) | ( n969 & n3169 ) ;
  assign n3175 = n128 | n154 ;
  assign n3176 = n1676 | n3175 ;
  assign n3177 = n1806 | n3174 ;
  assign n3178 = n3173 | n3176 ;
  assign n3179 = ( ~n1454 & n2499 ) | ( ~n1454 & n3177 ) | ( n2499 & n3177 ) ;
  assign n3180 = n1454 | n3179 ;
  assign n3181 = n3046 | n3174 ;
  assign n3182 = n3102 | n3172 ;
  assign n3183 = n2001 | n2227 ;
  assign n3184 = n3182 | n3183 ;
  assign n3185 = n757 | n3164 ;
  assign n3186 = n2841 | n3150 ;
  assign n3187 = n88 | n967 ;
  assign n3188 = n759 | n3187 ;
  assign n3189 = n82 | n125 ;
  assign n3190 = n561 | n1860 ;
  assign n3191 = n169 | n415 ;
  assign n3192 = n3188 | n3189 ;
  assign n3193 = n3191 | n3192 ;
  assign n3194 = n111 | n2551 ;
  assign n3195 = n448 | n3194 ;
  assign n3196 = n3190 | n3193 ;
  assign n3197 = n86 | n434 ;
  assign n3198 = n283 | n503 ;
  assign n3199 = n2802 | n3196 ;
  assign n3200 = ( n794 & ~n2329 ) | ( n794 & n3199 ) | ( ~n2329 & n3199 ) ;
  assign n3201 = n147 | n846 ;
  assign n3202 = n124 | n969 ;
  assign n3203 = n3198 | n3201 ;
  assign n3204 = n1087 | n2589 ;
  assign n3205 = n3197 | n3203 ;
  assign n3206 = n953 | n3205 ;
  assign n3207 = n350 | n1661 ;
  assign n3208 = n1087 | n2694 ;
  assign n3209 = n425 | n3202 ;
  assign n3210 = n1661 | n3209 ;
  assign n3211 = n247 | n3209 ;
  assign n3212 = n1288 | n3211 ;
  assign n3213 = n1529 | n3206 ;
  assign n3214 = n3208 | n3213 ;
  assign n3215 = n3195 | n3212 ;
  assign n3216 = n3214 | n3215 ;
  assign n3217 = ( ~n180 & n561 ) | ( ~n180 & n3216 ) | ( n561 & n3216 ) ;
  assign n3218 = n180 | n3217 ;
  assign n3219 = ( ~n420 & n1712 ) | ( ~n420 & n3218 ) | ( n1712 & n3218 ) ;
  assign n3220 = n206 | n829 ;
  assign n3221 = n2923 | n3220 ;
  assign n3222 = n420 | n3219 ;
  assign n3223 = ( n367 & ~n788 ) | ( n367 & n3222 ) | ( ~n788 & n3222 ) ;
  assign n3224 = n788 | n3223 ;
  assign n3225 = n203 | n3224 ;
  assign n3226 = ( ~n1243 & n2764 ) | ( ~n1243 & n3225 ) | ( n2764 & n3225 ) ;
  assign n3227 = n3142 | n3225 ;
  assign n3228 = ~n3225 & n3226 ;
  assign n3229 = n494 | n3220 ;
  assign n3230 = n2045 | n3229 ;
  assign n3231 = n223 | n3220 ;
  assign n3232 = n1285 | n3231 ;
  assign n3233 = n222 | n660 ;
  assign n3234 = n601 | n3232 ;
  assign n3235 = n3220 | n3233 ;
  assign n3236 = n3028 & ~n3235 ;
  assign n3237 = n2795 | n3233 ;
  assign n3238 = n3193 | n3227 ;
  assign n3239 = n3063 | n3238 ;
  assign n3240 = n344 | n2266 ;
  assign n3241 = ( n966 & ~n1745 ) | ( n966 & n3239 ) | ( ~n1745 & n3239 ) ;
  assign n3242 = n631 | n693 ;
  assign n3243 = n313 | n1019 ;
  assign n3244 = n3240 | n3242 ;
  assign n3245 = n1245 | n3244 ;
  assign n3246 = n3237 | n3243 ;
  assign n3247 = n3245 | n3246 ;
  assign n3248 = ( ~n125 & n1774 ) | ( ~n125 & n3247 ) | ( n1774 & n3247 ) ;
  assign n3249 = n116 | n1192 ;
  assign n3250 = n585 | n731 ;
  assign n3251 = n286 | n3249 ;
  assign n3252 = n288 | n593 ;
  assign n3253 = n246 | n306 ;
  assign n3254 = n3252 | n3253 ;
  assign n3255 = n371 | n955 ;
  assign n3256 = n3250 | n3255 ;
  assign n3257 = ( ~n1894 & n2367 ) | ( ~n1894 & n3256 ) | ( n2367 & n3256 ) ;
  assign n3258 = ~n3256 & n3257 ;
  assign n3259 = ~n1566 & n3258 ;
  assign n3260 = n473 | n2837 ;
  assign n3261 = n473 | n3233 ;
  assign n3262 = n3251 | n3261 ;
  assign n3263 = n2776 | n3262 ;
  assign n3264 = n161 | n336 ;
  assign n3265 = n3254 | n3264 ;
  assign n3266 = n184 | n348 ;
  assign n3267 = ( n210 & ~n442 ) | ( n210 & n3265 ) | ( ~n442 & n3265 ) ;
  assign n3268 = n442 | n3267 ;
  assign n3269 = ( ~n1146 & n3263 ) | ( ~n1146 & n3268 ) | ( n3263 & n3268 ) ;
  assign n3270 = n1146 | n3269 ;
  assign n3271 = ( n550 & ~n3266 ) | ( n550 & n3270 ) | ( ~n3266 & n3270 ) ;
  assign n3272 = n3266 | n3271 ;
  assign n3273 = ( ~n101 & n3250 ) | ( ~n101 & n3272 ) | ( n3250 & n3272 ) ;
  assign n3274 = n101 | n3273 ;
  assign n3275 = ( ~n649 & n1333 ) | ( ~n649 & n3274 ) | ( n1333 & n3274 ) ;
  assign n3276 = n649 | n3275 ;
  assign n3277 = n1465 | n3276 ;
  assign n3278 = n348 | n786 ;
  assign n3279 = n910 | n3276 ;
  assign n3280 = n105 | n3278 ;
  assign n3281 = n2277 | n3280 ;
  assign n3282 = n2670 | n3256 ;
  assign n3283 = n3281 | n3282 ;
  assign n3284 = ( ~n207 & n349 ) | ( ~n207 & n3283 ) | ( n349 & n3283 ) ;
  assign n3285 = n207 | n3284 ;
  assign n3286 = ( ~n145 & n965 ) | ( ~n145 & n3285 ) | ( n965 & n3285 ) ;
  assign n3287 = n145 | n3286 ;
  assign n3288 = ( n416 & ~n555 ) | ( n416 & n3287 ) | ( ~n555 & n3287 ) ;
  assign n3289 = n555 | n3288 ;
  assign n3290 = n206 | n3289 ;
  assign n3291 = n1508 | n3290 ;
  assign n3292 = n1783 | n3291 ;
  assign n3293 = n214 | n1051 ;
  assign n3294 = n3260 | n3292 ;
  assign n3295 = n607 | n693 ;
  assign n3296 = n3293 | n3295 ;
  assign n3297 = n345 | n2127 ;
  assign n3298 = n3296 | n3297 ;
  assign n3299 = n717 | n3298 ;
  assign n3300 = n3290 | n3299 ;
  assign n3301 = n204 | n3300 ;
  assign n3302 = n2112 | n3301 ;
  assign n3303 = n532 | n1136 ;
  assign n3304 = ( ~n82 & n3302 ) | ( ~n82 & n3303 ) | ( n3302 & n3303 ) ;
  assign n3305 = n82 | n3304 ;
  assign n3306 = ( ~n522 & n754 ) | ( ~n522 & n3305 ) | ( n754 & n3305 ) ;
  assign n3307 = n522 | n3306 ;
  assign n3308 = ( n497 & ~n719 ) | ( n497 & n3307 ) | ( ~n719 & n3307 ) ;
  assign n3309 = n719 | n3308 ;
  assign n3310 = ( n188 & ~n651 ) | ( n188 & n3309 ) | ( ~n651 & n3309 ) ;
  assign n3311 = n2595 | n3310 ;
  assign n3312 = n2045 | n3311 ;
  assign n3313 = n3146 | n3312 ;
  assign n3314 = ( n2801 & ~n3206 ) | ( n2801 & n3313 ) | ( ~n3206 & n3313 ) ;
  assign n3315 = n3206 | n3314 ;
  assign n3316 = n362 | n372 ;
  assign n3317 = n168 | n955 ;
  assign n3318 = n336 | n3316 ;
  assign n3319 = n2694 | n3318 ;
  assign n3320 = n1587 | n3319 ;
  assign n3321 = n757 | n3317 ;
  assign n3322 = n84 | n245 ;
  assign n3323 = n122 | n145 ;
  assign n3324 = n3322 | n3323 ;
  assign n3325 = n183 | n1846 ;
  assign n3326 = n3324 | n3325 ;
  assign n3327 = n3321 | n3326 ;
  assign n3328 = n3320 | n3327 ;
  assign n3329 = ( n456 & ~n565 ) | ( n456 & n3328 ) | ( ~n565 & n3328 ) ;
  assign n3330 = n88 | n1088 ;
  assign n3331 = n565 | n3329 ;
  assign n3332 = ( n154 & ~n693 ) | ( n154 & n3331 ) | ( ~n693 & n3331 ) ;
  assign n3333 = n693 | n3332 ;
  assign n3334 = ( n872 & ~n923 ) | ( n872 & n3333 ) | ( ~n923 & n3333 ) ;
  assign n3335 = n1740 | n3330 ;
  assign n3336 = n390 | n3334 ;
  assign n3337 = n2508 | n3334 ;
  assign n3338 = n234 | n532 ;
  assign n3339 = n3335 | n3338 ;
  assign n3340 = n229 | n862 ;
  assign n3341 = n612 | n3340 ;
  assign n3342 = n2095 | n3318 ;
  assign n3343 = n1204 | n3341 ;
  assign n3344 = n3339 | n3343 ;
  assign n3345 = ( ~n175 & n1333 ) | ( ~n175 & n3344 ) | ( n1333 & n3344 ) ;
  assign n3346 = n2694 | n3185 ;
  assign n3347 = n175 | n3345 ;
  assign n3348 = n93 | n653 ;
  assign n3349 = n3321 | n3348 ;
  assign n3350 = n1370 | n3349 ;
  assign n3351 = n3341 | n3348 ;
  assign n3352 = n3178 | n3351 ;
  assign n3353 = n608 | n715 ;
  assign n3354 = n249 | n2957 ;
  assign n3355 = ( n271 & ~n953 ) | ( n271 & n3347 ) | ( ~n953 & n3347 ) ;
  assign n3356 = n2447 | n3342 ;
  assign n3357 = n3354 | n3356 ;
  assign n3358 = n133 | n3353 ;
  assign n3359 = n224 | n585 ;
  assign n3360 = n953 | n3355 ;
  assign n3361 = ( n3185 & n3236 ) | ( n3185 & ~n3360 ) | ( n3236 & ~n3360 ) ;
  assign n3362 = n3358 | n3360 ;
  assign n3363 = n2533 | n3362 ;
  assign n3364 = n1770 | n3359 ;
  assign n3365 = n1770 | n2127 ;
  assign n3366 = n249 | n2429 ;
  assign n3367 = n559 | n3359 ;
  assign n3368 = n3366 | n3367 ;
  assign n3369 = n2882 | n3363 ;
  assign n3370 = n2629 | n3368 ;
  assign n3371 = ~n3185 & n3361 ;
  assign n3372 = n81 | n250 ;
  assign n3373 = n414 | n3372 ;
  assign n3374 = n1186 | n3373 ;
  assign n3375 = n2877 & ~n3374 ;
  assign n3376 = n183 | n1552 ;
  assign n3377 = n86 | n91 ;
  assign n3378 = n3376 | n3377 ;
  assign n3379 = n341 | n416 ;
  assign n3380 = n149 | n3379 ;
  assign n3381 = n3373 | n3380 ;
  assign n3382 = n3378 | n3381 ;
  assign n3383 = ( n247 & ~n279 ) | ( n247 & n3382 ) | ( ~n279 & n3382 ) ;
  assign n3384 = n279 | n3383 ;
  assign n3385 = n367 | n3384 ;
  assign n3386 = n843 | n3385 ;
  assign n3387 = n702 | n1577 ;
  assign n3388 = n343 | n3387 ;
  assign n3389 = n3364 | n3386 ;
  assign n3390 = n288 | n547 ;
  assign n3391 = n846 | n3390 ;
  assign n3392 = n3326 | n3388 ;
  assign n3393 = n3388 | n3391 ;
  assign n3394 = n2854 | n3393 ;
  assign n3395 = n172 | n210 ;
  assign n3396 = n1170 | n3394 ;
  assign n3397 = n1156 | n3380 ;
  assign n3398 = n1156 | n1666 ;
  assign n3399 = n715 | n963 ;
  assign n3400 = n587 | n3399 ;
  assign n3401 = n3395 | n3400 ;
  assign n3402 = n1552 | n3233 ;
  assign n3403 = n375 | n3175 ;
  assign n3404 = n3359 | n3401 ;
  assign n3405 = n279 | n1666 ;
  assign n3406 = n3404 | n3405 ;
  assign n3407 = n294 | n832 ;
  assign n3408 = n361 | n3407 ;
  assign n3409 = n1186 | n3408 ;
  assign n3410 = n1026 | n3408 ;
  assign n3411 = n182 | n3403 ;
  assign n3412 = n2763 | n3411 ;
  assign n3413 = n3409 | n3412 ;
  assign n3414 = n400 | n605 ;
  assign n3415 = n105 | n367 ;
  assign n3416 = n3414 | n3415 ;
  assign n3417 = n659 | n3415 ;
  assign n3418 = n3402 | n3417 ;
  assign n3419 = n1634 | n3417 ;
  assign n3420 = n2991 | n3416 ;
  assign n3421 = n2113 | n3420 ;
  assign n3422 = n83 | n97 ;
  assign n3423 = n1514 | n3422 ;
  assign n3424 = n902 | n3423 ;
  assign n3425 = n3406 | n3424 ;
  assign n3426 = n360 | n3337 ;
  assign n3427 = n617 | n3423 ;
  assign n3428 = n3421 | n3427 ;
  assign n3429 = n175 | n578 ;
  assign n3430 = n735 | n961 ;
  assign n3431 = n293 | n3429 ;
  assign n3432 = n3430 | n3431 ;
  assign n3433 = n1497 | n3330 ;
  assign n3434 = n3432 | n3433 ;
  assign n3435 = n3398 | n3432 ;
  assign n3436 = n1897 | n3434 ;
  assign n3437 = n221 | n628 ;
  assign n3438 = n304 | n552 ;
  assign n3439 = n3437 | n3438 ;
  assign n3440 = n182 | n841 ;
  assign n3441 = n3439 | n3440 ;
  assign n3442 = n713 | n942 ;
  assign n3443 = n3330 | n3442 ;
  assign n3444 = n3397 | n3443 ;
  assign n3445 = ( ~n678 & n3441 ) | ( ~n678 & n3444 ) | ( n3441 & n3444 ) ;
  assign n3446 = n3110 & ~n3445 ;
  assign n3447 = n420 | n841 ;
  assign n3448 = ~n678 & n3446 ;
  assign n3449 = n103 | n306 ;
  assign n3450 = n3447 | n3449 ;
  assign n3451 = n286 | n415 ;
  assign n3452 = n3450 | n3451 ;
  assign n3453 = ( ~n757 & n3436 ) | ( ~n757 & n3452 ) | ( n3436 & n3452 ) ;
  assign n3454 = n2991 | n3452 ;
  assign n3455 = n228 | n318 ;
  assign n3456 = n731 | n1738 ;
  assign n3457 = n3455 | n3456 ;
  assign n3458 = n757 | n3453 ;
  assign n3459 = n651 | n3458 ;
  assign n3460 = n3310 | n3459 ;
  assign n3461 = n580 | n942 ;
  assign n3462 = n2994 | n3461 ;
  assign n3463 = n3457 | n3462 ;
  assign n3464 = ( n502 & ~n943 ) | ( n502 & n3463 ) | ( ~n943 & n3463 ) ;
  assign n3465 = n943 | n3464 ;
  assign n3466 = ( ~n417 & n778 ) | ( ~n417 & n3465 ) | ( n778 & n3465 ) ;
  assign n3467 = n417 | n3466 ;
  assign n3468 = ( n89 & ~n651 ) | ( n89 & n3467 ) | ( ~n651 & n3467 ) ;
  assign n3469 = n651 | n3468 ;
  assign n3470 = n3188 | n3469 ;
  assign n3471 = n2424 & ~n3470 ;
  assign n3472 = n3441 | n3469 ;
  assign n3473 = ( ~n555 & n1379 ) | ( ~n555 & n3471 ) | ( n1379 & n3471 ) ;
  assign n3474 = n91 | n296 ;
  assign n3475 = n169 | n3090 ;
  assign n3476 = n628 | n715 ;
  assign n3477 = n3475 | n3476 ;
  assign n3478 = n757 | n3477 ;
  assign n3479 = n3391 | n3478 ;
  assign n3480 = n3454 | n3479 ;
  assign n3481 = n578 | n841 ;
  assign n3482 = ( ~n651 & n2647 ) | ( ~n651 & n3480 ) | ( n2647 & n3480 ) ;
  assign n3483 = n318 | n422 ;
  assign n3484 = n3477 | n3483 ;
  assign n3485 = n788 | n3474 ;
  assign n3486 = n2807 | n3484 ;
  assign n3487 = n362 | n444 ;
  assign n3488 = n3024 | n3486 ;
  assign n3489 = n2961 | n3487 ;
  assign n3490 = n3435 | n3489 ;
  assign n3491 = n116 | n719 ;
  assign n3492 = ( ~n850 & n2809 ) | ( ~n850 & n3491 ) | ( n2809 & n3491 ) ;
  assign n3493 = n850 | n3492 ;
  assign n3494 = ( ~n1230 & n2909 ) | ( ~n1230 & n3493 ) | ( n2909 & n3493 ) ;
  assign n3495 = n1230 | n3494 ;
  assign n3496 = ( ~n367 & n759 ) | ( ~n367 & n3495 ) | ( n759 & n3495 ) ;
  assign n3497 = n367 | n3496 ;
  assign n3498 = ( n697 & ~n2937 ) | ( n697 & n3490 ) | ( ~n2937 & n3490 ) ;
  assign n3499 = ( ~n271 & n2792 ) | ( ~n271 & n3497 ) | ( n2792 & n3497 ) ;
  assign n3500 = ~n3497 & n3499 ;
  assign n3501 = n271 | n3481 ;
  assign n3502 = n3485 | n3497 ;
  assign n3503 = n3501 | n3502 ;
  assign n3504 = n1603 | n3503 ;
  assign n3505 = ( n1686 & ~n1833 ) | ( n1686 & n3504 ) | ( ~n1833 & n3504 ) ;
  assign n3506 = n1833 | n3505 ;
  assign n3507 = ( ~n2041 & n3483 ) | ( ~n2041 & n3506 ) | ( n3483 & n3506 ) ;
  assign n3508 = n2041 | n3507 ;
  assign n3509 = ( n1754 & ~n2329 ) | ( n1754 & n3508 ) | ( ~n2329 & n3508 ) ;
  assign n3510 = ~n1621 & n3500 ;
  assign n3511 = n585 | n608 ;
  assign n3512 = n448 | n3511 ;
  assign n3513 = n499 | n786 ;
  assign n3514 = n3512 | n3513 ;
  assign n3515 = n2404 | n3514 ;
  assign n3516 = n125 | n969 ;
  assign n3517 = n702 | n3515 ;
  assign n3518 = n705 | n3517 ;
  assign n3519 = n86 | n164 ;
  assign n3520 = ( n1844 & n3477 ) | ( n1844 & ~n3512 ) | ( n3477 & ~n3512 ) ;
  assign n3521 = n3516 | n3519 ;
  assign n3522 = n245 | n250 ;
  assign n3523 = n3277 | n3521 ;
  assign n3524 = n1460 | n3487 ;
  assign n3525 = n2223 | n3522 ;
  assign n3526 = n3524 | n3525 ;
  assign n3527 = n225 | n757 ;
  assign n3528 = n1035 | n3527 ;
  assign n3529 = ( n2837 & n3228 ) | ( n2837 & ~n3481 ) | ( n3228 & ~n3481 ) ;
  assign n3530 = n3472 | n3526 ;
  assign n3531 = n3513 | n3528 ;
  assign n3532 = n3523 | n3531 ;
  assign n3533 = n206 | n647 ;
  assign n3534 = ( ~n785 & n3234 ) | ( ~n785 & n3530 ) | ( n3234 & n3530 ) ;
  assign n3535 = ( ~n1958 & n3234 ) | ( ~n1958 & n3532 ) | ( n3234 & n3532 ) ;
  assign n3536 = n1045 | n3533 ;
  assign n3537 = n3109 | n3536 ;
  assign n3538 = ~n1733 & n3510 ;
  assign n3539 = n81 | n754 ;
  assign n3540 = n1958 | n3535 ;
  assign n3541 = n1733 | n3006 ;
  assign n3542 = ( ~n98 & n3448 ) | ( ~n98 & n3539 ) | ( n3448 & n3539 ) ;
  assign n3543 = ~n3539 & n3542 ;
  assign n3544 = ( n229 & ~n825 ) | ( n229 & n3543 ) | ( ~n825 & n3543 ) ;
  assign n3545 = ~n229 & n3544 ;
  assign n3546 = ( n209 & ~n381 ) | ( n209 & n3545 ) | ( ~n381 & n3545 ) ;
  assign n3547 = n203 | n342 ;
  assign n3548 = ~n209 & n3546 ;
  assign n3549 = ( ~n3123 & n3540 ) | ( ~n3123 & n3548 ) | ( n3540 & n3548 ) ;
  assign n3550 = ~n3540 & n3549 ;
  assign n3551 = ~n2837 & n3529 ;
  assign n3552 = n234 | n796 ;
  assign n3553 = n2939 | n3547 ;
  assign n3554 = n2837 | n3533 ;
  assign n3555 = n3552 | n3553 ;
  assign n3556 = ~n530 & n3548 ;
  assign n3557 = ~n1338 & n3556 ;
  assign n3558 = ~n3533 & n3557 ;
  assign n3559 = ~n2970 & n3558 ;
  assign n3560 = ~n2270 & n3559 ;
  assign n3561 = ( n2829 & ~n3555 ) | ( n2829 & n3560 ) | ( ~n3555 & n3560 ) ;
  assign n3562 = n149 | n1111 ;
  assign n3563 = ~n2829 & n3561 ;
  assign n3564 = ( ~n1388 & n3268 ) | ( ~n1388 & n3563 ) | ( n3268 & n3563 ) ;
  assign n3565 = ~n3268 & n3564 ;
  assign n3566 = ~n1083 & n3565 ;
  assign n3567 = n701 | n3562 ;
  assign n3568 = n224 | n349 ;
  assign n3569 = n304 | n3568 ;
  assign n3570 = ( ~n1512 & n2909 ) | ( ~n1512 & n3537 ) | ( n2909 & n3537 ) ;
  assign n3571 = n2970 | n3569 ;
  assign n3572 = n2425 | n3571 ;
  assign n3573 = n3541 | n3572 ;
  assign n3574 = n3567 | n3569 ;
  assign n3575 = n2818 | n3569 ;
  assign n3576 = n1952 | n3574 ;
  assign n3577 = ( ~n256 & n3555 ) | ( ~n256 & n3576 ) | ( n3555 & n3576 ) ;
  assign n3578 = n256 | n3577 ;
  assign n3579 = n702 | n891 ;
  assign n3580 = n608 | n2879 ;
  assign n3581 = n1145 | n2507 ;
  assign n3582 = n644 | n1192 ;
  assign n3583 = n341 | n3491 ;
  assign n3584 = ( ~n608 & n3579 ) | ( ~n608 & n3583 ) | ( n3579 & n3583 ) ;
  assign n3585 = n1512 | n3570 ;
  assign n3586 = n351 | n965 ;
  assign n3587 = n813 | n3584 ;
  assign n3588 = n3580 | n3581 ;
  assign n3589 = n825 | n3582 ;
  assign n3590 = n2593 | n3589 ;
  assign n3591 = n3588 | n3590 ;
  assign n3592 = n3584 | n3591 ;
  assign n3593 = n552 | n649 ;
  assign n3594 = ( ~n1045 & n1920 ) | ( ~n1045 & n3592 ) | ( n1920 & n3592 ) ;
  assign n3595 = n1045 | n3594 ;
  assign n3596 = n1723 | n3593 ;
  assign n3597 = n3512 | n3520 ;
  assign n3598 = ~n1379 & n3473 ;
  assign n3599 = n94 | n437 ;
  assign n3600 = n3596 | n3599 ;
  assign n3601 = n1492 | n3600 ;
  assign n3602 = n1818 | n3442 ;
  assign n3603 = n3163 & ~n3602 ;
  assign n3604 = n282 | n1354 ;
  assign n3605 = n607 | n3604 ;
  assign n3606 = n1723 | n3604 ;
  assign n3607 = n306 | n3586 ;
  assign n3608 = ( ~n281 & n422 ) | ( ~n281 & n3585 ) | ( n422 & n3585 ) ;
  assign n3609 = n1431 | n3605 ;
  assign n3610 = n281 | n3608 ;
  assign n3611 = ( ~n306 & n2324 ) | ( ~n306 & n3597 ) | ( n2324 & n3597 ) ;
  assign n3612 = n306 | n3611 ;
  assign n3613 = ( ~n427 & n658 ) | ( ~n427 & n3610 ) | ( n658 & n3610 ) ;
  assign n3614 = ( ~n605 & n1333 ) | ( ~n605 & n3612 ) | ( n1333 & n3612 ) ;
  assign n3615 = n427 | n3613 ;
  assign n3616 = n3603 & ~n3609 ;
  assign n3617 = n153 | n1777 ;
  assign n3618 = n3606 | n3617 ;
  assign n3619 = n1304 | n3618 ;
  assign n3620 = n530 | n3522 ;
  assign n3621 = n1312 | n1593 ;
  assign n3622 = n555 | n1379 ;
  assign n3623 = n3589 | n3615 ;
  assign n3624 = n3620 | n3621 ;
  assign n3625 = n303 | n593 ;
  assign n3626 = n3623 | n3624 ;
  assign n3627 = n125 | n209 ;
  assign n3628 = n645 | n3626 ;
  assign n3629 = n3607 | n3627 ;
  assign n3630 = n756 | n3625 ;
  assign n3631 = n3141 | n3628 ;
  assign n3632 = n608 | n3593 ;
  assign n3633 = n3485 | n3629 ;
  assign n3634 = n3629 | n3630 ;
  assign n3635 = n3632 | n3634 ;
  assign n3636 = n3587 | n3635 ;
  assign n3637 = n183 | n945 ;
  assign n3638 = ( ~n82 & n2990 ) | ( ~n82 & n3637 ) | ( n2990 & n3637 ) ;
  assign n3639 = n2957 | n3636 ;
  assign n3640 = n82 | n3638 ;
  assign n3641 = ( ~n1973 & n3622 ) | ( ~n1973 & n3639 ) | ( n3622 & n3639 ) ;
  assign n3642 = n1973 | n3641 ;
  assign n3643 = ( ~n234 & n250 ) | ( ~n234 & n3640 ) | ( n250 & n3640 ) ;
  assign n3644 = ( n115 & ~n888 ) | ( n115 & n3642 ) | ( ~n888 & n3642 ) ;
  assign n3645 = ( ~n1111 & n3184 ) | ( ~n1111 & n3637 ) | ( n3184 & n3637 ) ;
  assign n3646 = n1111 | n3645 ;
  assign n3647 = n888 | n3644 ;
  assign n3648 = ( ~n295 & n1111 ) | ( ~n295 & n3647 ) | ( n1111 & n3647 ) ;
  assign n3649 = n234 | n3643 ;
  assign n3650 = n502 | n3649 ;
  assign n3651 = n605 | n3614 ;
  assign n3652 = n290 | n490 ;
  assign n3653 = n969 | n3652 ;
  assign n3654 = n1497 | n3652 ;
  assign n3655 = n1248 | n3653 ;
  assign n3656 = n583 & ~n953 ;
  assign n3657 = ~n1193 & n3656 ;
  assign n3658 = ~n3655 & n3657 ;
  assign n3659 = ~n3207 & n3658 ;
  assign n3660 = n177 | n943 ;
  assign n3661 = n416 | n3660 ;
  assign n3662 = ( ~n360 & n701 ) | ( ~n360 & n3651 ) | ( n701 & n3651 ) ;
  assign n3663 = n3426 | n3662 ;
  assign n3664 = n360 | n3662 ;
  assign n3665 = ( ~n270 & n3659 ) | ( ~n270 & n3664 ) | ( n3659 & n3664 ) ;
  assign n3666 = n1258 | n1381 ;
  assign n3667 = n3655 | n3666 ;
  assign n3668 = n3605 | n3666 ;
  assign n3669 = n3661 | n3666 ;
  assign n3670 = n3244 | n3586 ;
  assign n3671 = n3100 | n3667 ;
  assign n3672 = n223 | n3487 ;
  assign n3673 = ~n1398 & n3656 ;
  assign n3674 = ~n3661 & n3673 ;
  assign n3675 = ~n3670 & n3674 ;
  assign n3676 = n2512 | n3607 ;
  assign n3677 = n188 | n372 ;
  assign n3678 = n3637 | n3677 ;
  assign n3679 = n341 | n3678 ;
  assign n3680 = n3411 | n3679 ;
  assign n3681 = n649 | n955 ;
  assign n3682 = n747 | n3681 ;
  assign n3683 = n3139 | n3678 ;
  assign n3684 = n3676 | n3682 ;
  assign n3685 = n3668 | n3684 ;
  assign n3686 = n228 | n422 ;
  assign n3687 = n3683 | n3686 ;
  assign n3688 = ( ~n961 & n1879 ) | ( ~n961 & n3595 ) | ( n1879 & n3595 ) ;
  assign n3689 = ( ~n629 & n3650 ) | ( ~n629 & n3685 ) | ( n3650 & n3685 ) ;
  assign n3690 = n153 | n300 ;
  assign n3691 = n629 | n3689 ;
  assign n3692 = n2664 | n3690 ;
  assign n3693 = n3687 | n3692 ;
  assign n3694 = ( n501 & ~n643 ) | ( n501 & n3693 ) | ( ~n643 & n3693 ) ;
  assign n3695 = n643 | n3694 ;
  assign n3696 = ( ~n2589 & n3675 ) | ( ~n2589 & n3695 ) | ( n3675 & n3695 ) ;
  assign n3697 = ~n3695 & n3696 ;
  assign n3698 = ( ~n961 & n1879 ) | ( ~n961 & n3697 ) | ( n1879 & n3697 ) ;
  assign n3699 = n276 | n290 ;
  assign n3700 = n3548 & ~n3695 ;
  assign n3701 = ~n1879 & n3698 ;
  assign n3702 = ~n3006 & n3700 ;
  assign n3703 = n1369 | n3699 ;
  assign n3704 = n2370 | n3699 ;
  assign n3705 = n3702 & ~n3703 ;
  assign n3706 = ( ~n713 & n1123 ) | ( ~n713 & n3701 ) | ( n1123 & n3701 ) ;
  assign n3707 = n283 | n546 ;
  assign n3708 = ~n1123 & n3706 ;
  assign n3709 = ( n2232 & ~n2666 ) | ( n2232 & n3708 ) | ( ~n2666 & n3708 ) ;
  assign n3710 = n3704 | n3707 ;
  assign n3711 = n3672 | n3710 ;
  assign n3712 = n886 | n2041 ;
  assign n3713 = n1135 | n2939 ;
  assign n3714 = n3712 | n3713 ;
  assign n3715 = n530 | n829 ;
  assign n3716 = n2895 | n3714 ;
  assign n3717 = n285 | n900 ;
  assign n3718 = n2669 | n3715 ;
  assign n3719 = n3717 | n3718 ;
  assign n3720 = n1777 | n3719 ;
  assign n3721 = n3195 | n3720 ;
  assign n3722 = n397 | n961 ;
  assign n3723 = n2973 | n3721 ;
  assign n3724 = n3664 | n3722 ;
  assign n3725 = n3391 | n3722 ;
  assign n3726 = n3586 | n3722 ;
  assign n3727 = n1466 | n3401 ;
  assign n3728 = n207 | n283 ;
  assign n3729 = n107 | n3029 ;
  assign n3730 = ~n3664 & n3665 ;
  assign n3731 = n823 | n3728 ;
  assign n3732 = n229 | n490 ;
  assign n3733 = n886 | n3732 ;
  assign n3734 = n95 | n145 ;
  assign n3735 = n3726 | n3733 ;
  assign n3736 = n3731 | n3733 ;
  assign n3737 = ~n425 & n3656 ;
  assign n3738 = n561 | n3731 ;
  assign n3739 = n3737 & ~n3738 ;
  assign n3740 = n290 | n342 ;
  assign n3741 = n2030 | n3734 ;
  assign n3742 = n3682 | n3740 ;
  assign n3743 = n3719 | n3741 ;
  assign n3744 = n536 | n3741 ;
  assign n3745 = n167 | n187 ;
  assign n3746 = n533 | n3745 ;
  assign n3747 = n321 | n2507 ;
  assign n3748 = n3746 | n3747 ;
  assign n3749 = n125 | n149 ;
  assign n3750 = n1622 | n3749 ;
  assign n3751 = n1821 | n3745 ;
  assign n3752 = ~n2695 & n3739 ;
  assign n3753 = ~n1395 & n3752 ;
  assign n3754 = ~n3751 & n3753 ;
  assign n3755 = n103 | n969 ;
  assign n3756 = n3744 | n3750 ;
  assign n3757 = n3740 | n3755 ;
  assign n3758 = n967 | n3729 ;
  assign n3759 = n3757 | n3758 ;
  assign n3760 = n1730 | n3759 ;
  assign n3761 = n3756 | n3760 ;
  assign n3762 = ( n1975 & ~n2266 ) | ( n1975 & n3761 ) | ( ~n2266 & n3761 ) ;
  assign n3763 = n2266 | n3762 ;
  assign n3764 = ( n352 & ~n520 ) | ( n352 & n3763 ) | ( ~n520 & n3763 ) ;
  assign n3765 = n520 | n3764 ;
  assign n3766 = ( n375 & ~n941 ) | ( n375 & n3765 ) | ( ~n941 & n3765 ) ;
  assign n3767 = n941 | n3766 ;
  assign n3768 = ( ~n89 & n172 ) | ( ~n89 & n3767 ) | ( n172 & n3767 ) ;
  assign n3769 = n89 | n3768 ;
  assign n3770 = ( ~n219 & n578 ) | ( ~n219 & n3769 ) | ( n578 & n3769 ) ;
  assign n3771 = n219 | n3770 ;
  assign n3772 = n1466 | n3771 ;
  assign n3773 = n3735 | n3772 ;
  assign n3774 = ( ~n1496 & n2565 ) | ( ~n1496 & n3773 ) | ( n2565 & n3773 ) ;
  assign n3775 = n2329 | n3200 ;
  assign n3776 = ( n373 & ~n602 ) | ( n373 & n3775 ) | ( ~n602 & n3775 ) ;
  assign n3777 = n3348 | n3513 ;
  assign n3778 = n255 | n532 ;
  assign n3779 = n397 | n3778 ;
  assign n3780 = n480 | n3779 ;
  assign n3781 = n1769 | n2670 ;
  assign n3782 = n285 | n3781 ;
  assign n3783 = n1059 | n3779 ;
  assign n3784 = n602 | n3776 ;
  assign n3785 = n284 | n1467 ;
  assign n3786 = n400 | n3593 ;
  assign n3787 = ( ~n547 & n683 ) | ( ~n547 & n3784 ) | ( n683 & n3784 ) ;
  assign n3788 = n547 | n3787 ;
  assign n3789 = ( n357 & ~n650 ) | ( n357 & n3788 ) | ( ~n650 & n3788 ) ;
  assign n3790 = n650 | n3789 ;
  assign n3791 = n3680 | n3785 ;
  assign n3792 = n3783 | n3786 ;
  assign n3793 = n872 | n3790 ;
  assign n3794 = n103 | n735 ;
  assign n3795 = n3358 | n3794 ;
  assign n3796 = n345 | n788 ;
  assign n3797 = n3792 | n3795 ;
  assign n3798 = n529 | n3796 ;
  assign n3799 = n3782 | n3798 ;
  assign n3800 = ( ~n220 & n955 ) | ( ~n220 & n3791 ) | ( n955 & n3791 ) ;
  assign n3801 = n3793 | n3798 ;
  assign n3802 = n3418 | n3801 ;
  assign n3803 = n220 | n3800 ;
  assign n3804 = n810 | n841 ;
  assign n3805 = n111 | n3804 ;
  assign n3806 = ( ~n1853 & n3699 ) | ( ~n1853 & n3802 ) | ( n3699 & n3802 ) ;
  assign n3807 = n1853 | n3806 ;
  assign n3808 = n957 | n2490 ;
  assign n3809 = n3805 | n3808 ;
  assign n3810 = n3145 | n3809 ;
  assign n3811 = ( ~n288 & n585 ) | ( ~n288 & n3810 ) | ( n585 & n3810 ) ;
  assign n3812 = n288 | n3811 ;
  assign n3813 = ( ~n461 & n589 ) | ( ~n461 & n3812 ) | ( n589 & n3812 ) ;
  assign n3814 = ( n139 & ~n653 ) | ( n139 & n3803 ) | ( ~n653 & n3803 ) ;
  assign n3815 = n653 | n3814 ;
  assign n3816 = n433 | n891 ;
  assign n3817 = n461 | n3813 ;
  assign n3818 = n3348 | n3816 ;
  assign n3819 = ( n146 & ~n400 ) | ( n146 & n3817 ) | ( ~n400 & n3817 ) ;
  assign n3820 = n3797 | n3819 ;
  assign n3821 = ( ~n439 & n1620 ) | ( ~n439 & n3820 ) | ( n1620 & n3820 ) ;
  assign n3822 = n2688 | n3816 ;
  assign n3823 = n439 | n3821 ;
  assign n3824 = ( ~n1902 & n2663 ) | ( ~n1902 & n3823 ) | ( n2663 & n3823 ) ;
  assign n3825 = n1902 | n3824 ;
  assign n3826 = ( n225 & ~n282 ) | ( n225 & n3825 ) | ( ~n282 & n3825 ) ;
  assign n3827 = n282 | n3826 ;
  assign n3828 = ( n173 & ~n631 ) | ( n173 & n3827 ) | ( ~n631 & n3827 ) ;
  assign n3829 = n631 | n3828 ;
  assign n3830 = ( ~n653 & n779 ) | ( ~n653 & n3829 ) | ( n779 & n3829 ) ;
  assign n3831 = n653 | n3830 ;
  assign n3832 = n204 | n3831 ;
  assign n3833 = ( n2119 & n3754 ) | ( n2119 & ~n3831 ) | ( n3754 & ~n3831 ) ;
  assign n3834 = n3816 | n3831 ;
  assign n3835 = n721 | n3815 ;
  assign n3836 = ~n2119 & n3833 ;
  assign n3837 = n3204 | n3834 ;
  assign n3838 = n3816 | n3835 ;
  assign n3839 = n2758 | n3838 ;
  assign n3840 = ( ~n677 & n1621 ) | ( ~n677 & n3839 ) | ( n1621 & n3839 ) ;
  assign n3841 = n3799 | n3837 ;
  assign n3842 = ( ~n1475 & n2293 ) | ( ~n1475 & n3841 ) | ( n2293 & n3841 ) ;
  assign n3843 = n1475 | n3842 ;
  assign n3844 = n149 | n721 ;
  assign n3845 = n583 & ~n3139 ;
  assign n3846 = ~n1382 & n3845 ;
  assign n3847 = n439 | n2942 ;
  assign n3848 = n2390 | n3844 ;
  assign n3849 = ~n318 & n3846 ;
  assign n3850 = ~n3848 & n3849 ;
  assign n3851 = ~n3847 & n3850 ;
  assign n3852 = n1496 | n3774 ;
  assign n3853 = n133 | n367 ;
  assign n3854 = ( n162 & ~n433 ) | ( n162 & n3851 ) | ( ~n433 & n3851 ) ;
  assign n3855 = n362 | n3853 ;
  assign n3856 = ~n162 & n3854 ;
  assign n3857 = ~n578 & n3856 ;
  assign n3858 = ( ~n1496 & n3094 ) | ( ~n1496 & n3857 ) | ( n3094 & n3857 ) ;
  assign n3859 = ~n3094 & n3858 ;
  assign n3860 = ~n1663 & n3557 ;
  assign n3861 = n211 | n248 ;
  assign n3862 = n3855 | n3861 ;
  assign n3863 = n282 | n719 ;
  assign n3864 = ~n1833 & n3857 ;
  assign n3865 = ~n2537 & n3864 ;
  assign n3866 = n177 | n714 ;
  assign n3867 = n3863 | n3866 ;
  assign n3868 = n1391 | n3848 ;
  assign n3869 = n1403 | n3862 ;
  assign n3870 = n419 | n3867 ;
  assign n3871 = n2170 | n3867 ;
  assign n3872 = n3869 | n3871 ;
  assign n3873 = n2879 | n3862 ;
  assign n3874 = n3725 | n3872 ;
  assign n3875 = ( ~n1035 & n1146 ) | ( ~n1035 & n3874 ) | ( n1146 & n3874 ) ;
  assign n3876 = n1035 | n3875 ;
  assign n3877 = n303 | n417 ;
  assign n3878 = n3868 | n3873 ;
  assign n3879 = ( ~n758 & n3876 ) | ( ~n758 & n3877 ) | ( n3876 & n3877 ) ;
  assign n3880 = n758 | n3879 ;
  assign n3881 = ( ~n167 & n532 ) | ( ~n167 & n3880 ) | ( n532 & n3880 ) ;
  assign n3882 = n188 | n631 ;
  assign n3883 = n3175 | n3882 ;
  assign n3884 = n530 | n2947 ;
  assign n3885 = n167 | n3881 ;
  assign n3886 = ( n378 & ~n476 ) | ( n378 & n3885 ) | ( ~n476 & n3885 ) ;
  assign n3887 = n476 | n3886 ;
  assign n3888 = n717 | n3887 ;
  assign n3889 = n1059 | n3888 ;
  assign n3890 = n3860 & ~n3889 ;
  assign n3891 = n144 | n846 ;
  assign n3892 = ~n1213 & n3890 ;
  assign n3893 = n788 | n3891 ;
  assign n3894 = n3615 | n3893 ;
  assign n3895 = n284 | n3883 ;
  assign n3896 = n3884 | n3895 ;
  assign n3897 = n3894 | n3896 ;
  assign n3898 = n1044 & ~n3897 ;
  assign n3899 = ( n123 & ~n1410 ) | ( n123 & n3898 ) | ( ~n1410 & n3898 ) ;
  assign n3900 = ~n123 & n3899 ;
  assign n3901 = ( n2911 & n3512 ) | ( n2911 & ~n3877 ) | ( n3512 & ~n3877 ) ;
  assign n3902 = n296 | n422 ;
  assign n3903 = n183 | n3512 ;
  assign n3904 = n3902 | n3903 ;
  assign n3905 = n2425 | n3904 ;
  assign n3906 = n2040 & ~n3905 ;
  assign n3907 = n420 | n503 ;
  assign n3908 = n965 | n2575 ;
  assign n3909 = n2333 | n3907 ;
  assign n3910 = n2326 | n3909 ;
  assign n3911 = n2879 | n3909 ;
  assign n3912 = n124 | n281 ;
  assign n3913 = n3908 | n3912 ;
  assign n3914 = n93 | n3487 ;
  assign n3915 = n3913 | n3914 ;
  assign n3916 = n381 | n580 ;
  assign n3917 = ( ~n953 & n955 ) | ( ~n953 & n3915 ) | ( n955 & n3915 ) ;
  assign n3918 = n953 | n3917 ;
  assign n3919 = n701 | n1318 ;
  assign n3920 = n3904 | n3918 ;
  assign n3921 = n3870 | n3920 ;
  assign n3922 = n124 | n555 ;
  assign n3923 = n2028 | n3922 ;
  assign n3924 = n3919 | n3923 ;
  assign n3925 = n3883 | n3924 ;
  assign n3926 = n2420 & ~n3925 ;
  assign n3927 = n433 | n546 ;
  assign n3928 = n3916 | n3927 ;
  assign n3929 = n1901 | n3928 ;
  assign n3930 = n3910 | n3929 ;
  assign n3931 = n83 | n288 ;
  assign n3932 = n756 | n758 ;
  assign n3933 = ( n94 & ~n461 ) | ( n94 & n3930 ) | ( ~n461 & n3930 ) ;
  assign n3934 = n2481 | n3931 ;
  assign n3935 = n461 | n3933 ;
  assign n3936 = ( n103 & ~n175 ) | ( n103 & n3935 ) | ( ~n175 & n3935 ) ;
  assign n3937 = n175 | n3936 ;
  assign n3938 = n600 | n3937 ;
  assign n3939 = n2179 | n3938 ;
  assign n3940 = n3934 | n3938 ;
  assign n3941 = n3921 | n3939 ;
  assign n3942 = n342 | n1712 ;
  assign n3943 = n3932 | n3942 ;
  assign n3944 = n3934 | n3943 ;
  assign n3945 = n3926 & ~n3944 ;
  assign n3946 = ( ~n655 & n2363 ) | ( ~n655 & n3945 ) | ( n2363 & n3945 ) ;
  assign n3947 = n3724 | n3940 ;
  assign n3948 = n2299 | n3947 ;
  assign n3949 = n3793 | n3943 ;
  assign n3950 = ~n2363 & n3946 ;
  assign n3951 = ( ~n655 & n2363 ) | ( ~n655 & n3941 ) | ( n2363 & n3941 ) ;
  assign n3952 = n107 | n601 ;
  assign n3953 = n1709 | n3952 ;
  assign n3954 = n3528 | n3953 ;
  assign n3955 = n350 | n3953 ;
  assign n3956 = n3805 | n3955 ;
  assign n3957 = n83 | n744 ;
  assign n3958 = n350 | n559 ;
  assign n3959 = n3957 | n3958 ;
  assign n3960 = n3233 | n3539 ;
  assign n3961 = n92 | n834 ;
  assign n3962 = n164 | n3961 ;
  assign n3963 = n3959 | n3960 ;
  assign n3964 = n1308 | n3877 ;
  assign n3965 = n1632 | n3964 ;
  assign n3966 = n3729 | n3962 ;
  assign n3967 = n3965 | n3966 ;
  assign n3968 = ( ~n522 & n747 ) | ( ~n522 & n3967 ) | ( n747 & n3967 ) ;
  assign n3969 = n522 | n3968 ;
  assign n3970 = ( ~n235 & n756 ) | ( ~n235 & n3969 ) | ( n756 & n3969 ) ;
  assign n3971 = n203 | n822 ;
  assign n3972 = n677 | n3840 ;
  assign n3973 = n235 | n3970 ;
  assign n3974 = n271 | n3973 ;
  assign n3975 = ( n3971 & n3972 ) | ( n3971 & ~n3974 ) | ( n3972 & ~n3974 ) ;
  assign n3976 = n3974 | n3975 ;
  assign n3977 = ( n1076 & ~n2939 ) | ( n1076 & n3976 ) | ( ~n2939 & n3976 ) ;
  assign n3978 = n133 | n303 ;
  assign n3979 = n101 | n846 ;
  assign n3980 = n81 | n293 ;
  assign n3981 = n3979 | n3980 ;
  assign n3982 = n444 | n580 ;
  assign n3983 = n3981 | n3982 ;
  assign n3984 = n2170 | n3442 ;
  assign n3985 = n3251 | n3984 ;
  assign n3986 = n294 | n302 ;
  assign n3987 = n503 | n3986 ;
  assign n3988 = n162 | n3978 ;
  assign n3989 = n3924 | n3983 ;
  assign n3990 = n3442 | n3988 ;
  assign n3991 = n2517 | n3983 ;
  assign n3992 = n1456 | n3987 ;
  assign n3993 = n2064 & ~n3992 ;
  assign n3994 = ~n3991 & n3993 ;
  assign n3995 = n283 | n422 ;
  assign n3996 = n3990 | n3995 ;
  assign n3997 = n2535 | n3996 ;
  assign n3998 = ( ~n3771 & n3994 ) | ( ~n3771 & n3996 ) | ( n3994 & n3996 ) ;
  assign n3999 = ~n3996 & n3998 ;
  assign n4000 = ~n2106 & n3999 ;
  assign n4001 = n3956 | n3997 ;
  assign n4002 = n1169 | n1250 ;
  assign n4003 = n100 | n731 ;
  assign n4004 = n447 | n4003 ;
  assign n4005 = n4002 | n4004 ;
  assign n4006 = n865 | n4004 ;
  assign n4007 = n415 | n502 ;
  assign n4008 = n2481 | n4007 ;
  assign n4009 = n789 | n4008 ;
  assign n4010 = n3988 | n4009 ;
  assign n4011 = n128 | n489 ;
  assign n4012 = n3148 & ~n4006 ;
  assign n4013 = n210 | n289 ;
  assign n4014 = n4011 | n4013 ;
  assign n4015 = n212 | n547 ;
  assign n4016 = n3522 | n4015 ;
  assign n4017 = n4005 | n4016 ;
  assign n4018 = n147 | n651 ;
  assign n4019 = ( n2541 & n4017 ) | ( n2541 & ~n4018 ) | ( n4017 & ~n4018 ) ;
  assign n4020 = n4018 | n4019 ;
  assign n4021 = ( ~n203 & n822 ) | ( ~n203 & n4020 ) | ( n822 & n4020 ) ;
  assign n4022 = n510 | n779 ;
  assign n4023 = n4014 | n4022 ;
  assign n4024 = n276 | n841 ;
  assign n4025 = ( ~n579 & n3369 ) | ( ~n579 & n3962 ) | ( n3369 & n3962 ) ;
  assign n4026 = n2293 | n4023 ;
  assign n4027 = n2836 | n4026 ;
  assign n4028 = n565 | n602 ;
  assign n4029 = n3575 | n4028 ;
  assign n4030 = n579 | n4025 ;
  assign n4031 = n565 | n4015 ;
  assign n4032 = n3521 | n4031 ;
  assign n4033 = n2086 | n4024 ;
  assign n4034 = n4029 | n4033 ;
  assign n4035 = n1738 | n3794 ;
  assign n4036 = n4032 | n4035 ;
  assign n4037 = n557 | n4018 ;
  assign n4038 = ( ~n547 & n644 ) | ( ~n547 & n4034 ) | ( n644 & n4034 ) ;
  assign n4039 = n547 | n4038 ;
  assign n4040 = ( n139 & ~n955 ) | ( n139 & n4039 ) | ( ~n955 & n4039 ) ;
  assign n4041 = n955 | n4040 ;
  assign n4042 = n1911 | n2405 ;
  assign n4043 = n3794 | n4041 ;
  assign n4044 = n4023 | n4043 ;
  assign n4045 = n229 | n969 ;
  assign n4046 = n4037 | n4045 ;
  assign n4047 = n4042 | n4046 ;
  assign n4048 = n3818 | n4044 ;
  assign n4049 = ( ~n307 & n579 ) | ( ~n307 & n4048 ) | ( n579 & n4048 ) ;
  assign n4050 = n307 | n4049 ;
  assign n4051 = n1243 | n4046 ;
  assign n4052 = ( n557 & ~n2481 ) | ( n557 & n4050 ) | ( ~n2481 & n4050 ) ;
  assign n4053 = n3911 | n4047 ;
  assign n4054 = n2481 | n4052 ;
  assign n4055 = ( ~n420 & n510 ) | ( ~n420 & n4036 ) | ( n510 & n4036 ) ;
  assign n4056 = n321 | n1299 ;
  assign n4057 = n420 | n4055 ;
  assign n4058 = n653 | n1312 ;
  assign n4059 = n650 | n4057 ;
  assign n4060 = n3987 | n4059 ;
  assign n4061 = n416 | n923 ;
  assign n4062 = n967 | n4061 ;
  assign n4063 = n3745 | n4058 ;
  assign n4064 = n3745 | n3877 ;
  assign n4065 = n4060 | n4064 ;
  assign n4066 = n1371 | n4062 ;
  assign n4067 = n3878 | n4066 ;
  assign n4068 = n125 | n427 ;
  assign n4069 = n827 | n4068 ;
  assign n4070 = n4062 | n4069 ;
  assign n4071 = n3091 | n4070 ;
  assign n4072 = n98 | n241 ;
  assign n4073 = ( n677 & n4001 ) | ( n677 & ~n4072 ) | ( n4001 & ~n4072 ) ;
  assign n4074 = n4072 | n4073 ;
  assign n4075 = ( n1318 & ~n1382 ) | ( n1318 & n4074 ) | ( ~n1382 & n4074 ) ;
  assign n4076 = n1382 | n4075 ;
  assign n4077 = ( ~n144 & n150 ) | ( ~n144 & n4076 ) | ( n150 & n4076 ) ;
  assign n4078 = n144 | n4077 ;
  assign n4079 = ( n415 & ~n941 ) | ( n415 & n4078 ) | ( ~n941 & n4078 ) ;
  assign n4080 = ( ~n271 & n3973 ) | ( ~n271 & n4067 ) | ( n3973 & n4067 ) ;
  assign n4081 = n941 | n4079 ;
  assign n4082 = n759 | n4081 ;
  assign n4083 = ( ~n759 & n2151 ) | ( ~n759 & n4081 ) | ( n2151 & n4081 ) ;
  assign n4084 = n759 | n4083 ;
  assign n4085 = ( n1818 & n4071 ) | ( n1818 & ~n4072 ) | ( n4071 & ~n4072 ) ;
  assign n4086 = n589 | n747 ;
  assign n4087 = ( n877 & ~n2664 ) | ( n877 & n4084 ) | ( ~n2664 & n4084 ) ;
  assign n4088 = n177 | n790 ;
  assign n4089 = n4086 | n4088 ;
  assign n4090 = n2712 | n4089 ;
  assign n4091 = n109 | n225 ;
  assign n4092 = n235 | n4091 ;
  assign n4093 = n4069 | n4092 ;
  assign n4094 = n2170 | n4092 ;
  assign n4095 = n4051 | n4094 ;
  assign n4096 = n4072 | n4085 ;
  assign n4097 = ( n2224 & n3172 ) | ( n2224 & ~n4096 ) | ( n3172 & ~n4096 ) ;
  assign n4098 = n2574 | n4093 ;
  assign n4099 = n4096 | n4097 ;
  assign n4100 = n894 | n4090 ;
  assign n4101 = n4095 | n4100 ;
  assign n4102 = ( n950 & ~n4082 ) | ( n950 & n4101 ) | ( ~n4082 & n4101 ) ;
  assign n4103 = ~n4101 & n4102 ;
  assign n4104 = n246 | n423 ;
  assign n4105 = n250 | n651 ;
  assign n4106 = n4104 | n4105 ;
  assign n4107 = n92 | n693 ;
  assign n4108 = n2947 | n4107 ;
  assign n4109 = n4106 | n4108 ;
  assign n4110 = n4086 | n4109 ;
  assign n4111 = n4065 | n4110 ;
  assign n4112 = n228 | n887 ;
  assign n4113 = n3654 | n4112 ;
  assign n4114 = ~n1410 & n2774 ;
  assign n4115 = n150 | n221 ;
  assign n4116 = n293 | n4115 ;
  assign n4117 = ( ~n1187 & n2670 ) | ( ~n1187 & n3538 ) | ( n2670 & n3538 ) ;
  assign n4118 = n982 | n4109 ;
  assign n4119 = n101 | n148 ;
  assign n4120 = n146 | n4119 ;
  assign n4121 = n2282 | n4118 ;
  assign n4122 = n3483 | n4120 ;
  assign n4123 = n4113 | n4122 ;
  assign n4124 = ( ~n647 & n713 ) | ( ~n647 & n4123 ) | ( n713 & n4123 ) ;
  assign n4125 = n647 | n4124 ;
  assign n4126 = n343 | n4125 ;
  assign n4127 = ( ~n1410 & n3294 ) | ( ~n1410 & n4126 ) | ( n3294 & n4126 ) ;
  assign n4128 = n1410 | n4127 ;
  assign n4129 = n87 | n89 ;
  assign n4130 = n203 | n4021 ;
  assign n4131 = n2369 | n4120 ;
  assign n4132 = n109 | n414 ;
  assign n4133 = n4129 | n4132 ;
  assign n4134 = n1310 | n4116 ;
  assign n4135 = ( n1307 & ~n1514 ) | ( n1307 & n4130 ) | ( ~n1514 & n4130 ) ;
  assign n4136 = n1514 | n4135 ;
  assign n4137 = n4133 | n4134 ;
  assign n4138 = ( n332 & ~n336 ) | ( n332 & n4136 ) | ( ~n336 & n4136 ) ;
  assign n4139 = n336 | n4138 ;
  assign n4140 = n124 | n4139 ;
  assign n4141 = n1187 | n4140 ;
  assign n4142 = n1838 | n4131 ;
  assign n4143 = n3927 | n4116 ;
  assign n4144 = n1299 | n4086 ;
  assign n4145 = n4126 | n4143 ;
  assign n4146 = n3730 & ~n4137 ;
  assign n4147 = ~n1001 & n4146 ;
  assign n4148 = ~n4141 & n4147 ;
  assign n4149 = ~n4107 & n4148 ;
  assign n4150 = ( ~n300 & n3916 ) | ( ~n300 & n4121 ) | ( n3916 & n4121 ) ;
  assign n4151 = n300 | n4150 ;
  assign n4152 = ( n103 & ~n128 ) | ( n103 & n4151 ) | ( ~n128 & n4151 ) ;
  assign n4153 = n2664 | n4087 ;
  assign n4154 = n128 | n4152 ;
  assign n4155 = ( ~n547 & n719 ) | ( ~n547 & n4154 ) | ( n719 & n4154 ) ;
  assign n4156 = n547 | n4155 ;
  assign n4157 = ( ~n210 & n969 ) | ( ~n210 & n4156 ) | ( n969 & n4156 ) ;
  assign n4158 = n210 | n4157 ;
  assign n4159 = n2821 | n4158 ;
  assign n4160 = n2769 | n4159 ;
  assign n4161 = ( n2718 & n3607 ) | ( n2718 & ~n4160 ) | ( n3607 & ~n4160 ) ;
  assign n4162 = n4160 | n4161 ;
  assign n4163 = ( n2664 & ~n3483 ) | ( n2664 & n4162 ) | ( ~n3483 & n4162 ) ;
  assign n4164 = n197 | n650 ;
  assign n4165 = n361 | n2230 ;
  assign n4166 = n4164 | n4165 ;
  assign n4167 = n1740 | n4024 ;
  assign n4168 = ~n3481 & n3739 ;
  assign n4169 = n1089 | n1309 ;
  assign n4170 = n4166 | n4167 ;
  assign n4171 = n3481 | n4169 ;
  assign n4172 = n489 | n501 ;
  assign n4173 = n3065 | n4024 ;
  assign n4174 = n2429 | n4024 ;
  assign n4175 = n1964 | n4174 ;
  assign n4176 = n289 | n644 ;
  assign n4177 = ( n3481 & n3807 ) | ( n3481 & ~n4172 ) | ( n3807 & ~n4172 ) ;
  assign n4178 = n1902 | n3893 ;
  assign n4179 = n2230 | n3481 ;
  assign n4180 = n143 | n2535 ;
  assign n4181 = ( n90 & ~n175 ) | ( n90 & n4170 ) | ( ~n175 & n4170 ) ;
  assign n4182 = n2718 | n4172 ;
  assign n4183 = n4176 | n4182 ;
  assign n4184 = n4178 | n4183 ;
  assign n4185 = n720 | n4172 ;
  assign n4186 = n4145 | n4185 ;
  assign n4187 = n4172 | n4177 ;
  assign n4188 = ( ~n2669 & n3963 ) | ( ~n2669 & n4186 ) | ( n3963 & n4186 ) ;
  assign n4189 = n2669 | n4188 ;
  assign n4190 = n82 | n241 ;
  assign n4191 = n3593 | n4190 ;
  assign n4192 = ( n143 & ~n2232 ) | ( n143 & n4187 ) | ( ~n2232 & n4187 ) ;
  assign n4193 = n4189 | n4190 ;
  assign n4194 = ( ~n169 & n173 ) | ( ~n169 & n4193 ) | ( n173 & n4193 ) ;
  assign n4195 = n169 | n4194 ;
  assign n4196 = ( ~n612 & n1333 ) | ( ~n612 & n4195 ) | ( n1333 & n4195 ) ;
  assign n4197 = n175 | n4181 ;
  assign n4198 = ( n351 & ~n862 ) | ( n351 & n4197 ) | ( ~n862 & n4197 ) ;
  assign n4199 = n862 | n4198 ;
  assign n4200 = n2660 | n4199 ;
  assign n4201 = n1456 | n4199 ;
  assign n4202 = n612 | n4196 ;
  assign n4203 = ( ~n210 & n973 ) | ( ~n210 & n4202 ) | ( n973 & n4202 ) ;
  assign n4204 = n210 | n4203 ;
  assign n4205 = n2821 | n4204 ;
  assign n4206 = n4180 | n4205 ;
  assign n4207 = n2903 | n4206 ;
  assign n4208 = n90 | n942 ;
  assign n4209 = n923 | n1145 ;
  assign n4210 = n646 | n4208 ;
  assign n4211 = n4191 | n4210 ;
  assign n4212 = n360 | n965 ;
  assign n4213 = n3483 | n4163 ;
  assign n4214 = ( ~n1174 & n4211 ) | ( ~n1174 & n4213 ) | ( n4211 & n4213 ) ;
  assign n4215 = n1174 | n4214 ;
  assign n4216 = n585 | n591 ;
  assign n4217 = n4212 | n4216 ;
  assign n4218 = n348 | n425 ;
  assign n4219 = ( n2246 & ~n2333 ) | ( n2246 & n3051 ) | ( ~n2333 & n3051 ) ;
  assign n4220 = n4209 | n4217 ;
  assign n4221 = n3336 | n4220 ;
  assign n4222 = n231 | n759 ;
  assign n4223 = n870 & ~n4222 ;
  assign n4224 = ( ~n4204 & n4221 ) | ( ~n4204 & n4223 ) | ( n4221 & n4223 ) ;
  assign n4225 = ~n4221 & n4224 ;
  assign n4226 = n97 | n224 ;
  assign n4227 = n4015 | n4226 ;
  assign n4228 = n660 | n4222 ;
  assign n4229 = n2232 | n4192 ;
  assign n4230 = n2333 | n4228 ;
  assign n4231 = n4171 | n4230 ;
  assign n4232 = n255 | n943 ;
  assign n4233 = ( n1184 & n4225 ) | ( n1184 & ~n4232 ) | ( n4225 & ~n4232 ) ;
  assign n4234 = ~n1184 & n4233 ;
  assign n4235 = ( ~n1125 & n2663 ) | ( ~n1125 & n4234 ) | ( n2663 & n4234 ) ;
  assign n4236 = ( ~n97 & n415 ) | ( ~n97 & n4231 ) | ( n415 & n4231 ) ;
  assign n4237 = ( ~n2266 & n4229 ) | ( ~n2266 & n4232 ) | ( n4229 & n4232 ) ;
  assign n4238 = n288 | n552 ;
  assign n4239 = ~n2663 & n4235 ;
  assign n4240 = ( n211 & ~n2351 ) | ( n211 & n4239 ) | ( ~n2351 & n4239 ) ;
  assign n4241 = n2266 | n4237 ;
  assign n4242 = n97 | n4236 ;
  assign n4243 = ( ~n224 & n1679 ) | ( ~n224 & n4241 ) | ( n1679 & n4241 ) ;
  assign n4244 = n224 | n4243 ;
  assign n4245 = ~n211 & n4240 ;
  assign n4246 = n963 | n4242 ;
  assign n4247 = n1512 | n4246 ;
  assign n4248 = n2613 | n4238 ;
  assign n4249 = n4218 | n4248 ;
  assign n4250 = n2264 | n4247 ;
  assign n4251 = ~n1997 & n4245 ;
  assign n4252 = n488 | n4249 ;
  assign n4253 = ( ~n677 & n3550 ) | ( ~n677 & n4232 ) | ( n3550 & n4232 ) ;
  assign n4254 = n3954 | n4252 ;
  assign n4255 = ~n4232 & n4253 ;
  assign n4256 = ( n285 & ~n345 ) | ( n285 & n4255 ) | ( ~n345 & n4255 ) ;
  assign n4257 = ( n3299 & ~n4246 ) | ( n3299 & n4254 ) | ( ~n4246 & n4254 ) ;
  assign n4258 = n4246 | n4257 ;
  assign n4259 = ~n285 & n4256 ;
  assign n4260 = ( n553 & ~n1246 ) | ( n553 & n3488 ) | ( ~n1246 & n3488 ) ;
  assign n4261 = n247 | n552 ;
  assign n4262 = n1246 | n4260 ;
  assign n4263 = ( ~n336 & n1056 ) | ( ~n336 & n4262 ) | ( n1056 & n4262 ) ;
  assign n4264 = n336 | n4263 ;
  assign n4265 = ( n95 & ~n823 ) | ( n95 & n4264 ) | ( ~n823 & n4264 ) ;
  assign n4266 = n1623 | n1914 ;
  assign n4267 = n3796 | n4261 ;
  assign n4268 = n823 | n4265 ;
  assign n4269 = n128 | n295 ;
  assign n4270 = ( n125 & ~n649 ) | ( n125 & n4268 ) | ( ~n649 & n4268 ) ;
  assign n4271 = n649 | n4270 ;
  assign n4272 = ( n221 & ~n348 ) | ( n221 & n4271 ) | ( ~n348 & n4271 ) ;
  assign n4273 = n348 | n4272 ;
  assign n4274 = ( ~n360 & n362 ) | ( ~n360 & n4273 ) | ( n362 & n4273 ) ;
  assign n4275 = n360 | n4274 ;
  assign n4276 = n360 | n2603 ;
  assign n4277 = n4269 | n4276 ;
  assign n4278 = n222 | n810 ;
  assign n4279 = n2593 | n4278 ;
  assign n4280 = n1914 | n4278 ;
  assign n4281 = n497 | n4278 ;
  assign n4282 = n4267 | n4281 ;
  assign n4283 = n823 | n2490 ;
  assign n4284 = n4277 | n4283 ;
  assign n4285 = n296 | n607 ;
  assign n4286 = n2490 | n4285 ;
  assign n4287 = ( ~n188 & n2755 ) | ( ~n188 & n4275 ) | ( n2755 & n4275 ) ;
  assign n4288 = n2606 | n4286 ;
  assign n4289 = ( ~n1417 & n3631 ) | ( ~n1417 & n3835 ) | ( n3631 & n3835 ) ;
  assign n4290 = n97 | n147 ;
  assign n4291 = n592 | n4290 ;
  assign n4292 = n4173 | n4291 ;
  assign n4293 = n1088 | n1391 ;
  assign n4294 = n4279 | n4292 ;
  assign n4295 = ( ~n188 & n4275 ) | ( ~n188 & n4294 ) | ( n4275 & n4294 ) ;
  assign n4296 = n611 | n4288 ;
  assign n4297 = n371 | n1764 ;
  assign n4298 = n4280 | n4297 ;
  assign n4299 = n1195 | n4298 ;
  assign n4300 = n4293 | n4299 ;
  assign n4301 = n1417 | n4289 ;
  assign n4302 = ( n611 & ~n1349 ) | ( n611 & n4301 ) | ( ~n1349 & n4301 ) ;
  assign n4303 = n3230 | n4296 ;
  assign n4304 = n3888 | n4298 ;
  assign n4305 = ( ~n1902 & n2446 ) | ( ~n1902 & n4303 ) | ( n2446 & n4303 ) ;
  assign n4306 = n1902 | n4305 ;
  assign n4307 = n433 | n489 ;
  assign n4308 = n188 | n4287 ;
  assign n4309 = ( ~n97 & n1679 ) | ( ~n97 & n4054 ) | ( n1679 & n4054 ) ;
  assign n4310 = n97 | n4309 ;
  assign n4311 = n1395 | n4307 ;
  assign n4312 = ( ~n165 & n220 ) | ( ~n165 & n4310 ) | ( n220 & n4310 ) ;
  assign n4313 = n2217 | n4311 ;
  assign n4314 = n165 | n4312 ;
  assign n4315 = ( n148 & ~n416 ) | ( n148 & n4314 ) | ( ~n416 & n4314 ) ;
  assign n4316 = n416 | n4315 ;
  assign n4317 = n3389 | n4313 ;
  assign n4318 = ( ~n2217 & n4308 ) | ( ~n2217 & n4316 ) | ( n4308 & n4316 ) ;
  assign n4319 = n188 | n4295 ;
  assign n4320 = ( ~n92 & n154 ) | ( ~n92 & n4317 ) | ( n154 & n4317 ) ;
  assign n4321 = n92 | n4320 ;
  assign n4322 = n735 | n810 ;
  assign n4323 = ( ~n116 & n960 ) | ( ~n116 & n4321 ) | ( n960 & n4321 ) ;
  assign n4324 = n116 | n4323 ;
  assign n4325 = ( n172 & ~n659 ) | ( n172 & n4324 ) | ( ~n659 & n4324 ) ;
  assign n4326 = ( n101 & ~n220 ) | ( n101 & n3350 ) | ( ~n220 & n3350 ) ;
  assign n4327 = n220 | n4326 ;
  assign n4328 = ( n583 & n829 ) | ( n583 & ~n4327 ) | ( n829 & ~n4327 ) ;
  assign n4329 = n2217 | n4318 ;
  assign n4330 = ~n829 & n4328 ;
  assign n4331 = n694 | n823 ;
  assign n4332 = n4322 | n4331 ;
  assign n4333 = n659 | n4325 ;
  assign n4334 = ( n2417 & ~n4018 ) | ( n2417 & n4332 ) | ( ~n4018 & n4332 ) ;
  assign n4335 = n4018 | n4334 ;
  assign n4336 = ( n796 & ~n2549 ) | ( n796 & n4335 ) | ( ~n2549 & n4335 ) ;
  assign n4337 = ( ~n580 & n655 ) | ( ~n580 & n4333 ) | ( n655 & n4333 ) ;
  assign n4338 = n580 | n4337 ;
  assign n4339 = ( ~n4319 & n4330 ) | ( ~n4319 & n4338 ) | ( n4330 & n4338 ) ;
  assign n4340 = n2549 | n4336 ;
  assign n4341 = ( ~n100 & n229 ) | ( ~n100 & n4340 ) | ( n229 & n4340 ) ;
  assign n4342 = n100 | n4341 ;
  assign n4343 = n849 | n4342 ;
  assign n4344 = ( n1965 & n4338 ) | ( n1965 & ~n4343 ) | ( n4338 & ~n4343 ) ;
  assign n4345 = n4343 | n4344 ;
  assign n4346 = ( ~n1781 & n3846 ) | ( ~n1781 & n4345 ) | ( n3846 & n4345 ) ;
  assign n4347 = n3607 | n4338 ;
  assign n4348 = ( ~n849 & n1786 ) | ( ~n849 & n4342 ) | ( n1786 & n4342 ) ;
  assign n4349 = ~n4338 & n4339 ;
  assign n4350 = ~n3759 & n4349 ;
  assign n4351 = n849 | n4348 ;
  assign n4352 = ( ~n3749 & n4204 ) | ( ~n3749 & n4351 ) | ( n4204 & n4351 ) ;
  assign n4353 = ~n4345 & n4346 ;
  assign n4354 = n88 | n248 ;
  assign n4355 = n172 | n222 ;
  assign n4356 = n1460 | n4355 ;
  assign n4357 = n4354 | n4356 ;
  assign n4358 = ( n351 & ~n963 ) | ( n351 & n4357 ) | ( ~n963 & n4357 ) ;
  assign n4359 = n426 | n941 ;
  assign n4360 = n4285 | n4359 ;
  assign n4361 = ( n491 & ~n3396 ) | ( n491 & n3749 ) | ( ~n3396 & n3749 ) ;
  assign n4362 = n3396 | n4361 ;
  assign n4363 = ( n1230 & ~n2028 ) | ( n1230 & n4362 ) | ( ~n2028 & n4362 ) ;
  assign n4364 = n2028 | n4363 ;
  assign n4365 = ( ~n133 & n3266 ) | ( ~n133 & n4364 ) | ( n3266 & n4364 ) ;
  assign n4366 = n133 | n4365 ;
  assign n4367 = ( ~n534 & n612 ) | ( ~n534 & n4366 ) | ( n612 & n4366 ) ;
  assign n4368 = n785 | n3534 ;
  assign n4369 = n534 | n4367 ;
  assign n4370 = ( n111 & ~n735 ) | ( n111 & n4369 ) | ( ~n735 & n4369 ) ;
  assign n4371 = n735 | n4370 ;
  assign n4372 = n963 | n4358 ;
  assign n4373 = n520 | n790 ;
  assign n4374 = ( ~n1855 & n4368 ) | ( ~n1855 & n4371 ) | ( n4368 & n4371 ) ;
  assign n4375 = n146 | n4373 ;
  assign n4376 = n4360 | n4371 ;
  assign n4377 = n3210 | n4376 ;
  assign n4378 = n4372 | n4375 ;
  assign n4379 = n4175 | n4378 ;
  assign n4380 = ( n2329 & ~n2663 ) | ( n2329 & n4379 ) | ( ~n2663 & n4379 ) ;
  assign n4381 = ~n1001 & n4330 ;
  assign n4382 = n2663 | n4380 ;
  assign n4383 = ( ~n293 & n336 ) | ( ~n293 & n4382 ) | ( n336 & n4382 ) ;
  assign n4384 = n961 | n3688 ;
  assign n4385 = n293 | n4383 ;
  assign n4386 = ( ~n211 & n348 ) | ( ~n211 & n4385 ) | ( n348 & n4385 ) ;
  assign n4387 = n211 | n4386 ;
  assign n4388 = ( n425 & ~n605 ) | ( n425 & n4387 ) | ( ~n605 & n4387 ) ;
  assign n4389 = n605 | n4388 ;
  assign n4390 = n400 | n4389 ;
  assign n4391 = n275 | n4390 ;
  assign n4392 = n4381 & ~n4391 ;
  assign n4393 = ~n3736 & n4392 ;
  assign n4394 = ( ~n1855 & n2830 ) | ( ~n1855 & n4393 ) | ( n2830 & n4393 ) ;
  assign n4395 = ( ~n2128 & n4384 ) | ( ~n2128 & n4390 ) | ( n4384 & n4390 ) ;
  assign n4396 = n1855 | n3429 ;
  assign n4397 = ~n2830 & n4394 ;
  assign n4398 = n1855 | n4374 ;
  assign n4399 = n2128 | n4395 ;
  assign n4400 = ( ~n3916 & n4059 ) | ( ~n3916 & n4399 ) | ( n4059 & n4399 ) ;
  assign n4401 = n659 | n735 ;
  assign n4402 = n754 | n4401 ;
  assign n4403 = n4249 | n4402 ;
  assign n4404 = n2177 | n4360 ;
  assign n4405 = n2429 | n4402 ;
  assign n4406 = n4250 | n4405 ;
  assign n4407 = n998 | n1818 ;
  assign n4408 = n4404 | n4407 ;
  assign n4409 = n300 | n381 ;
  assign n4410 = n961 | n4409 ;
  assign n4411 = n4347 | n4410 ;
  assign n4412 = n1740 | n4410 ;
  assign n4413 = n4408 | n4412 ;
  assign n4414 = n713 | n788 ;
  assign n4415 = ( n2909 & n4406 ) | ( n2909 & ~n4414 ) | ( n4406 & ~n4414 ) ;
  assign n4416 = n4414 | n4415 ;
  assign n4417 = ( ~n165 & n1088 ) | ( ~n165 & n4416 ) | ( n1088 & n4416 ) ;
  assign n4418 = n165 | n4417 ;
  assign n4419 = ( ~n207 & n293 ) | ( ~n207 & n4418 ) | ( n293 & n4418 ) ;
  assign n4420 = n207 | n4419 ;
  assign n4421 = ( n56 & ~n1340 ) | ( n56 & n4420 ) | ( ~n1340 & n4420 ) ;
  assign n4422 = ( ~n100 & n552 ) | ( ~n100 & n4098 ) | ( n552 & n4098 ) ;
  assign n4423 = n100 | n4422 ;
  assign n4424 = n3949 | n4411 ;
  assign n4425 = ( ~n1251 & n3691 ) | ( ~n1251 & n4421 ) | ( n3691 & n4421 ) ;
  assign n4426 = ( n203 & ~n872 ) | ( n203 & n4423 ) | ( ~n872 & n4423 ) ;
  assign n4427 = n872 | n4426 ;
  assign n4428 = n444 | n4427 ;
  assign n4429 = n202 | n4428 ;
  assign n4430 = n534 | n953 ;
  assign n4431 = ( n2778 & ~n4072 ) | ( n2778 & n4421 ) | ( ~n4072 & n4421 ) ;
  assign n4432 = n4072 | n4431 ;
  assign n4433 = ( n1745 & ~n3491 ) | ( n1745 & n4432 ) | ( ~n3491 & n4432 ) ;
  assign n4434 = n3491 | n4433 ;
  assign n4435 = ( ~n796 & n2908 ) | ( ~n796 & n4434 ) | ( n2908 & n4434 ) ;
  assign n4436 = n332 | n823 ;
  assign n4437 = n4430 | n4436 ;
  assign n4438 = n4421 | n4437 ;
  assign n4439 = ~n2613 & n3846 ;
  assign n4440 = ~n4438 & n4439 ;
  assign n4441 = ~n4304 & n4440 ;
  assign n4442 = ~n4428 & n4441 ;
  assign n4443 = ~n1094 & n4442 ;
  assign n4444 = n585 | n631 ;
  assign n4445 = n967 | n4444 ;
  assign n4446 = n2617 | n4445 ;
  assign n4447 = n318 | n715 ;
  assign n4448 = n1193 | n3927 ;
  assign n4449 = n1193 | n3278 ;
  assign n4450 = n4446 | n4449 ;
  assign n4451 = n3780 | n4450 ;
  assign n4452 = n655 | n778 ;
  assign n4453 = ( ~n1630 & n3663 ) | ( ~n1630 & n4452 ) | ( n3663 & n4452 ) ;
  assign n4454 = n1630 | n4453 ;
  assign n4455 = ( n303 & ~n2939 ) | ( n303 & n4454 ) | ( ~n2939 & n4454 ) ;
  assign n4456 = n2939 | n4455 ;
  assign n4457 = ( n648 & ~n786 ) | ( n648 & n4456 ) | ( ~n786 & n4456 ) ;
  assign n4458 = n2549 | n3491 ;
  assign n4459 = n4447 | n4458 ;
  assign n4460 = n1859 | n4452 ;
  assign n4461 = n1251 | n4425 ;
  assign n4462 = ( ~n180 & n213 ) | ( ~n180 & n4451 ) | ( n213 & n4451 ) ;
  assign n4463 = n180 | n4462 ;
  assign n4464 = ( ~n82 & n207 ) | ( ~n82 & n4463 ) | ( n207 & n4463 ) ;
  assign n4465 = n82 | n4464 ;
  assign n4466 = ( n502 & ~n960 ) | ( n502 & n4465 ) | ( ~n960 & n4465 ) ;
  assign n4467 = n960 | n4466 ;
  assign n4468 = ( n583 & n754 ) | ( n583 & ~n4467 ) | ( n754 & ~n4467 ) ;
  assign n4469 = ~n754 & n4468 ;
  assign n4470 = ( n245 & ~n645 ) | ( n245 & n4469 ) | ( ~n645 & n4469 ) ;
  assign n4471 = ( ~n180 & n4284 ) | ( ~n180 & n4461 ) | ( n4284 & n4461 ) ;
  assign n4472 = ( ~n351 & n961 ) | ( ~n351 & n4459 ) | ( n961 & n4459 ) ;
  assign n4473 = ~n245 & n4470 ;
  assign n4474 = ~n1003 & n4473 ;
  assign n4475 = n3671 | n4472 ;
  assign n4476 = ( n4316 & n4473 ) | ( n4316 & ~n4475 ) | ( n4473 & ~n4475 ) ;
  assign n4477 = ~n4316 & n4476 ;
  assign n4478 = n341 | n887 ;
  assign n4479 = n4460 | n4478 ;
  assign n4480 = n2669 | n2681 ;
  assign n4481 = n4479 | n4480 ;
  assign n4482 = ( ~n612 & n756 ) | ( ~n612 & n4481 ) | ( n756 & n4481 ) ;
  assign n4483 = n612 | n4482 ;
  assign n4484 = ( n717 & ~n953 ) | ( n717 & n4483 ) | ( ~n953 & n4483 ) ;
  assign n4485 = n953 | n4484 ;
  assign n4486 = n1922 | n4414 ;
  assign n4487 = n372 | n4485 ;
  assign n4488 = ( ~n1417 & n4477 ) | ( ~n1417 & n4487 ) | ( n4477 & n4487 ) ;
  assign n4489 = n4284 | n4487 ;
  assign n4490 = ~n4487 & n4488 ;
  assign n4491 = n1159 | n2994 ;
  assign n4492 = n4486 | n4491 ;
  assign n4493 = ( ~n1514 & n2413 ) | ( ~n1514 & n3551 ) | ( n2413 & n3551 ) ;
  assign n4494 = n4489 | n4492 ;
  assign n4495 = n351 | n4472 ;
  assign n4496 = ( ~n1125 & n2324 ) | ( ~n1125 & n4494 ) | ( n2324 & n4494 ) ;
  assign n4497 = n1125 | n4496 ;
  assign n4498 = ( ~n153 & n302 ) | ( ~n153 & n4497 ) | ( n302 & n4497 ) ;
  assign n4499 = n153 | n4498 ;
  assign n4500 = n165 | n281 ;
  assign n4501 = ( ~n94 & n352 ) | ( ~n94 & n4499 ) | ( n352 & n4499 ) ;
  assign n4502 = n375 | n448 ;
  assign n4503 = n94 | n4501 ;
  assign n4504 = ( n89 & ~n546 ) | ( n89 & n4503 ) | ( ~n546 & n4503 ) ;
  assign n4505 = n1315 | n4500 ;
  assign n4506 = n546 | n4504 ;
  assign n4507 = n4502 | n4506 ;
  assign n4508 = n1959 | n4507 ;
  assign n4509 = n4474 & ~n4508 ;
  assign n4510 = ~n3989 & n4509 ;
  assign n4511 = ~n4041 & n4510 ;
  assign n4512 = ~n1136 & n4511 ;
  assign n4513 = n1460 | n4507 ;
  assign n4514 = ( ~n1349 & n1744 ) | ( ~n1349 & n4506 ) | ( n1744 & n4506 ) ;
  assign n4515 = ~n4506 & n4514 ;
  assign n4516 = ( n1514 & ~n4018 ) | ( n1514 & n4512 ) | ( ~n4018 & n4512 ) ;
  assign n4517 = n4505 | n4513 ;
  assign n4518 = n3777 | n4517 ;
  assign n4519 = ( ~n4140 & n4495 ) | ( ~n4140 & n4518 ) | ( n4495 & n4518 ) ;
  assign n4520 = n4140 | n4519 ;
  assign n4521 = ~n1514 & n4516 ;
  assign n4522 = ( n424 & ~n998 ) | ( n424 & n4521 ) | ( ~n998 & n4521 ) ;
  assign n4523 = n3036 & ~n4222 ;
  assign n4524 = n1384 | n1403 ;
  assign n4525 = n271 | n4080 ;
  assign n4526 = ( ~n225 & n4452 ) | ( ~n225 & n4525 ) | ( n4452 & n4525 ) ;
  assign n4527 = n225 | n4526 ;
  assign n4528 = ( ~n2266 & n4111 ) | ( ~n2266 & n4452 ) | ( n4111 & n4452 ) ;
  assign n4529 = n2266 | n4528 ;
  assign n4530 = ( ~n97 & n1367 ) | ( ~n97 & n4529 ) | ( n1367 & n4529 ) ;
  assign n4531 = n97 | n4530 ;
  assign n4532 = ( n583 & n1333 ) | ( n583 & ~n4527 ) | ( n1333 & ~n4527 ) ;
  assign n4533 = ~n1333 & n4532 ;
  assign n4534 = ~n945 & n4533 ;
  assign n4535 = ~n3181 & n4534 ;
  assign n4536 = n651 | n3482 ;
  assign n4537 = ( ~n2098 & n3916 ) | ( ~n2098 & n4536 ) | ( n3916 & n4536 ) ;
  assign n4538 = ~n95 & n4534 ;
  assign n4539 = ( n1738 & ~n3916 ) | ( n1738 & n4535 ) | ( ~n3916 & n4535 ) ;
  assign n4540 = n3916 | n4400 ;
  assign n4541 = ~n1920 & n4538 ;
  assign n4542 = ~n4524 & n4541 ;
  assign n4543 = n565 | n2613 ;
  assign n4544 = n81 | n375 ;
  assign n4545 = n942 | n4544 ;
  assign n4546 = n4543 | n4545 ;
  assign n4547 = n1764 | n4222 ;
  assign n4548 = n3749 | n4222 ;
  assign n4549 = n4546 | n4548 ;
  assign n4550 = n148 | n717 ;
  assign n4551 = n1251 | n4545 ;
  assign n4552 = ( ~n97 & n943 ) | ( ~n97 & n4549 ) | ( n943 & n4549 ) ;
  assign n4553 = n731 | n4550 ;
  assign n4554 = n97 | n4552 ;
  assign n4555 = n203 | n591 ;
  assign n4556 = ( n4053 & n4372 ) | ( n4053 & ~n4555 ) | ( n4372 & ~n4555 ) ;
  assign n4557 = n351 | n832 ;
  assign n4558 = n4553 | n4557 ;
  assign n4559 = n1467 | n2028 ;
  assign n4560 = n3365 | n4559 ;
  assign n4561 = ~n2413 & n4493 ;
  assign n4562 = n4551 | n4558 ;
  assign n4563 = n2477 | n2681 ;
  assign n4564 = n555 | n2551 ;
  assign n4565 = n796 | n4564 ;
  assign n4566 = ( n248 & ~n608 ) | ( n248 & n4554 ) | ( ~n608 & n4554 ) ;
  assign n4567 = n608 | n4566 ;
  assign n4568 = n343 | n4567 ;
  assign n4569 = n2720 | n4562 ;
  assign n4570 = n747 | n834 ;
  assign n4571 = n2477 | n4558 ;
  assign n4572 = n713 | n4570 ;
  assign n4573 = n2650 | n4572 ;
  assign n4574 = n2447 | n4573 ;
  assign n4575 = n672 | n4565 ;
  assign n4576 = n4560 | n4571 ;
  assign n4577 = n3186 | n4574 ;
  assign n4578 = ( ~n1195 & n2367 ) | ( ~n1195 & n4577 ) | ( n2367 & n4577 ) ;
  assign n4579 = n4565 | n4568 ;
  assign n4580 = n2956 & ~n4579 ;
  assign n4581 = ~n4577 & n4578 ;
  assign n4582 = ( n1833 & ~n3385 ) | ( n1833 & n4581 ) | ( ~n3385 & n4581 ) ;
  assign n4583 = ~n1833 & n4582 ;
  assign n4584 = n2866 & ~n4568 ;
  assign n4585 = ( n2413 & ~n4555 ) | ( n2413 & n4583 ) | ( ~n4555 & n4583 ) ;
  assign n4586 = ~n784 & n4580 ;
  assign n4587 = ~n2413 & n4586 ;
  assign n4588 = ~n2413 & n4585 ;
  assign n4589 = n122 | n1349 ;
  assign n4590 = n553 | n757 ;
  assign n4591 = n4589 | n4590 ;
  assign n4592 = n4547 | n4591 ;
  assign n4593 = n107 | n287 ;
  assign n4594 = n175 | n827 ;
  assign n4595 = ( ~n1248 & n1709 ) | ( ~n1248 & n4584 ) | ( n1709 & n4584 ) ;
  assign n4596 = n343 | n4593 ;
  assign n4597 = n553 | n4594 ;
  assign n4598 = n4596 | n4597 ;
  assign n4599 = n2126 | n4598 ;
  assign n4600 = n1113 | n4598 ;
  assign n4601 = n887 | n4228 ;
  assign n4602 = n4599 | n4601 ;
  assign n4603 = n3410 | n4602 ;
  assign n4604 = n228 | n520 ;
  assign n4605 = n180 | n476 ;
  assign n4606 = n4604 | n4605 ;
  assign n4607 = n211 | n887 ;
  assign n4608 = n2869 & ~n4600 ;
  assign n4609 = n318 | n341 ;
  assign n4610 = n646 | n2095 ;
  assign n4611 = n646 | n4606 ;
  assign n4612 = n4596 | n4611 ;
  assign n4613 = n229 | n448 ;
  assign n4614 = n4607 | n4613 ;
  assign n4615 = n4448 | n4614 ;
  assign n4616 = n271 | n4615 ;
  assign n4617 = n4555 | n4616 ;
  assign n4618 = n336 | n759 ;
  assign n4619 = n3749 | n4616 ;
  assign n4620 = ( n225 & ~n503 ) | ( n225 & n4576 ) | ( ~n503 & n4576 ) ;
  assign n4621 = n503 | n4620 ;
  assign n4622 = n3749 | n4352 ;
  assign n4623 = n303 | n410 ;
  assign n4624 = ( ~n210 & n647 ) | ( ~n210 & n4621 ) | ( n647 & n4621 ) ;
  assign n4625 = n210 | n4624 ;
  assign n4626 = n4609 | n4623 ;
  assign n4627 = n4618 | n4626 ;
  assign n4628 = n2125 | n4627 ;
  assign n4629 = n3669 | n4628 ;
  assign n4630 = n2878 | n4629 ;
  assign n4631 = ( ~n428 & n1620 ) | ( ~n428 & n4630 ) | ( n1620 & n4630 ) ;
  assign n4632 = ( n203 & ~n414 ) | ( n203 & n4625 ) | ( ~n414 & n4625 ) ;
  assign n4633 = n428 | n4631 ;
  assign n4634 = n4377 | n4617 ;
  assign n4635 = n414 | n4632 ;
  assign n4636 = n231 | n4635 ;
  assign n4637 = ( ~n4018 & n4633 ) | ( ~n4018 & n4636 ) | ( n4633 & n4636 ) ;
  assign n4638 = n4018 | n4637 ;
  assign n4639 = ( n502 & ~n916 ) | ( n502 & n4638 ) | ( ~n916 & n4638 ) ;
  assign n4640 = n916 | n4639 ;
  assign n4641 = ( ~n866 & n4608 ) | ( ~n866 & n4640 ) | ( n4608 & n4640 ) ;
  assign n4642 = ~n4640 & n4641 ;
  assign n4643 = n548 | n4606 ;
  assign n4644 = ~n2670 & n4117 ;
  assign n4645 = ~n1709 & n4595 ;
  assign n4646 = ( n1709 & ~n1833 ) | ( n1709 & n4642 ) | ( ~n1833 & n4642 ) ;
  assign n4647 = ~n1709 & n4646 ;
  assign n4648 = n1920 | n4640 ;
  assign n4649 = ( ~n373 & n2670 ) | ( ~n373 & n4647 ) | ( n2670 & n4647 ) ;
  assign n4650 = ~n2670 & n4649 ;
  assign n4651 = n4619 | n4648 ;
  assign n4652 = n547 | n659 ;
  assign n4653 = n3742 | n4652 ;
  assign n4654 = n144 | n756 ;
  assign n4655 = ( n561 & ~n846 ) | ( n561 & n3352 ) | ( ~n846 & n3352 ) ;
  assign n4656 = n846 | n4655 ;
  assign n4657 = ( n235 & ~n723 ) | ( n235 & n4656 ) | ( ~n723 & n4656 ) ;
  assign n4658 = n723 | n4657 ;
  assign n4659 = ( ~n476 & n489 ) | ( ~n476 & n4658 ) | ( n489 & n4658 ) ;
  assign n4660 = n476 | n4659 ;
  assign n4661 = ( n2509 & n4653 ) | ( n2509 & ~n4660 ) | ( n4653 & ~n4660 ) ;
  assign n4662 = n4660 | n4661 ;
  assign n4663 = n4636 | n4662 ;
  assign n4664 = n81 | n721 ;
  assign n4665 = n2551 | n4664 ;
  assign n4666 = n4610 | n4665 ;
  assign n4667 = n3221 | n4666 ;
  assign n4668 = n203 | n747 ;
  assign n4669 = n150 | n1125 ;
  assign n4670 = n4668 | n4669 ;
  assign n4671 = n2575 | n4654 ;
  assign n4672 = n4217 | n4671 ;
  assign n4673 = n1398 | n1992 ;
  assign n4674 = n4672 | n4673 ;
  assign n4675 = ~n2300 & n2367 ;
  assign n4676 = ( n565 & ~n1738 ) | ( n565 & n4674 ) | ( ~n1738 & n4674 ) ;
  assign n4677 = n4643 | n4670 ;
  assign n4678 = n1738 | n4676 ;
  assign n4679 = ( ~n286 & n1520 ) | ( ~n286 & n4678 ) | ( n1520 & n4678 ) ;
  assign n4680 = n286 | n4679 ;
  assign n4681 = n96 | n2300 ;
  assign n4682 = n3859 & ~n4653 ;
  assign n4683 = n1777 | n1846 ;
  assign n4684 = ( n1846 & n4072 ) | ( n1846 & ~n4667 ) | ( n4072 & ~n4667 ) ;
  assign n4685 = n468 | n1777 ;
  assign n4686 = ( n220 & ~n281 ) | ( n220 & n4680 ) | ( ~n281 & n4680 ) ;
  assign n4687 = n281 | n4686 ;
  assign n4688 = n4667 | n4684 ;
  assign n4689 = ( ~n414 & n683 ) | ( ~n414 & n4687 ) | ( n683 & n4687 ) ;
  assign n4690 = n172 | n960 ;
  assign n4691 = n414 | n4689 ;
  assign n4692 = n4685 | n4690 ;
  assign n4693 = n422 | n2657 ;
  assign n4694 = n231 | n4691 ;
  assign n4695 = n1574 | n2811 ;
  assign n4696 = n2367 & ~n4695 ;
  assign n4697 = ( ~n1303 & n4694 ) | ( ~n1303 & n4696 ) | ( n4694 & n4696 ) ;
  assign n4698 = ~n4694 & n4697 ;
  assign n4699 = ( n1230 & ~n2613 ) | ( n1230 & n4698 ) | ( ~n2613 & n4698 ) ;
  assign n4700 = ( n1230 & ~n1246 ) | ( n1230 & n4663 ) | ( ~n1246 & n4663 ) ;
  assign n4701 = ~n1230 & n4699 ;
  assign n4702 = ~n4693 & n4701 ;
  assign n4703 = ( ~n141 & n4207 ) | ( ~n141 & n4694 ) | ( n4207 & n4694 ) ;
  assign n4704 = n141 | n4703 ;
  assign n4705 = n4681 | n4692 ;
  assign n4706 = ~n2378 & n4702 ;
  assign n4707 = n4403 | n4677 ;
  assign n4708 = ( n3256 & n3483 ) | ( n3256 & ~n4688 ) | ( n3483 & ~n4688 ) ;
  assign n4709 = ( ~n281 & n295 ) | ( ~n281 & n2886 ) | ( n295 & n2886 ) ;
  assign n4710 = n4688 | n4708 ;
  assign n4711 = ( n2324 & ~n2939 ) | ( n2324 & n4645 ) | ( ~n2939 & n4645 ) ;
  assign n4712 = ( ~n1095 & n2460 ) | ( ~n1095 & n3491 ) | ( n2460 & n3491 ) ;
  assign n4713 = n1095 | n4712 ;
  assign n4714 = ( n2551 & ~n3175 ) | ( n2551 & n4713 ) | ( ~n3175 & n4713 ) ;
  assign n4715 = n3175 | n4714 ;
  assign n4716 = ( n165 & ~n420 ) | ( n165 & n4715 ) | ( ~n420 & n4715 ) ;
  assign n4717 = n420 | n4716 ;
  assign n4718 = ( ~n372 & n4397 ) | ( ~n372 & n4717 ) | ( n4397 & n4717 ) ;
  assign n4719 = ~n4717 & n4718 ;
  assign n4720 = ( ~n161 & n3113 ) | ( ~n161 & n4719 ) | ( n3113 & n4719 ) ;
  assign n4721 = ~n3113 & n4720 ;
  assign n4722 = n101 | n643 ;
  assign n4723 = n2937 | n3498 ;
  assign n4724 = ( n528 & ~n2611 ) | ( n528 & n4723 ) | ( ~n2611 & n4723 ) ;
  assign n4725 = n608 | n4705 ;
  assign n4726 = ( n1001 & ~n1144 ) | ( n1001 & n2751 ) | ( ~n1144 & n2751 ) ;
  assign n4727 = ( ~n2098 & n4710 ) | ( ~n2098 & n4725 ) | ( n4710 & n4725 ) ;
  assign n4728 = ( ~n372 & n4634 ) | ( ~n372 & n4717 ) | ( n4634 & n4717 ) ;
  assign n4729 = ~n2324 & n4711 ;
  assign n4730 = n372 | n4728 ;
  assign n4731 = ( ~n213 & n528 ) | ( ~n213 & n4730 ) | ( n528 & n4730 ) ;
  assign n4732 = n304 | n1333 ;
  assign n4733 = n4722 | n4732 ;
  assign n4734 = n84 | n2575 ;
  assign n4735 = n2575 | n4500 ;
  assign n4736 = n4733 | n4734 ;
  assign n4737 = n206 | n872 ;
  assign n4738 = n3782 | n4736 ;
  assign n4739 = n3083 | n4738 ;
  assign n4740 = n3303 | n4737 ;
  assign n4741 = n2476 | n4332 ;
  assign n4742 = n4429 | n4735 ;
  assign n4743 = n144 | n345 ;
  assign n4744 = ( ~n4725 & n4739 ) | ( ~n4725 & n4743 ) | ( n4739 & n4743 ) ;
  assign n4745 = n4725 | n4744 ;
  assign n4746 = ( ~n306 & n1307 ) | ( ~n306 & n4745 ) | ( n1307 & n4745 ) ;
  assign n4747 = n306 | n4746 ;
  assign n4748 = ( ~n149 & n683 ) | ( ~n149 & n4747 ) | ( n683 & n4747 ) ;
  assign n4749 = n149 | n4748 ;
  assign n4750 = n1144 | n4726 ;
  assign n4751 = n4740 | n4749 ;
  assign n4752 = n714 | n4749 ;
  assign n4753 = ( ~n1035 & n4750 ) | ( ~n1035 & n4752 ) | ( n4750 & n4752 ) ;
  assign n4754 = n2530 | n4751 ;
  assign n4755 = ( ~n4211 & n4741 ) | ( ~n4211 & n4754 ) | ( n4741 & n4754 ) ;
  assign n4756 = n4211 | n4755 ;
  assign n4757 = ( ~n372 & n4717 ) | ( ~n372 & n4756 ) | ( n4717 & n4756 ) ;
  assign n4758 = n372 | n4757 ;
  assign n4759 = ( n758 & ~n2324 ) | ( n758 & n4758 ) | ( ~n2324 & n4758 ) ;
  assign n4760 = n1035 | n4753 ;
  assign n4761 = n2324 | n4759 ;
  assign n4762 = ( n1712 & ~n2446 ) | ( n1712 & n4707 ) | ( ~n2446 & n4707 ) ;
  assign n4763 = n2446 | n4762 ;
  assign n4764 = ( ~n83 & n95 ) | ( ~n83 & n4763 ) | ( n95 & n4763 ) ;
  assign n4765 = ( ~n1051 & n1859 ) | ( ~n1051 & n4215 ) | ( n1859 & n4215 ) ;
  assign n4766 = n2098 | n4727 ;
  assign n4767 = n83 | n4764 ;
  assign n4768 = ( n437 & ~n605 ) | ( n437 & n4767 ) | ( ~n605 & n4767 ) ;
  assign n4769 = n605 | n4768 ;
  assign n4770 = ( n416 & ~n420 ) | ( n416 & n4769 ) | ( ~n420 & n4769 ) ;
  assign n4771 = n420 | n4770 ;
  assign n4772 = ( n88 & ~n578 ) | ( n88 & n4771 ) | ( ~n578 & n4771 ) ;
  assign n4773 = n578 | n4772 ;
  assign n4774 = n1798 | n1859 ;
  assign n4775 = n1467 | n3461 ;
  assign n4776 = n559 | n4773 ;
  assign n4777 = ( ~n2366 & n3906 ) | ( ~n2366 & n4776 ) | ( n3906 & n4776 ) ;
  assign n4778 = n2936 | n4776 ;
  assign n4779 = n652 & ~n4778 ;
  assign n4780 = n653 | n963 ;
  assign n4781 = n652 & ~n4704 ;
  assign n4782 = n433 | n943 ;
  assign n4783 = n4780 | n4782 ;
  assign n4784 = n4665 | n4783 ;
  assign n4785 = n4742 | n4784 ;
  assign n4786 = n150 | n3278 ;
  assign n4787 = n643 | n790 ;
  assign n4788 = n4786 | n4787 ;
  assign n4789 = n3554 | n4788 ;
  assign n4790 = n102 | n433 ;
  assign n4791 = n165 | n559 ;
  assign n4792 = ( n247 & ~n591 ) | ( n247 & n4789 ) | ( ~n591 & n4789 ) ;
  assign n4793 = n4790 | n4791 ;
  assign n4794 = n414 | n3461 ;
  assign n4795 = n591 | n4792 ;
  assign n4796 = ( n434 & ~n744 ) | ( n434 & n4795 ) | ( ~n744 & n4795 ) ;
  assign n4797 = n744 | n4796 ;
  assign n4798 = n580 | n4797 ;
  assign n4799 = n4783 | n4798 ;
  assign n4800 = n4228 | n4798 ;
  assign n4801 = n2278 & ~n4799 ;
  assign n4802 = ( n1485 & n4414 ) | ( n1485 & ~n4766 ) | ( n4414 & ~n4766 ) ;
  assign n4803 = n4766 | n4802 ;
  assign n4804 = ( n300 & ~n723 ) | ( n300 & n4803 ) | ( ~n723 & n4803 ) ;
  assign n4805 = n723 | n4804 ;
  assign n4806 = n232 | n4805 ;
  assign n4807 = n1722 | n4806 ;
  assign n4808 = ~n2476 & n4801 ;
  assign n4809 = ~n4776 & n4777 ;
  assign n4810 = n4793 | n4794 ;
  assign n4811 = ( ~n2480 & n4806 ) | ( ~n2480 & n4810 ) | ( n4806 & n4810 ) ;
  assign n4812 = n2480 | n4811 ;
  assign n4813 = ( n677 & ~n1258 ) | ( n677 & n4812 ) | ( ~n1258 & n4812 ) ;
  assign n4814 = n1258 | n4813 ;
  assign n4815 = ( n1859 & ~n2041 ) | ( n1859 & n4814 ) | ( ~n2041 & n4814 ) ;
  assign n4816 = ( n133 & ~n153 ) | ( n133 & n4531 ) | ( ~n153 & n4531 ) ;
  assign n4817 = n153 | n4816 ;
  assign n4818 = ( ~n94 & n255 ) | ( ~n94 & n4817 ) | ( n255 & n4817 ) ;
  assign n4819 = n94 | n4818 ;
  assign n4820 = ( n351 & ~n841 ) | ( n351 & n4819 ) | ( ~n841 & n4819 ) ;
  assign n4821 = n841 | n4820 ;
  assign n4822 = n827 | n4821 ;
  assign n4823 = ( ~n1740 & n4128 ) | ( ~n1740 & n4822 ) | ( n4128 & n4822 ) ;
  assign n4824 = n1740 | n4823 ;
  assign n4825 = ( ~n2028 & n4660 ) | ( ~n2028 & n4824 ) | ( n4660 & n4824 ) ;
  assign n4826 = ( n1986 & ~n2368 ) | ( n1986 & n4660 ) | ( ~n2368 & n4660 ) ;
  assign n4827 = n2368 | n4826 ;
  assign n4828 = n82 | n891 ;
  assign n4829 = n4822 | n4828 ;
  assign n4830 = n503 | n923 ;
  assign n4831 = n4396 | n4830 ;
  assign n4832 = n2158 | n4831 ;
  assign n4833 = ( n173 & ~n447 ) | ( n173 & n3711 ) | ( ~n447 & n3711 ) ;
  assign n4834 = n447 | n4833 ;
  assign n4835 = n4396 | n4829 ;
  assign n4836 = ( n90 & ~n605 ) | ( n90 & n4834 ) | ( ~n605 & n4834 ) ;
  assign n4837 = n605 | n4836 ;
  assign n4838 = ( n601 & ~n645 ) | ( n601 & n4837 ) | ( ~n645 & n4837 ) ;
  assign n4839 = n241 | n659 ;
  assign n4840 = n757 | n4839 ;
  assign n4841 = n645 | n4838 ;
  assign n4842 = n1250 | n4841 ;
  assign n4843 = n4829 | n4842 ;
  assign n4844 = n4807 | n4843 ;
  assign n4845 = n343 | n714 ;
  assign n4846 = n4840 | n4845 ;
  assign n4847 = n168 | n658 ;
  assign n4848 = ( n4258 & ~n4654 ) | ( n4258 & n4847 ) | ( ~n4654 & n4847 ) ;
  assign n4849 = n4800 | n4846 ;
  assign n4850 = n4563 | n4849 ;
  assign n4851 = ( ~n1248 & n1508 ) | ( ~n1248 & n4850 ) | ( n1508 & n4850 ) ;
  assign n4852 = n1248 | n4851 ;
  assign n4853 = ( ~n1308 & n4847 ) | ( ~n1308 & n4852 ) | ( n4847 & n4852 ) ;
  assign n4854 = ~n1417 & n4350 ;
  assign n4855 = ( ~n720 & n2541 ) | ( ~n720 & n4854 ) | ( n2541 & n4854 ) ;
  assign n4856 = n1308 | n4853 ;
  assign n4857 = n4654 | n4848 ;
  assign n4858 = ( ~n286 & n2937 ) | ( ~n286 & n4857 ) | ( n2937 & n4857 ) ;
  assign n4859 = ( ~n1478 & n2128 ) | ( ~n1478 & n4844 ) | ( n2128 & n4844 ) ;
  assign n4860 = n1478 | n4859 ;
  assign n4861 = ( ~n109 & n184 ) | ( ~n109 & n4856 ) | ( n184 & n4856 ) ;
  assign n4862 = ( ~n161 & n287 ) | ( ~n161 & n4860 ) | ( n287 & n4860 ) ;
  assign n4863 = n161 | n4862 ;
  assign n4864 = n109 | n4861 ;
  assign n4865 = ( ~n600 & n969 ) | ( ~n600 & n4864 ) | ( n969 & n4864 ) ;
  assign n4866 = n600 | n4865 ;
  assign n4867 = n651 | n4866 ;
  assign n4868 = n2659 | n4867 ;
  assign n4869 = n1828 | n4868 ;
  assign n4870 = ( ~n617 & n4841 ) | ( ~n617 & n4869 ) | ( n4841 & n4869 ) ;
  assign n4871 = n617 | n4870 ;
  assign n4872 = ( n720 & ~n2613 ) | ( n720 & n4871 ) | ( ~n2613 & n4871 ) ;
  assign n4873 = ( ~n116 & n1567 ) | ( ~n116 & n4863 ) | ( n1567 & n4863 ) ;
  assign n4874 = n954 | n4291 ;
  assign n4875 = n162 | n397 ;
  assign n4876 = n4311 | n4875 ;
  assign n4877 = n4300 | n4876 ;
  assign n4878 = ( n313 & ~n693 ) | ( n313 & n4877 ) | ( ~n693 & n4877 ) ;
  assign n4879 = n693 | n4878 ;
  assign n4880 = ( ~n288 & n499 ) | ( ~n288 & n4879 ) | ( n499 & n4879 ) ;
  assign n4881 = ~n918 & n4781 ;
  assign n4882 = n288 | n4880 ;
  assign n4883 = ( n375 & ~n522 ) | ( n375 & n4882 ) | ( ~n522 & n4882 ) ;
  assign n4884 = n522 | n4883 ;
  assign n4885 = ( n175 & ~n744 ) | ( n175 & n4884 ) | ( ~n744 & n4884 ) ;
  assign n4886 = n744 | n4885 ;
  assign n4887 = n2070 & ~n4886 ;
  assign n4888 = n229 | n559 ;
  assign n4889 = ( ~n918 & n2635 ) | ( ~n918 & n4887 ) | ( n2635 & n4887 ) ;
  assign n4890 = n145 | n2139 ;
  assign n4891 = n4888 | n4890 ;
  assign n4892 = n3633 | n4891 ;
  assign n4893 = n4867 | n4892 ;
  assign n4894 = n173 | n222 ;
  assign n4895 = n352 | n649 ;
  assign n4896 = n1318 | n4894 ;
  assign n4897 = n1248 | n2965 ;
  assign n4898 = n3832 | n4893 ;
  assign n4899 = n1756 | n2139 ;
  assign n4900 = n4895 | n4896 ;
  assign n4901 = n954 | n2541 ;
  assign n4902 = n1910 | n4414 ;
  assign n4903 = n4900 | n4902 ;
  assign n4904 = ( ~n414 & n778 ) | ( ~n414 & n4903 ) | ( n778 & n4903 ) ;
  assign n4905 = n414 | n4904 ;
  assign n4906 = n601 | n4905 ;
  assign n4907 = n2611 | n4724 ;
  assign n4908 = ( n1191 & ~n1630 ) | ( n1191 & n4907 ) | ( ~n1630 & n4907 ) ;
  assign n4909 = n1986 | n4906 ;
  assign n4910 = n2473 | n4909 ;
  assign n4911 = n4899 | n4901 ;
  assign n4912 = ( ~n3835 & n3948 ) | ( ~n3835 & n4906 ) | ( n3948 & n4906 ) ;
  assign n4913 = n3835 | n4912 ;
  assign n4914 = ( n1191 & ~n1248 ) | ( n1191 & n4913 ) | ( ~n1248 & n4913 ) ;
  assign n4915 = n1248 | n4914 ;
  assign n4916 = n744 | n2125 ;
  assign n4917 = n3699 | n4885 ;
  assign n4918 = n4916 | n4917 ;
  assign n4919 = n3392 | n4918 ;
  assign n4920 = ( n1382 & ~n2611 ) | ( n1382 & n2838 ) | ( ~n2611 & n2838 ) ;
  assign n4921 = ~n1382 & n4920 ;
  assign n4922 = ( ~n133 & n2663 ) | ( ~n133 & n4921 ) | ( n2663 & n4921 ) ;
  assign n4923 = ~n2663 & n4922 ;
  assign n4924 = ( ~n520 & n701 ) | ( ~n520 & n4923 ) | ( n701 & n4923 ) ;
  assign n4925 = ( ~n2098 & n3460 ) | ( ~n2098 & n4654 ) | ( n3460 & n4654 ) ;
  assign n4926 = ~n701 & n4924 ;
  assign n4927 = n2613 | n4872 ;
  assign n4928 = ( ~n489 & n555 ) | ( ~n489 & n4926 ) | ( n555 & n4926 ) ;
  assign n4929 = n2098 | n4925 ;
  assign n4930 = ~n555 & n4928 ;
  assign n4931 = ( n4332 & ~n4927 ) | ( n4332 & n4930 ) | ( ~n4927 & n4930 ) ;
  assign n4932 = ~n4332 & n4931 ;
  assign n4933 = ~n4785 & n4930 ;
  assign n4934 = n1388 | n2098 ;
  assign n4935 = ( n133 & ~n2549 ) | ( n133 & n4929 ) | ( ~n2549 & n4929 ) ;
  assign n4936 = n4282 | n4934 ;
  assign n4937 = n2246 | n3278 ;
  assign n4938 = n4200 | n4936 ;
  assign n4939 = n357 | n497 ;
  assign n4940 = n1910 | n4939 ;
  assign n4941 = n205 | n4939 ;
  assign n4942 = n787 | n4939 ;
  assign n4943 = n4937 | n4942 ;
  assign n4944 = n428 | n491 ;
  assign n4945 = n4941 | n4944 ;
  assign n4946 = n4874 | n4945 ;
  assign n4947 = n552 | n715 ;
  assign n4948 = ( ~n883 & n1382 ) | ( ~n883 & n4946 ) | ( n1382 & n4946 ) ;
  assign n4949 = n98 | n735 ;
  assign n4950 = n4947 | n4949 ;
  assign n4951 = n2729 | n4950 ;
  assign n4952 = n973 | n4951 ;
  assign n4953 = ( ~n957 & n4910 ) | ( ~n957 & n4952 ) | ( n4910 & n4952 ) ;
  assign n4954 = ( ~n1001 & n4424 ) | ( ~n1001 & n4952 ) | ( n4424 & n4952 ) ;
  assign n4955 = n1001 | n4954 ;
  assign n4956 = n957 | n4953 ;
  assign n4957 = ( ~n2613 & n4555 ) | ( ~n2613 & n4956 ) | ( n4555 & n4956 ) ;
  assign n4958 = n883 | n942 ;
  assign n4959 = n2613 | n4957 ;
  assign n4960 = n4930 & ~n4959 ;
  assign n4961 = ~n1388 & n4960 ;
  assign n4962 = ( ~n1349 & n2086 ) | ( ~n1349 & n4961 ) | ( n2086 & n4961 ) ;
  assign n4963 = n133 | n585 ;
  assign n4964 = n4958 | n4963 ;
  assign n4965 = ~n2086 & n4962 ;
  assign n4966 = n2961 | n4964 ;
  assign n4967 = ( n787 & ~n1159 ) | ( n787 & n4955 ) | ( ~n1159 & n4955 ) ;
  assign n4968 = n883 | n4948 ;
  assign n4969 = n4651 | n4966 ;
  assign n4970 = ( n88 & ~n358 ) | ( n88 & n4184 ) | ( ~n358 & n4184 ) ;
  assign n4971 = n358 | n4970 ;
  assign n4972 = ( n559 & ~n589 ) | ( n559 & n4971 ) | ( ~n589 & n4971 ) ;
  assign n4973 = n589 | n4972 ;
  assign n4974 = n271 | n4973 ;
  assign n4975 = n2390 | n4974 ;
  assign n4976 = n4964 | n4975 ;
  assign n4977 = n128 | n357 ;
  assign n4978 = n139 | n4977 ;
  assign n4979 = n3416 | n4978 ;
  assign n4980 = n4775 | n4979 ;
  assign n4981 = n302 | n643 ;
  assign n4982 = n693 | n4981 ;
  assign n4983 = n4316 | n4982 ;
  assign n4984 = n4978 | n4982 ;
  assign n4985 = n4976 | n4984 ;
  assign n4986 = n282 | n4500 ;
  assign n4987 = n313 | n422 ;
  assign n4988 = n731 | n4987 ;
  assign n4989 = n4986 | n4988 ;
  assign n4990 = ( ~n241 & n415 ) | ( ~n241 & n4989 ) | ( n415 & n4989 ) ;
  assign n4991 = n241 | n4990 ;
  assign n4992 = ( n147 & ~n810 ) | ( n147 & n4991 ) | ( ~n810 & n4991 ) ;
  assign n4993 = n810 | n4992 ;
  assign n4994 = ( ~n231 & n578 ) | ( ~n231 & n4993 ) | ( n578 & n4993 ) ;
  assign n4995 = n231 | n4994 ;
  assign n4996 = ( n2189 & ~n2713 ) | ( n2189 & n4995 ) | ( ~n2713 & n4995 ) ;
  assign n4997 = n2713 | n4996 ;
  assign n4998 = n248 | n965 ;
  assign n4999 = n420 | n4998 ;
  assign n5000 = ( ~n161 & n1518 ) | ( ~n161 & n4999 ) | ( n1518 & n4999 ) ;
  assign n5001 = n161 | n5000 ;
  assign n5002 = ( ~n197 & n593 ) | ( ~n197 & n5001 ) | ( n593 & n5001 ) ;
  assign n5003 = n197 | n5002 ;
  assign n5004 = ( n122 & ~n717 ) | ( n122 & n5003 ) | ( ~n717 & n5003 ) ;
  assign n5005 = n717 | n5004 ;
  assign n5006 = n601 | n5005 ;
  assign n5007 = n154 | n161 ;
  assign n5008 = ( n3212 & n4985 ) | ( n3212 & ~n5006 ) | ( n4985 & ~n5006 ) ;
  assign n5009 = n148 | n719 ;
  assign n5010 = n2603 | n4500 ;
  assign n5011 = n111 | n4572 ;
  assign n5012 = n4875 | n5009 ;
  assign n5013 = ( n1818 & ~n4997 ) | ( n1818 & n5006 ) | ( ~n4997 & n5006 ) ;
  assign n5014 = n5011 | n5012 ;
  assign n5015 = n4997 | n5013 ;
  assign n5016 = n197 | n357 ;
  assign n5017 = n5007 | n5016 ;
  assign n5018 = n5006 | n5008 ;
  assign n5019 = n1151 | n5017 ;
  assign n5020 = ( ~n2669 & n3699 ) | ( ~n2669 & n5018 ) | ( n3699 & n5018 ) ;
  assign n5021 = n3346 | n5019 ;
  assign n5022 = n4983 | n5021 ;
  assign n5023 = n1008 | n5017 ;
  assign n5024 = n4898 | n5023 ;
  assign n5025 = n2669 | n5020 ;
  assign n5026 = n1251 | n4875 ;
  assign n5027 = ~n1663 & n3616 ;
  assign n5028 = ( ~n1136 & n2994 ) | ( ~n1136 & n5027 ) | ( n2994 & n5027 ) ;
  assign n5029 = ~n2994 & n5028 ;
  assign n5030 = ( ~n287 & n1860 ) | ( ~n287 & n5029 ) | ( n1860 & n5029 ) ;
  assign n5031 = ~n1860 & n5030 ;
  assign n5032 = ( n96 & ~n167 ) | ( n96 & n5031 ) | ( ~n167 & n5031 ) ;
  assign n5033 = n232 | n247 ;
  assign n5034 = ( ~n1338 & n3962 ) | ( ~n1338 & n5015 ) | ( n3962 & n5015 ) ;
  assign n5035 = n102 | n5033 ;
  assign n5036 = ( n1134 & n3370 ) | ( n1134 & ~n5035 ) | ( n3370 & ~n5035 ) ;
  assign n5037 = n5035 | n5036 ;
  assign n5038 = ( ~n888 & n3962 ) | ( ~n888 & n5037 ) | ( n3962 & n5037 ) ;
  assign n5039 = n888 | n5038 ;
  assign n5040 = ( n1071 & ~n1136 ) | ( n1071 & n5039 ) | ( ~n1136 & n5039 ) ;
  assign n5041 = n650 | n1520 ;
  assign n5042 = ~n96 & n5032 ;
  assign n5043 = n499 | n5041 ;
  assign n5044 = ( n88 & ~n721 ) | ( n88 & n5042 ) | ( ~n721 & n5042 ) ;
  assign n5045 = ~n88 & n5044 ;
  assign n5046 = n4892 | n5043 ;
  assign n5047 = n1224 | n5046 ;
  assign n5048 = n461 | n593 ;
  assign n5049 = n757 | n5048 ;
  assign n5050 = ( ~n116 & n943 ) | ( ~n116 & n3601 ) | ( n943 & n3601 ) ;
  assign n5051 = n116 | n5050 ;
  assign n5052 = ( n111 & ~n162 ) | ( n111 & n5051 ) | ( ~n162 & n5051 ) ;
  assign n5053 = ~n146 & n5045 ;
  assign n5054 = n4587 & ~n4654 ;
  assign n5055 = ~n888 & n5054 ;
  assign n5056 = n342 | n601 ;
  assign n5057 = n4144 | n5041 ;
  assign n5058 = n4974 | n5049 ;
  assign n5059 = n1134 | n2429 ;
  assign n5060 = n162 | n5052 ;
  assign n5061 = n4896 | n5035 ;
  assign n5062 = n2817 | n5052 ;
  assign n5063 = n4010 | n5061 ;
  assign n5064 = n175 | n5049 ;
  assign n5065 = n197 | n248 ;
  assign n5066 = n5056 | n5065 ;
  assign n5067 = n5064 | n5066 ;
  assign n5068 = ( ~n2998 & n4172 ) | ( ~n2998 & n5063 ) | ( n4172 & n5063 ) ;
  assign n5069 = n2998 | n5068 ;
  assign n5070 = ( ~n5035 & n5047 ) | ( ~n5035 & n5053 ) | ( n5047 & n5053 ) ;
  assign n5071 = ( ~n2515 & n5053 ) | ( ~n2515 & n5067 ) | ( n5053 & n5067 ) ;
  assign n5072 = ~n5067 & n5071 ;
  assign n5073 = ( n1134 & ~n5060 ) | ( n1134 & n5072 ) | ( ~n5060 & n5072 ) ;
  assign n5074 = ~n1134 & n5073 ;
  assign n5075 = ~n5047 & n5070 ;
  assign n5076 = ~n4736 & n5075 ;
  assign n5077 = ( n491 & ~n1922 ) | ( n491 & n5074 ) | ( ~n1922 & n5074 ) ;
  assign n5078 = ( ~n1485 & n3266 ) | ( ~n1485 & n4897 ) | ( n3266 & n4897 ) ;
  assign n5079 = ( ~n84 & n796 ) | ( ~n84 & n5025 ) | ( n796 & n5025 ) ;
  assign n5080 = n1485 | n5078 ;
  assign n5081 = ( n288 & ~n437 ) | ( n288 & n5080 ) | ( ~n437 & n5080 ) ;
  assign n5082 = n84 | n5079 ;
  assign n5083 = ( n288 & ~n790 ) | ( n288 & n5082 ) | ( ~n790 & n5082 ) ;
  assign n5084 = n147 | n532 ;
  assign n5085 = n91 | n5084 ;
  assign n5086 = n2220 | n5085 ;
  assign n5087 = n4943 | n5086 ;
  assign n5088 = ( ~n84 & n289 ) | ( ~n84 & n5087 ) | ( n289 & n5087 ) ;
  assign n5089 = n84 | n5088 ;
  assign n5090 = n87 | n499 ;
  assign n5091 = ( ~n84 & n1318 ) | ( ~n84 & n4398 ) | ( n1318 & n4398 ) ;
  assign n5092 = n84 | n5091 ;
  assign n5093 = ( n1529 & n5062 ) | ( n1529 & ~n5085 ) | ( n5062 & ~n5085 ) ;
  assign n5094 = ( ~n561 & n1529 ) | ( ~n561 & n4622 ) | ( n1529 & n4622 ) ;
  assign n5095 = n109 | n211 ;
  assign n5096 = n93 | n5095 ;
  assign n5097 = n5090 | n5096 ;
  assign n5098 = n786 | n2795 ;
  assign n5099 = n2128 | n5098 ;
  assign n5100 = n125 | n351 ;
  assign n5101 = n694 | n5100 ;
  assign n5102 = n2001 | n5101 ;
  assign n5103 = n5097 | n5102 ;
  assign n5104 = n5099 | n5103 ;
  assign n5105 = n2572 | n5104 ;
  assign n5106 = ( ~n1308 & n4232 ) | ( ~n1308 & n5105 ) | ( n4232 & n5105 ) ;
  assign n5107 = n1308 | n5106 ;
  assign n5108 = ( n3637 & ~n5085 ) | ( n3637 & n5107 ) | ( ~n5085 & n5107 ) ;
  assign n5109 = n5085 | n5108 ;
  assign n5110 = ( ~n81 & n289 ) | ( ~n81 & n5109 ) | ( n289 & n5109 ) ;
  assign n5111 = n81 | n5110 ;
  assign n5112 = ( ~n161 & n607 ) | ( ~n161 & n5111 ) | ( n607 & n5111 ) ;
  assign n5113 = n161 | n5112 ;
  assign n5114 = ( n295 & ~n420 ) | ( n295 & n5113 ) | ( ~n420 & n5113 ) ;
  assign n5115 = n420 | n5114 ;
  assign n5116 = ( ~n100 & n148 ) | ( ~n100 & n5115 ) | ( n148 & n5115 ) ;
  assign n5117 = n100 | n5116 ;
  assign n5118 = ( n3723 & ~n4158 ) | ( n3723 & n5117 ) | ( ~n4158 & n5117 ) ;
  assign n5119 = n1593 | n5117 ;
  assign n5120 = n4158 | n5118 ;
  assign n5121 = n1816 | n5103 ;
  assign n5122 = n4575 | n5119 ;
  assign n5123 = n3822 | n5122 ;
  assign n5124 = ( ~n4090 & n5067 ) | ( ~n4090 & n5120 ) | ( n5067 & n5120 ) ;
  assign n5125 = n4090 | n5124 ;
  assign n5126 = n561 | n5094 ;
  assign n5127 = ( ~n93 & n3637 ) | ( ~n93 & n5126 ) | ( n3637 & n5126 ) ;
  assign n5128 = n362 | n602 ;
  assign n5129 = n510 | n5128 ;
  assign n5130 = n1051 | n5129 ;
  assign n5131 = ( ~n714 & n3539 ) | ( ~n714 & n4413 ) | ( n3539 & n4413 ) ;
  assign n5132 = n714 | n5131 ;
  assign n5133 = ( n653 & ~n756 ) | ( n653 & n5132 ) | ( ~n756 & n5132 ) ;
  assign n5134 = n756 | n5133 ;
  assign n5135 = n701 | n5134 ;
  assign n5136 = n4627 | n5135 ;
  assign n5137 = n5130 | n5136 ;
  assign n5138 = n5121 | n5137 ;
  assign n5139 = ( ~n212 & n234 ) | ( ~n212 & n5138 ) | ( n234 & n5138 ) ;
  assign n5140 = n212 | n5139 ;
  assign n5141 = ( n683 & ~n829 ) | ( n683 & n5140 ) | ( ~n829 & n5140 ) ;
  assign n5142 = n829 | n5141 ;
  assign n5143 = ( ~n503 & n1333 ) | ( ~n503 & n5142 ) | ( n1333 & n5142 ) ;
  assign n5144 = n503 | n5143 ;
  assign n5145 = ( n345 & ~n723 ) | ( n345 & n5144 ) | ( ~n723 & n5144 ) ;
  assign n5146 = n723 | n5145 ;
  assign n5147 = ( ~n580 & n833 ) | ( ~n580 & n5146 ) | ( n833 & n5146 ) ;
  assign n5148 = n580 | n5147 ;
  assign n5149 = n530 | n5148 ;
  assign n5150 = n2535 | n5149 ;
  assign n5151 = n5026 | n5150 ;
  assign n5152 = n5058 | n5151 ;
  assign n5153 = n1192 | n3637 ;
  assign n5154 = n2635 | n5129 ;
  assign n5155 = n3865 & ~n5154 ;
  assign n5156 = n2218 | n4446 ;
  assign n5157 = n790 | n5083 ;
  assign n5158 = ( n417 & ~n735 ) | ( n417 & n5157 ) | ( ~n735 & n5157 ) ;
  assign n5159 = n735 | n5158 ;
  assign n5160 = n378 | n5159 ;
  assign n5161 = n4437 | n5149 ;
  assign n5162 = n4612 | n5161 ;
  assign n5163 = ( n2218 & ~n4995 ) | ( n2218 & n5162 ) | ( ~n4995 & n5162 ) ;
  assign n5164 = n4995 | n5163 ;
  assign n5165 = n5160 | n5164 ;
  assign n5166 = ( n677 & ~n1144 ) | ( n677 & n5165 ) | ( ~n1144 & n5165 ) ;
  assign n5167 = n1144 | n5166 ;
  assign n5168 = ( n557 & ~n2994 ) | ( n557 & n5167 ) | ( ~n2994 & n5167 ) ;
  assign n5169 = n2994 | n5168 ;
  assign n5170 = ( ~n916 & n3637 ) | ( ~n916 & n5169 ) | ( n3637 & n5169 ) ;
  assign n5171 = n180 | n4471 ;
  assign n5172 = ( n2275 & ~n2939 ) | ( n2275 & n4414 ) | ( ~n2939 & n4414 ) ;
  assign n5173 = ( n546 & ~n960 ) | ( n546 & n3716 ) | ( ~n960 & n3716 ) ;
  assign n5174 = ( n879 & ~n1345 ) | ( n879 & n5171 ) | ( ~n1345 & n5171 ) ;
  assign n5175 = n1345 | n5174 ;
  assign n5176 = n960 | n5173 ;
  assign n5177 = n1345 | n4999 ;
  assign n5178 = ( ~n279 & n647 ) | ( ~n279 & n5176 ) | ( n647 & n5176 ) ;
  assign n5179 = ( ~n489 & n701 ) | ( ~n489 & n4832 ) | ( n701 & n4832 ) ;
  assign n5180 = n3425 | n5178 ;
  assign n5181 = n279 | n5178 ;
  assign n5182 = ( ~n2613 & n5155 ) | ( ~n2613 & n5181 ) | ( n5155 & n5181 ) ;
  assign n5183 = ~n5181 & n5182 ;
  assign n5184 = ( n550 & ~n4018 ) | ( n550 & n5183 ) | ( ~n4018 & n5183 ) ;
  assign n5185 = n220 | n250 ;
  assign n5186 = n489 | n5179 ;
  assign n5187 = ~n550 & n5184 ;
  assign n5188 = n203 | n247 ;
  assign n5189 = n400 | n3819 ;
  assign n5190 = n5185 | n5188 ;
  assign n5191 = n5043 | n5190 ;
  assign n5192 = n3985 | n5191 ;
  assign n5193 = n184 | n422 ;
  assign n5194 = n105 | n356 ;
  assign n5195 = n220 | n433 ;
  assign n5196 = n5194 | n5195 ;
  assign n5197 = n417 | n786 ;
  assign n5198 = ( n245 & ~n372 ) | ( n245 & n5186 ) | ( ~n372 & n5186 ) ;
  assign n5199 = n5193 | n5197 ;
  assign n5200 = n5177 | n5199 ;
  assign n5201 = n228 | n293 ;
  assign n5202 = n4227 | n5201 ;
  assign n5203 = ( ~n90 & n973 ) | ( ~n90 & n5202 ) | ( n973 & n5202 ) ;
  assign n5204 = n90 | n5203 ;
  assign n5205 = ( n2743 & ~n4232 ) | ( n2743 & n5204 ) | ( ~n4232 & n5204 ) ;
  assign n5206 = ( n56 & ~n1340 ) | ( n56 & n5200 ) | ( ~n1340 & n5200 ) ;
  assign n5207 = ( ~n4414 & n5123 ) | ( ~n4414 & n5204 ) | ( n5123 & n5204 ) ;
  assign n5208 = ~n4414 & n5172 ;
  assign n5209 = n4414 | n5207 ;
  assign n5210 = n4774 | n5196 ;
  assign n5211 = n372 | n5198 ;
  assign n5212 = n5190 | n5211 ;
  assign n5213 = ( n3413 & ~n5117 ) | ( n3413 & n5212 ) | ( ~n5117 & n5212 ) ;
  assign n5214 = n5117 | n5213 ;
  assign n5215 = ( ~n1745 & n5189 ) | ( ~n1745 & n5214 ) | ( n5189 & n5214 ) ;
  assign n5216 = ( n116 & ~n342 ) | ( n116 & n4542 ) | ( ~n342 & n4542 ) ;
  assign n5217 = ~n116 & n5216 ;
  assign n5218 = ( ~n714 & n786 ) | ( ~n714 & n5217 ) | ( n786 & n5217 ) ;
  assign n5219 = ~n786 & n5218 ;
  assign n5220 = ( n111 & ~n827 ) | ( n111 & n5219 ) | ( ~n827 & n5219 ) ;
  assign n5221 = ~n111 & n5220 ;
  assign n5222 = ~n2827 & n5221 ;
  assign n5223 = ~n5205 & n5221 ;
  assign n5224 = n100 | n650 ;
  assign n5225 = n497 | n5224 ;
  assign n5226 = n5101 | n5225 ;
  assign n5227 = n4911 | n5226 ;
  assign n5228 = n212 | n520 ;
  assign n5229 = ~n1417 & n5222 ;
  assign n5230 = n289 | n371 ;
  assign n5231 = n96 | n336 ;
  assign n5232 = ( ~n83 & n341 ) | ( ~n83 & n5227 ) | ( n341 & n5227 ) ;
  assign n5233 = n83 | n5232 ;
  assign n5234 = ( ~n532 & n628 ) | ( ~n532 & n5233 ) | ( n628 & n5233 ) ;
  assign n5235 = n532 | n5234 ;
  assign n5236 = n759 | n846 ;
  assign n5237 = n1190 | n5135 ;
  assign n5238 = ( ~n1712 & n5187 ) | ( ~n1712 & n5236 ) | ( n5187 & n5236 ) ;
  assign n5239 = ( n410 & ~n580 ) | ( n410 & n5235 ) | ( ~n580 & n5235 ) ;
  assign n5240 = n2122 | n5239 ;
  assign n5241 = ~n5236 & n5238 ;
  assign n5242 = ( n139 & ~n823 ) | ( n139 & n5241 ) | ( ~n823 & n5241 ) ;
  assign n5243 = n5228 | n5230 ;
  assign n5244 = n5231 | n5243 ;
  assign n5245 = n2169 | n5239 ;
  assign n5246 = ( n719 & ~n778 ) | ( n719 & n5244 ) | ( ~n778 & n5244 ) ;
  assign n5247 = n778 | n5246 ;
  assign n5248 = n2101 | n5247 ;
  assign n5249 = ( n3836 & ~n5211 ) | ( n3836 & n5247 ) | ( ~n5211 & n5247 ) ;
  assign n5250 = ~n139 & n5242 ;
  assign n5251 = ( ~n90 & n148 ) | ( ~n90 & n5250 ) | ( n148 & n5250 ) ;
  assign n5252 = ~n148 & n5251 ;
  assign n5253 = ~n5247 & n5249 ;
  assign n5254 = ( n5245 & ~n5248 ) | ( n5245 & n5252 ) | ( ~n5248 & n5252 ) ;
  assign n5255 = ~n5245 & n5254 ;
  assign n5256 = ~n2170 & n5252 ;
  assign n5257 = ~n5237 & n5256 ;
  assign n5258 = ~n5156 & n5257 ;
  assign n5259 = ( n1095 & ~n4172 ) | ( n1095 & n5024 ) | ( ~n4172 & n5024 ) ;
  assign n5260 = ( ~n650 & n702 ) | ( ~n650 & n5210 ) | ( n702 & n5210 ) ;
  assign n5261 = n372 | n3578 ;
  assign n5262 = ( ~n304 & n3963 ) | ( ~n304 & n4099 ) | ( n3963 & n4099 ) ;
  assign n5263 = n650 | n5260 ;
  assign n5264 = ( n206 & ~n372 ) | ( n206 & n5263 ) | ( ~n372 & n5263 ) ;
  assign n5265 = n5261 | n5264 ;
  assign n5266 = ( ~n180 & n607 ) | ( ~n180 & n5265 ) | ( n607 & n5265 ) ;
  assign n5267 = n180 | n5266 ;
  assign n5268 = ( ~n1382 & n3117 ) | ( ~n1382 & n4743 ) | ( n3117 & n4743 ) ;
  assign n5269 = n1382 | n5268 ;
  assign n5270 = ( ~n105 & n221 ) | ( ~n105 & n4490 ) | ( n221 & n4490 ) ;
  assign n5271 = n2322 | n5099 ;
  assign n5272 = ( ~n128 & n520 ) | ( ~n128 & n5267 ) | ( n520 & n5267 ) ;
  assign n5273 = n128 | n5272 ;
  assign n5274 = ( ~n1088 & n2108 ) | ( ~n1088 & n2569 ) | ( n2108 & n2569 ) ;
  assign n5275 = n362 | n5273 ;
  assign n5276 = n4172 | n5259 ;
  assign n5277 = n1088 | n5274 ;
  assign n5278 = ( ~n105 & n2185 ) | ( ~n105 & n5277 ) | ( n2185 & n5277 ) ;
  assign n5279 = ( n424 & ~n2663 ) | ( n424 & n5269 ) | ( ~n2663 & n5269 ) ;
  assign n5280 = n105 | n5278 ;
  assign n5281 = ( n1382 & ~n2446 ) | ( n1382 & n5276 ) | ( ~n2446 & n5276 ) ;
  assign n5282 = n271 | n530 ;
  assign n5283 = n1056 | n5282 ;
  assign n5284 = n1926 | n5283 ;
  assign n5285 = n2310 & ~n5284 ;
  assign n5286 = n2322 | n5283 ;
  assign n5287 = n2663 | n5279 ;
  assign n5288 = ( n1975 & ~n5275 ) | ( n1975 & n5287 ) | ( ~n5275 & n5287 ) ;
  assign n5289 = n304 | n5262 ;
  assign n5290 = n5275 | n5288 ;
  assign n5291 = ( ~n683 & n2185 ) | ( ~n683 & n5290 ) | ( n2185 & n5290 ) ;
  assign n5292 = n206 | n601 ;
  assign n5293 = n5286 | n5292 ;
  assign n5294 = n683 | n5291 ;
  assign n5295 = ( n1975 & ~n2030 ) | ( n1975 & n5285 ) | ( ~n2030 & n5285 ) ;
  assign n5296 = ~n1975 & n5295 ;
  assign n5297 = ( n1712 & ~n2551 ) | ( n1712 & n5296 ) | ( ~n2551 & n5296 ) ;
  assign n5298 = ~n1712 & n5297 ;
  assign n5299 = ( ~n128 & n649 ) | ( ~n128 & n5289 ) | ( n649 & n5289 ) ;
  assign n5300 = n128 | n5299 ;
  assign n5301 = ( ~n1309 & n4063 ) | ( ~n1309 & n5180 ) | ( n4063 & n5180 ) ;
  assign n5302 = n1309 | n5301 ;
  assign n5303 = ( ~n796 & n2541 ) | ( ~n796 & n5302 ) | ( n2541 & n5302 ) ;
  assign n5304 = n796 | n5303 ;
  assign n5305 = ( ~n290 & n3539 ) | ( ~n290 & n5304 ) | ( n3539 & n5304 ) ;
  assign n5306 = n290 | n5305 ;
  assign n5307 = n796 | n4435 ;
  assign n5308 = n184 | n891 ;
  assign n5309 = n5010 | n5308 ;
  assign n5310 = ( ~n211 & n246 ) | ( ~n211 & n5306 ) | ( n246 & n5306 ) ;
  assign n5311 = n631 | n810 ;
  assign n5312 = n5309 | n5311 ;
  assign n5313 = n4779 & ~n5312 ;
  assign n5314 = n211 | n5310 ;
  assign n5315 = ( ~n644 & n1333 ) | ( ~n644 & n5314 ) | ( n1333 & n5314 ) ;
  assign n5316 = n644 | n5315 ;
  assign n5317 = n717 | n4153 ;
  assign n5318 = ( ~n2909 & n3539 ) | ( ~n2909 & n4760 ) | ( n3539 & n4760 ) ;
  assign n5319 = ~n2108 & n3892 ;
  assign n5320 = ( n88 & ~n717 ) | ( n88 & n5316 ) | ( ~n717 & n5316 ) ;
  assign n5321 = n717 | n3081 ;
  assign n5322 = n717 | n5320 ;
  assign n5323 = n2909 | n5318 ;
  assign n5324 = n5317 | n5320 ;
  assign n5325 = ( ~n659 & n4232 ) | ( ~n659 & n5324 ) | ( n4232 & n5324 ) ;
  assign n5326 = ( n246 & ~n423 ) | ( n246 & n5323 ) | ( ~n423 & n5323 ) ;
  assign n5327 = n1136 | n5040 ;
  assign n5328 = ( ~n1095 & n4452 ) | ( ~n1095 & n5152 ) | ( n4452 & n5152 ) ;
  assign n5329 = ~n4232 & n5223 ;
  assign n5330 = ( ~n428 & n1354 ) | ( ~n428 & n5313 ) | ( n1354 & n5313 ) ;
  assign n5331 = n4012 & ~n5322 ;
  assign n5332 = ( n332 & ~n631 ) | ( n332 & n5327 ) | ( ~n631 & n5327 ) ;
  assign n5333 = n631 | n5332 ;
  assign n5334 = ~n361 & n5319 ;
  assign n5335 = ( n173 & ~n631 ) | ( n173 & n4650 ) | ( ~n631 & n4650 ) ;
  assign n5336 = ( ~n424 & n4452 ) | ( ~n424 & n5334 ) | ( n4452 & n5334 ) ;
  assign n5337 = n5320 | n5321 ;
  assign n5338 = ~n4452 & n5336 ;
  assign n5339 = ( n1085 & ~n1630 ) | ( n1085 & n5337 ) | ( ~n1630 & n5337 ) ;
  assign n5340 = n655 | n3951 ;
  assign n5341 = ( ~n102 & n3598 ) | ( ~n102 & n5033 ) | ( n3598 & n5033 ) ;
  assign n5342 = ( n1745 & ~n1756 ) | ( n1745 & n5340 ) | ( ~n1756 & n5340 ) ;
  assign n5343 = n1756 | n5342 ;
  assign n5344 = n146 | n825 ;
  assign n5345 = ( n1756 & ~n4569 ) | ( n1756 & n5344 ) | ( ~n4569 & n5344 ) ;
  assign n5346 = n4569 | n5345 ;
  assign n5347 = n2041 | n4815 ;
  assign n5348 = ( ~n437 & n3175 ) | ( ~n437 & n5346 ) | ( n3175 & n5346 ) ;
  assign n5349 = ( ~n3491 & n5209 ) | ( ~n3491 & n5236 ) | ( n5209 & n5236 ) ;
  assign n5350 = ~n424 & n4522 ;
  assign n5351 = ( ~n1246 & n1860 ) | ( ~n1246 & n4968 ) | ( n1860 & n4968 ) ;
  assign n5352 = n437 | n5348 ;
  assign n5353 = ( ~n468 & n593 ) | ( ~n468 & n5352 ) | ( n593 & n5352 ) ;
  assign n5354 = n1246 | n4700 ;
  assign n5355 = ( n2549 & n4114 ) | ( n2549 & ~n4840 ) | ( n4114 & ~n4840 ) ;
  assign n5356 = n279 | n547 ;
  assign n5357 = n3491 | n5349 ;
  assign n5358 = n1860 | n5354 ;
  assign n5359 = ( n336 & ~n417 ) | ( n336 & n5357 ) | ( ~n417 & n5357 ) ;
  assign n5360 = ( n116 & ~n144 ) | ( n116 & n4965 ) | ( ~n144 & n4965 ) ;
  assign n5361 = n468 | n5353 ;
  assign n5362 = ( n1371 & ~n1983 ) | ( n1371 & n5361 ) | ( ~n1983 & n5361 ) ;
  assign n5363 = ( ~n4840 & n5329 ) | ( ~n4840 & n5361 ) | ( n5329 & n5361 ) ;
  assign n5364 = ~n5361 & n5363 ;
  assign n5365 = n109 | n111 ;
  assign n5366 = n1983 | n5362 ;
  assign n5367 = n188 | n468 ;
  assign n5368 = n5356 | n5367 ;
  assign n5369 = n5365 | n5368 ;
  assign n5370 = n4266 | n5369 ;
  assign n5371 = n3279 | n5370 ;
  assign n5372 = ~n5033 & n5341 ;
  assign n5373 = n98 | n872 ;
  assign n5374 = n444 | n5373 ;
  assign n5375 = n5369 | n5374 ;
  assign n5376 = n4142 | n5375 ;
  assign n5377 = ( ~n424 & n2997 ) | ( ~n424 & n5376 ) | ( n2997 & n5376 ) ;
  assign n5378 = n424 | n5377 ;
  assign n5379 = ( ~n1520 & n1860 ) | ( ~n1520 & n5378 ) | ( n1860 & n5378 ) ;
  assign n5380 = n1520 | n5379 ;
  assign n5381 = ( ~n82 & n336 ) | ( ~n82 & n5380 ) | ( n336 & n5380 ) ;
  assign n5382 = n82 | n5381 ;
  assign n5383 = ( ~n211 & n304 ) | ( ~n211 & n5382 ) | ( n304 & n5382 ) ;
  assign n5384 = n211 | n5383 ;
  assign n5385 = ( ~n559 & n4919 ) | ( ~n559 & n5384 ) | ( n4919 & n5384 ) ;
  assign n5386 = n559 | n5385 ;
  assign n5387 = n559 | n5384 ;
  assign n5388 = ( n1446 & n4980 ) | ( n1446 & ~n5387 ) | ( n4980 & ~n5387 ) ;
  assign n5389 = n5387 | n5388 ;
  assign n5390 = ( ~n559 & n5372 ) | ( ~n559 & n5384 ) | ( n5372 & n5384 ) ;
  assign n5391 = ~n5384 & n5390 ;
  assign n5392 = ( n2077 & ~n4840 ) | ( n2077 & n5386 ) | ( ~n4840 & n5386 ) ;
  assign n5393 = n3098 | n5374 ;
  assign n5394 = ( ~n1136 & n2041 ) | ( ~n1136 & n5391 ) | ( n2041 & n5391 ) ;
  assign n5395 = ~n2041 & n5394 ;
  assign n5396 = ( ~n144 & n786 ) | ( ~n144 & n5395 ) | ( n786 & n5395 ) ;
  assign n5397 = n4840 | n5392 ;
  assign n5398 = ( n860 & ~n4018 ) | ( n860 & n5397 ) | ( ~n4018 & n5397 ) ;
  assign n5399 = n1745 | n5215 ;
  assign n5400 = n1745 | n3241 ;
  assign n5401 = ~n1745 & n4933 ;
  assign n5402 = ~n2549 & n5355 ;
  assign n5403 = ( n1544 & ~n2939 ) | ( n1544 & n5402 ) | ( ~n2939 & n5402 ) ;
  assign n5404 = ~n1544 & n5403 ;
  assign n5405 = ( ~n2613 & n4654 ) | ( ~n2613 & n4969 ) | ( n4654 & n4969 ) ;
  assign n5406 = n2613 | n5405 ;
  assign n5407 = ( ~n1544 & n2541 ) | ( ~n1544 & n5406 ) | ( n2541 & n5406 ) ;
  assign n5408 = n1544 | n5407 ;
  assign n5409 = n222 | n349 ;
  assign n5410 = n214 | n846 ;
  assign n5411 = n5409 | n5410 ;
  assign n5412 = n2177 | n5409 ;
  assign n5413 = n183 | n965 ;
  assign n5414 = ~n2541 & n4855 ;
  assign n5415 = ~n1308 & n3259 ;
  assign n5416 = ( ~n1051 & n2108 ) | ( ~n1051 & n5399 ) | ( n2108 & n5399 ) ;
  assign n5417 = n2939 | n3977 ;
  assign n5418 = ~n161 & n4000 ;
  assign n5419 = n2098 | n2108 ;
  assign n5420 = ( ~n183 & n247 ) | ( ~n183 & n5418 ) | ( n247 & n5418 ) ;
  assign n5421 = n188 | n5413 ;
  assign n5422 = ( ~n225 & n5415 ) | ( ~n225 & n5421 ) | ( n5415 & n5421 ) ;
  assign n5423 = n1190 | n5421 ;
  assign n5424 = n5419 | n5423 ;
  assign n5425 = n3419 | n5424 ;
  assign n5426 = n3110 & ~n5425 ;
  assign n5427 = ~n1520 & n5426 ;
  assign n5428 = n234 | n448 ;
  assign n5429 = n5411 | n5428 ;
  assign n5430 = ( ~n182 & n434 ) | ( ~n182 & n5429 ) | ( n434 & n5429 ) ;
  assign n5431 = ( ~n342 & n923 ) | ( ~n342 & n5427 ) | ( n923 & n5427 ) ;
  assign n5432 = n182 | n5430 ;
  assign n5433 = n601 | n5432 ;
  assign n5434 = ~n923 & n5431 ;
  assign n5435 = ( ~n1001 & n5389 ) | ( ~n1001 & n5433 ) | ( n5389 & n5433 ) ;
  assign n5436 = ( n100 & ~n232 ) | ( n100 & n5434 ) | ( ~n232 & n5434 ) ;
  assign n5437 = ~n100 & n5436 ;
  assign n5438 = ~n111 & n5437 ;
  assign n5439 = ~n4375 & n5438 ;
  assign n5440 = ~n5433 & n5439 ;
  assign n5441 = ~n4835 & n5440 ;
  assign n5442 = n1001 | n5435 ;
  assign n5443 = ~n5022 & n5438 ;
  assign n5444 = ( ~n2053 & n4137 ) | ( ~n2053 & n5441 ) | ( n4137 & n5441 ) ;
  assign n5445 = ( n2541 & ~n2939 ) | ( n2541 & n5442 ) | ( ~n2939 & n5442 ) ;
  assign n5446 = ~n4137 & n5444 ;
  assign n5447 = n2939 | n5445 ;
  assign n5448 = ( ~n95 & n1367 ) | ( ~n95 & n5350 ) | ( n1367 & n5350 ) ;
  assign n5449 = ~n1367 & n5448 ;
  assign n5450 = ( ~n829 & n1333 ) | ( ~n829 & n5449 ) | ( n1333 & n5449 ) ;
  assign n5451 = ~n1333 & n5450 ;
  assign n5452 = ( n295 & ~n891 ) | ( n295 & n3619 ) | ( ~n891 & n3619 ) ;
  assign n5453 = n891 | n5452 ;
  assign n5454 = ( n232 & n583 ) | ( n232 & ~n5453 ) | ( n583 & ~n5453 ) ;
  assign n5455 = ~n232 & n5454 ;
  assign n5456 = ( ~n367 & n608 ) | ( ~n367 & n5455 ) | ( n608 & n5455 ) ;
  assign n5457 = ~n608 & n5456 ;
  assign n5458 = ( ~n4063 & n5371 ) | ( ~n4063 & n5457 ) | ( n5371 & n5457 ) ;
  assign n5459 = ~n5371 & n5458 ;
  assign n5460 = ~n5275 & n5459 ;
  assign n5461 = ( n2030 & ~n3175 ) | ( n2030 & n4561 ) | ( ~n3175 & n4561 ) ;
  assign n5462 = n4555 | n4556 ;
  assign n5463 = ( ~n1307 & n4063 ) | ( ~n1307 & n5462 ) | ( n4063 & n5462 ) ;
  assign n5464 = n1307 | n5463 ;
  assign n5465 = ( ~n313 & n593 ) | ( ~n313 & n5464 ) | ( n593 & n5464 ) ;
  assign n5466 = n313 | n5465 ;
  assign n5467 = ( n96 & ~n649 ) | ( n96 & n5466 ) | ( ~n649 & n5466 ) ;
  assign n5468 = n649 | n5467 ;
  assign n5469 = ( n139 & ~n547 ) | ( n139 & n5468 ) | ( ~n547 & n5468 ) ;
  assign n5470 = n547 | n5469 ;
  assign n5471 = ( ~n89 & n701 ) | ( ~n89 & n5470 ) | ( n701 & n5470 ) ;
  assign n5472 = n89 | n5471 ;
  assign n5473 = n4740 | n5472 ;
  assign n5474 = ~n356 & n5457 ;
  assign n5475 = ~n5059 & n5474 ;
  assign n5476 = ~n5473 & n5475 ;
  assign n5477 = ~n3918 & n5476 ;
  assign n5478 = ( ~n161 & n289 ) | ( ~n161 & n3573 ) | ( n289 & n3573 ) ;
  assign n5479 = n161 | n5478 ;
  assign n5480 = ( n90 & ~n891 ) | ( n90 & n5479 ) | ( ~n891 & n5479 ) ;
  assign n5481 = n891 | n5480 ;
  assign n5482 = n938 | n4008 ;
  assign n5483 = n3043 & ~n3175 ;
  assign n5484 = n2597 | n3568 ;
  assign n5485 = n5483 & ~n5484 ;
  assign n5486 = ~n5482 & n5485 ;
  assign n5487 = ( n2204 & ~n2597 ) | ( n2204 & n5472 ) | ( ~n2597 & n5472 ) ;
  assign n5488 = n2597 | n5487 ;
  assign n5489 = ( ~n591 & n987 ) | ( ~n591 & n5298 ) | ( n987 & n5298 ) ;
  assign n5490 = ~n987 & n5489 ;
  assign n5491 = ( n235 & ~n276 ) | ( n235 & n5490 ) | ( ~n276 & n5490 ) ;
  assign n5492 = ~n235 & n5491 ;
  assign n5493 = ~n759 & n5492 ;
  assign n5494 = ~n356 & n5493 ;
  assign n5495 = ~n3567 & n5494 ;
  assign n5496 = n2098 | n4537 ;
  assign n5497 = ( ~n1630 & n5275 ) | ( ~n1630 & n5496 ) | ( n5275 & n5496 ) ;
  assign n5498 = ~n5447 & n5493 ;
  assign n5499 = n312 | n4810 ;
  assign n5500 = n213 | n4731 ;
  assign n5501 = ( n95 & ~n723 ) | ( n95 & n5500 ) | ( ~n723 & n5500 ) ;
  assign n5502 = n95 | n207 ;
  assign n5503 = ( n1309 & ~n1381 ) | ( n1309 & n5488 ) | ( ~n1381 & n5488 ) ;
  assign n5504 = n1381 | n5503 ;
  assign n5505 = ( n561 & ~n1381 ) | ( n561 & n4027 ) | ( ~n1381 & n4027 ) ;
  assign n5506 = n93 | n5127 ;
  assign n5507 = ( ~n1367 & n4030 ) | ( ~n1367 & n5421 ) | ( n4030 & n5421 ) ;
  assign n5508 = ~n491 & n5477 ;
  assign n5509 = n723 | n5501 ;
  assign n5510 = n3877 | n3901 ;
  assign n5511 = ( ~n90 & n345 ) | ( ~n90 & n5509 ) | ( n345 & n5509 ) ;
  assign n5512 = n90 | n5511 ;
  assign n5513 = n276 | n2098 ;
  assign n5514 = ( ~n1318 & n1367 ) | ( ~n1318 & n5504 ) | ( n1367 & n5504 ) ;
  assign n5515 = n1318 | n5514 ;
  assign n5516 = ( n109 & ~n437 ) | ( n109 & n5515 ) | ( ~n437 & n5515 ) ;
  assign n5517 = n437 | n5516 ;
  assign n5518 = ( ~n304 & n422 ) | ( ~n304 & n5517 ) | ( n422 & n5517 ) ;
  assign n5519 = n304 | n5518 ;
  assign n5520 = ( ~n510 & n1808 ) | ( ~n510 & n5519 ) | ( n1808 & n5519 ) ;
  assign n5521 = n510 | n5520 ;
  assign n5522 = ( ~n1338 & n3877 ) | ( ~n1338 & n5508 ) | ( n3877 & n5508 ) ;
  assign n5523 = n437 | n5081 ;
  assign n5524 = ~n3877 & n5522 ;
  assign n5525 = n1381 | n5505 ;
  assign n5526 = ( n103 & ~n510 ) | ( n103 & n5506 ) | ( ~n510 & n5506 ) ;
  assign n5527 = n302 | n1485 ;
  assign n5528 = n1367 | n5527 ;
  assign n5529 = n5502 | n5528 ;
  assign n5530 = n2008 | n5529 ;
  assign n5531 = n510 | n5526 ;
  assign n5532 = ( ~n276 & n448 ) | ( ~n276 & n5531 ) | ( n448 & n5531 ) ;
  assign n5533 = n2405 | n5513 ;
  assign n5534 = n276 | n5532 ;
  assign n5535 = n4846 | n5513 ;
  assign n5536 = n5499 | n5535 ;
  assign n5537 = n5393 | n5536 ;
  assign n5538 = n5529 | n5533 ;
  assign n5539 = n1367 | n5507 ;
  assign n5540 = n5495 & ~n5530 ;
  assign n5541 = n1246 | n5351 ;
  assign n5542 = ( ~n86 & n2551 ) | ( ~n86 & n5541 ) | ( n2551 & n5541 ) ;
  assign n5543 = n86 | n5542 ;
  assign n5544 = ( n139 & ~n241 ) | ( n139 & n5543 ) | ( ~n241 & n5543 ) ;
  assign n5545 = n241 | n5544 ;
  assign n5546 = ( n188 & ~n232 ) | ( n188 & n5545 ) | ( ~n232 & n5545 ) ;
  assign n5547 = n232 | n5546 ;
  assign n5548 = n410 | n5547 ;
  assign n5549 = n785 | n5548 ;
  assign n5550 = n5538 | n5549 ;
  assign n5551 = ( n957 & ~n2635 ) | ( n957 & n5550 ) | ( ~n2635 & n5550 ) ;
  assign n5552 = n2635 | n5551 ;
  assign n5553 = n148 | n900 ;
  assign n5554 = n289 | n756 ;
  assign n5555 = n5553 | n5554 ;
  assign n5556 = n5412 | n5555 ;
  assign n5557 = ( n203 & ~n489 ) | ( n203 & n5556 ) | ( ~n489 & n5556 ) ;
  assign n5558 = n489 | n5557 ;
  assign n5559 = ( n5312 & ~n5552 ) | ( n5312 & n5558 ) | ( ~n5552 & n5558 ) ;
  assign n5560 = n5552 | n5559 ;
  assign n5561 = ( ~n91 & n290 ) | ( ~n91 & n3646 ) | ( n290 & n3646 ) ;
  assign n5562 = n91 | n5561 ;
  assign n5563 = ( n94 & ~n461 ) | ( n94 & n5562 ) | ( ~n461 & n5562 ) ;
  assign n5564 = n461 | n5563 ;
  assign n5565 = ( ~n145 & n713 ) | ( ~n145 & n5564 ) | ( n713 & n5564 ) ;
  assign n5566 = n145 | n5565 ;
  assign n5567 = n580 | n5566 ;
  assign n5568 = ( ~n3491 & n5510 ) | ( ~n3491 & n5567 ) | ( n5510 & n5567 ) ;
  assign n5569 = n3491 | n5568 ;
  assign n5570 = ( ~n2028 & n3539 ) | ( ~n2028 & n5569 ) | ( n3539 & n5569 ) ;
  assign n5571 = n2028 | n5570 ;
  assign n5572 = ( ~n180 & n1307 ) | ( ~n180 & n4306 ) | ( n1307 & n4306 ) ;
  assign n5573 = n180 | n5572 ;
  assign n5574 = ( ~n94 & n1427 ) | ( ~n94 & n5573 ) | ( n1427 & n5573 ) ;
  assign n5575 = n94 | n5574 ;
  assign n5576 = ( ~n2551 & n3539 ) | ( ~n2551 & n3900 ) | ( n3539 & n3900 ) ;
  assign n5577 = ~n3539 & n5576 ;
  assign n5578 = n2028 | n4825 ;
  assign n5579 = ( ~n1679 & n2551 ) | ( ~n1679 & n5578 ) | ( n2551 & n5578 ) ;
  assign n5580 = ~n2635 & n4889 ;
  assign n5581 = n1630 | n4908 ;
  assign n5582 = ( ~n289 & n5567 ) | ( ~n289 & n5581 ) | ( n5567 & n5581 ) ;
  assign n5583 = n289 | n5582 ;
  assign n5584 = ( n557 & n5331 ) | ( n557 & ~n5558 ) | ( n5331 & ~n5558 ) ;
  assign n5585 = ~n557 & n5584 ;
  assign n5586 = ( ~n145 & n5085 ) | ( ~n145 & n5585 ) | ( n5085 & n5585 ) ;
  assign n5587 = ~n3491 & n5443 ;
  assign n5588 = n2551 | n2657 ;
  assign n5589 = n5587 & ~n5588 ;
  assign n5590 = ~n3690 & n5589 ;
  assign n5591 = ( ~n180 & n5055 ) | ( ~n180 & n5344 ) | ( n5055 & n5344 ) ;
  assign n5592 = n5085 | n5093 ;
  assign n5593 = ~n1146 & n5076 ;
  assign n5594 = ( n125 & ~n241 ) | ( n125 & n5575 ) | ( ~n241 & n5575 ) ;
  assign n5595 = n1679 | n5579 ;
  assign n5596 = ( n602 & ~n790 ) | ( n602 & n5595 ) | ( ~n790 & n5595 ) ;
  assign n5597 = n790 | n5596 ;
  assign n5598 = ( ~n790 & n846 ) | ( ~n790 & n5525 ) | ( n846 & n5525 ) ;
  assign n5599 = n790 | n5598 ;
  assign n5600 = ( ~n116 & n184 ) | ( ~n116 & n5599 ) | ( n184 & n5599 ) ;
  assign n5601 = n116 | n5600 ;
  assign n5602 = ( n88 & ~n89 ) | ( n88 & n5601 ) | ( ~n89 & n5601 ) ;
  assign n5603 = n89 | n5602 ;
  assign n5604 = ( ~n313 & n5421 ) | ( ~n313 & n5537 ) | ( n5421 & n5537 ) ;
  assign n5605 = n313 | n5604 ;
  assign n5606 = ( n296 & ~n592 ) | ( n296 & n5605 ) | ( ~n592 & n5605 ) ;
  assign n5607 = n592 | n5606 ;
  assign n5608 = ( ~n547 & n735 ) | ( ~n547 & n5607 ) | ( n735 & n5607 ) ;
  assign n5609 = n547 | n5608 ;
  assign n5610 = ( n358 & ~n425 ) | ( n358 & n5609 ) | ( ~n425 & n5609 ) ;
  assign n5611 = n425 | n3518 ;
  assign n5612 = n5610 | n5611 ;
  assign n5613 = ( ~n953 & n5603 ) | ( ~n953 & n5612 ) | ( n5603 & n5612 ) ;
  assign n5614 = n953 | n5613 ;
  assign n5615 = ( ~n2611 & n4555 ) | ( ~n2611 & n5614 ) | ( n4555 & n5614 ) ;
  assign n5616 = ( n180 & ~n790 ) | ( n180 & n5255 ) | ( ~n790 & n5255 ) ;
  assign n5617 = ~n180 & n5616 ;
  assign n5618 = ( ~n1354 & n5253 ) | ( ~n1354 & n5421 ) | ( n5253 & n5421 ) ;
  assign n5619 = ~n5421 & n5618 ;
  assign n5620 = ( ~n953 & n5240 ) | ( ~n953 & n5603 ) | ( n5240 & n5603 ) ;
  assign n5621 = n953 | n5620 ;
  assign n5622 = ( n565 & ~n1146 ) | ( n565 & n5621 ) | ( ~n1146 & n5621 ) ;
  assign n5623 = n1146 | n5622 ;
  assign n5624 = n425 | n5610 ;
  assign n5625 = n3167 & ~n5624 ;
  assign n5626 = ~n5085 & n5586 ;
  assign n5627 = ( ~n953 & n3375 ) | ( ~n953 & n5603 ) | ( n3375 & n5603 ) ;
  assign n5628 = ~n5603 & n5627 ;
  assign n5629 = ~n5421 & n5422 ;
  assign n5630 = ( ~n2997 & n5548 ) | ( ~n2997 & n5628 ) | ( n5548 & n5628 ) ;
  assign n5631 = ~n5548 & n5630 ;
  assign n5632 = ( ~n916 & n1679 ) | ( ~n916 & n5592 ) | ( n1679 & n5592 ) ;
  assign n5633 = n916 | n5632 ;
  assign n5634 = n241 | n5594 ;
  assign n5635 = ( ~n82 & n731 ) | ( ~n82 & n5633 ) | ( n731 & n5633 ) ;
  assign n5636 = n82 | n5635 ;
  assign n5637 = ( n293 & ~n423 ) | ( n293 & n5636 ) | ( ~n423 & n5636 ) ;
  assign n5638 = n423 | n5637 ;
  assign n5639 = ( n149 & ~n520 ) | ( n149 & n5638 ) | ( ~n520 & n5638 ) ;
  assign n5640 = n520 | n5639 ;
  assign n5641 = ( n279 & ~n887 ) | ( n279 & n5640 ) | ( ~n887 & n5640 ) ;
  assign n5642 = ( ~n145 & n241 ) | ( ~n145 & n5523 ) | ( n241 & n5523 ) ;
  assign n5643 = n497 | n850 ;
  assign n5644 = n3630 | n5643 ;
  assign n5645 = n612 | n5236 ;
  assign n5646 = n5644 | n5645 ;
  assign n5647 = n87 | n1051 ;
  assign n5648 = n434 | n5647 ;
  assign n5649 = ( n255 & ~n823 ) | ( n255 & n5089 ) | ( ~n823 & n5089 ) ;
  assign n5650 = ( n1056 & ~n2611 ) | ( n1056 & n5229 ) | ( ~n2611 & n5229 ) ;
  assign n5651 = n2611 | n5615 ;
  assign n5652 = ( ~n258 & n293 ) | ( ~n258 & n5539 ) | ( n293 & n5539 ) ;
  assign n5653 = n823 | n5649 ;
  assign n5654 = ( n375 & ~n788 ) | ( n375 & n5653 ) | ( ~n788 & n5653 ) ;
  assign n5655 = n788 | n5654 ;
  assign n5656 = ( n754 & ~n810 ) | ( n754 & n5655 ) | ( ~n810 & n5655 ) ;
  assign n5657 = n810 | n5656 ;
  assign n5658 = ( n187 & ~n833 ) | ( n187 & n5646 ) | ( ~n833 & n5646 ) ;
  assign n5659 = ~n1390 & n3043 ;
  assign n5660 = ~n371 & n5486 ;
  assign n5661 = n203 | n850 ;
  assign n5662 = n833 | n5658 ;
  assign n5663 = n1390 | n5648 ;
  assign n5664 = n4603 | n5641 ;
  assign n5665 = ( n426 & ~n501 ) | ( n426 & n5657 ) | ( ~n501 & n5657 ) ;
  assign n5666 = ( n2829 & ~n2997 ) | ( n2829 & n5664 ) | ( ~n2997 & n5664 ) ;
  assign n5667 = n468 | n559 ;
  assign n5668 = n5663 | n5667 ;
  assign n5669 = n942 | n4172 ;
  assign n5670 = n967 | n5662 ;
  assign n5671 = n2852 | n5668 ;
  assign n5672 = n378 | n5671 ;
  assign n5673 = ~n491 & n5077 ;
  assign n5674 = n589 | n827 ;
  assign n5675 = n5672 | n5674 ;
  assign n5676 = n1398 | n5675 ;
  assign n5677 = n501 | n5665 ;
  assign n5678 = n2997 | n5666 ;
  assign n5679 = ( ~n587 & n5625 ) | ( ~n587 & n5670 ) | ( n5625 & n5670 ) ;
  assign n5680 = ( n1136 & ~n4172 ) | ( n1136 & n5678 ) | ( ~n4172 & n5678 ) ;
  assign n5681 = n4172 | n5680 ;
  assign n5682 = ( ~n1246 & n1307 ) | ( ~n1246 & n5681 ) | ( n1307 & n5681 ) ;
  assign n5683 = n3743 | n5676 ;
  assign n5684 = ~n5648 & n5660 ;
  assign n5685 = n2455 | n5661 ;
  assign n5686 = n5669 | n5685 ;
  assign n5687 = ~n5670 & n5679 ;
  assign n5688 = ( n561 & ~n1308 ) | ( n561 & n5687 ) | ( ~n1308 & n5687 ) ;
  assign n5689 = n3727 | n5683 ;
  assign n5690 = n887 | n5689 ;
  assign n5691 = ( n1309 & n5401 ) | ( n1309 & ~n5677 ) | ( n5401 & ~n5677 ) ;
  assign n5692 = ~n1309 & n5691 ;
  assign n5693 = n5641 | n5690 ;
  assign n5694 = ( n1574 & ~n2455 ) | ( n1574 & n5693 ) | ( ~n2455 & n5693 ) ;
  assign n5695 = ~n2773 & n5684 ;
  assign n5696 = n2455 | n5694 ;
  assign n5697 = ( ~n491 & n2369 ) | ( ~n491 & n5696 ) | ( n2369 & n5696 ) ;
  assign n5698 = n491 | n5697 ;
  assign n5699 = ( n587 & n3950 ) | ( n587 & ~n5677 ) | ( n3950 & ~n5677 ) ;
  assign n5700 = ~n587 & n5699 ;
  assign n5701 = ( ~n3357 & n3650 ) | ( ~n3357 & n5670 ) | ( n3650 & n5670 ) ;
  assign n5702 = ~n4201 & n5695 ;
  assign n5703 = ( n100 & ~n2611 ) | ( n100 & n5673 ) | ( ~n2611 & n5673 ) ;
  assign n5704 = n3357 | n5701 ;
  assign n5705 = ( n1738 & ~n2232 ) | ( n1738 & n5704 ) | ( ~n2232 & n5704 ) ;
  assign n5706 = ~n1738 & n4539 ;
  assign n5707 = ~n5057 & n5659 ;
  assign n5708 = ~n5271 & n5707 ;
  assign n5709 = n644 | n714 ;
  assign n5710 = n1051 | n5416 ;
  assign n5711 = ( ~n1740 & n4847 ) | ( ~n1740 & n5692 ) | ( n4847 & n5692 ) ;
  assign n5712 = ~n4847 & n5711 ;
  assign n5713 = ( ~n731 & n1088 ) | ( ~n731 & n5712 ) | ( n1088 & n5712 ) ;
  assign n5714 = ( n1909 & ~n3491 ) | ( n1909 & n4743 ) | ( ~n3491 & n4743 ) ;
  assign n5715 = ~n1088 & n5713 ;
  assign n5716 = ( ~n2351 & n4743 ) | ( ~n2351 & n5524 ) | ( n4743 & n5524 ) ;
  assign n5717 = ( ~n607 & n4743 ) | ( ~n607 & n5706 ) | ( n4743 & n5706 ) ;
  assign n5718 = ~n4743 & n5716 ;
  assign n5719 = ~n4743 & n5717 ;
  assign n5720 = n546 | n1051 ;
  assign n5721 = ( n234 & ~n757 ) | ( n234 & n5719 ) | ( ~n757 & n5719 ) ;
  assign n5722 = ( ~n82 & n1019 ) | ( ~n82 & n5710 ) | ( n1019 & n5710 ) ;
  assign n5723 = ( ~n1244 & n4520 ) | ( ~n1244 & n5236 ) | ( n4520 & n5236 ) ;
  assign n5724 = n87 | n649 ;
  assign n5725 = n1244 | n5723 ;
  assign n5726 = n5709 | n5724 ;
  assign n5727 = n122 | n345 ;
  assign n5728 = n1135 | n4018 ;
  assign n5729 = n5726 | n5727 ;
  assign n5730 = n434 | n5729 ;
  assign n5731 = n4018 | n5398 ;
  assign n5732 = ( n1246 & ~n2351 ) | ( n1246 & n5404 ) | ( ~n2351 & n5404 ) ;
  assign n5733 = ( ~n1577 & n5631 ) | ( ~n1577 & n5730 ) | ( n5631 & n5730 ) ;
  assign n5734 = ( n3852 & ~n4018 ) | ( n3852 & n5730 ) | ( ~n4018 & n5730 ) ;
  assign n5735 = ~n5730 & n5733 ;
  assign n5736 = ( n3483 & ~n5344 ) | ( n3483 & n5735 ) | ( ~n5344 & n5735 ) ;
  assign n5737 = n4018 | n5734 ;
  assign n5738 = ( n1019 & ~n4288 ) | ( n1019 & n5737 ) | ( ~n4288 & n5737 ) ;
  assign n5739 = ( ~n302 & n1244 ) | ( ~n302 & n5623 ) | ( n1244 & n5623 ) ;
  assign n5740 = ( ~n1095 & n4847 ) | ( ~n1095 & n5400 ) | ( n4847 & n5400 ) ;
  assign n5741 = n757 | n5720 ;
  assign n5742 = n4940 | n5741 ;
  assign n5743 = n4288 | n5738 ;
  assign n5744 = ( n1056 & ~n1244 ) | ( n1056 & n5208 ) | ( ~n1244 & n5208 ) ;
  assign n5745 = ( ~n93 & n423 ) | ( ~n93 & n5743 ) | ( n423 & n5743 ) ;
  assign n5746 = ~n3483 & n5736 ;
  assign n5747 = n93 | n5745 ;
  assign n5748 = ( n3705 & n4694 ) | ( n3705 & ~n5730 ) | ( n4694 & ~n5730 ) ;
  assign n5749 = n1642 | n5742 ;
  assign n5750 = ( ~n213 & n5236 ) | ( ~n213 & n5749 ) | ( n5236 & n5749 ) ;
  assign n5751 = n213 | n5750 ;
  assign n5752 = ~n4694 & n5748 ;
  assign n5753 = ~n4847 & n5752 ;
  assign n5754 = ( n1019 & ~n2942 ) | ( n1019 & n3180 ) | ( ~n2942 & n3180 ) ;
  assign n5755 = ( ~n520 & n2351 ) | ( ~n520 & n5751 ) | ( n2351 & n5751 ) ;
  assign n5756 = ~n2232 & n4682 ;
  assign n5757 = ( ~n92 & n342 ) | ( ~n92 & n4515 ) | ( n342 & n4515 ) ;
  assign n5758 = ( ~n1427 & n2663 ) | ( ~n1427 & n4103 ) | ( n2663 & n4103 ) ;
  assign n5759 = ~n2663 & n5758 ;
  assign n5760 = ( n154 & ~n916 ) | ( n154 & n5759 ) | ( ~n916 & n5759 ) ;
  assign n5761 = n258 | n5652 ;
  assign n5762 = ~n342 & n5757 ;
  assign n5763 = ~n154 & n5760 ;
  assign n5764 = ( ~n258 & n5413 ) | ( ~n258 & n5763 ) | ( n5413 & n5763 ) ;
  assign n5765 = ( ~n258 & n607 ) | ( ~n258 & n5762 ) | ( n607 & n5762 ) ;
  assign n5766 = n235 | n381 ;
  assign n5767 = n5206 | n5766 ;
  assign n5768 = n5728 | n5767 ;
  assign n5769 = n116 | n4873 ;
  assign n5770 = n87 | n373 ;
  assign n5771 = n3090 | n5770 ;
  assign n5772 = n552 | n721 ;
  assign n5773 = ~n116 & n5360 ;
  assign n5774 = ( ~n92 & n103 ) | ( ~n92 & n5731 ) | ( n103 & n5731 ) ;
  assign n5775 = ( ~n92 & n344 ) | ( ~n92 & n5756 ) | ( n344 & n5756 ) ;
  assign n5776 = ~n2030 & n5461 ;
  assign n5777 = ( ~n98 & n2942 ) | ( ~n98 & n5718 ) | ( n2942 & n5718 ) ;
  assign n5778 = ~n607 & n5765 ;
  assign n5779 = n92 | n5774 ;
  assign n5780 = n1446 | n5768 ;
  assign n5781 = ~n2942 & n5777 ;
  assign n5782 = ~n344 & n5775 ;
  assign n5783 = ~n5413 & n5764 ;
  assign n5784 = ( n344 & n5307 ) | ( n344 & ~n5344 ) | ( n5307 & ~n5344 ) ;
  assign n5785 = ( n165 & ~n342 ) | ( n165 & n5781 ) | ( ~n342 & n5781 ) ;
  assign n5786 = n5771 | n5772 ;
  assign n5787 = ( n378 & ~n945 ) | ( n378 & n5786 ) | ( ~n945 & n5786 ) ;
  assign n5788 = n945 | n5787 ;
  assign n5789 = n425 | n5788 ;
  assign n5790 = n2650 | n5789 ;
  assign n5791 = n4675 & ~n5790 ;
  assign n5792 = ~n5780 & n5791 ;
  assign n5793 = ~n4072 & n5792 ;
  assign n5794 = ( ~n1427 & n2030 ) | ( ~n1427 & n5793 ) | ( n2030 & n5793 ) ;
  assign n5795 = ~n2030 & n5794 ;
  assign n5796 = ( ~n282 & n546 ) | ( ~n282 & n5795 ) | ( n546 & n5795 ) ;
  assign n5797 = ( ~n116 & n825 ) | ( ~n116 & n5776 ) | ( n825 & n5776 ) ;
  assign n5798 = n1095 | n5740 ;
  assign n5799 = ( n501 & ~n580 ) | ( n501 & n5481 ) | ( ~n580 & n5481 ) ;
  assign n5800 = n580 | n5799 ;
  assign n5801 = ( n306 & ~n1384 ) | ( n306 & n5798 ) | ( ~n1384 & n5798 ) ;
  assign n5802 = n1384 | n5801 ;
  assign n5803 = ( ~n153 & n693 ) | ( ~n153 & n5802 ) | ( n693 & n5802 ) ;
  assign n5804 = n153 | n5803 ;
  assign n5805 = ( ~n522 & n534 ) | ( ~n522 & n5634 ) | ( n534 & n5634 ) ;
  assign n5806 = n124 | n589 ;
  assign n5807 = ( ~n361 & n1318 ) | ( ~n361 & n3843 ) | ( n1318 & n3843 ) ;
  assign n5808 = ~n2232 & n3709 ;
  assign n5809 = ( n161 & ~n1520 ) | ( n161 & n5560 ) | ( ~n1520 & n5560 ) ;
  assign n5810 = ~n3266 & n5808 ;
  assign n5811 = n1427 | n3266 ;
  assign n5812 = n647 | n702 ;
  assign n5813 = ( ~n1427 & n2795 ) | ( ~n1427 & n4938 ) | ( n2795 & n4938 ) ;
  assign n5814 = n1427 | n5813 ;
  assign n5815 = n756 | n778 ;
  assign n5816 = n5806 | n5815 ;
  assign n5817 = n5741 | n5812 ;
  assign n5818 = n4179 | n5816 ;
  assign n5819 = n600 | n759 ;
  assign n5820 = n532 | n559 ;
  assign n5821 = n107 | n5800 ;
  assign n5822 = ( n122 & ~n701 ) | ( n122 & n5818 ) | ( ~n701 & n5818 ) ;
  assign n5823 = n5819 | n5820 ;
  assign n5824 = n5817 | n5823 ;
  assign n5825 = ( ~n234 & n283 ) | ( ~n234 & n5583 ) | ( n283 & n5583 ) ;
  assign n5826 = n361 | n5807 ;
  assign n5827 = n182 | n5824 ;
  assign n5828 = n3491 | n5714 ;
  assign n5829 = ( n1095 & ~n2266 ) | ( n1095 & n5580 ) | ( ~n2266 & n5580 ) ;
  assign n5830 = n2431 | n5827 ;
  assign n5831 = ~n1095 & n5829 ;
  assign n5832 = ( ~n306 & n373 ) | ( ~n306 & n5831 ) | ( n373 & n5831 ) ;
  assign n5833 = n1520 | n5809 ;
  assign n5834 = ( n2909 & ~n3491 ) | ( n2909 & n5826 ) | ( ~n3491 & n5826 ) ;
  assign n5835 = n234 | n5825 ;
  assign n5836 = ( ~n86 & n823 ) | ( ~n86 & n5828 ) | ( n823 & n5828 ) ;
  assign n5837 = ~n373 & n5832 ;
  assign n5838 = n3491 | n5834 ;
  assign n5839 = n701 | n5822 ;
  assign n5840 = n963 | n5839 ;
  assign n5841 = n522 | n5805 ;
  assign n5842 = n1169 | n1195 ;
  assign n5843 = n5225 | n5840 ;
  assign n5844 = n5513 | n5821 ;
  assign n5845 = n303 | n1520 ;
  assign n5846 = n5842 | n5843 ;
  assign n5847 = ( n234 & ~n823 ) | ( n234 & n5698 ) | ( ~n823 & n5698 ) ;
  assign n5848 = n823 | n5847 ;
  assign n5849 = ( n229 & ~n823 ) | ( n229 & n4729 ) | ( ~n823 & n4729 ) ;
  assign n5850 = n1275 | n5768 ;
  assign n5851 = n373 | n5848 ;
  assign n5852 = ( n4168 & n5192 ) | ( n4168 & ~n5841 ) | ( n5192 & ~n5841 ) ;
  assign n5853 = n5811 | n5845 ;
  assign n5854 = ~n5192 & n5852 ;
  assign n5855 = n5789 | n5821 ;
  assign n5856 = n5846 | n5855 ;
  assign n5857 = ( ~n1630 & n5841 ) | ( ~n1630 & n5856 ) | ( n5841 & n5856 ) ;
  assign n5858 = n1630 | n5857 ;
  assign n5859 = n1095 | n5328 ;
  assign n5860 = n361 | n2098 ;
  assign n5861 = ~n234 & n5721 ;
  assign n5862 = n5686 | n5860 ;
  assign n5863 = n4683 | n5853 ;
  assign n5864 = n5830 | n5844 ;
  assign n5865 = n5850 | n5864 ;
  assign n5866 = ( ~n1740 & n5841 ) | ( ~n1740 & n5865 ) | ( n5841 & n5865 ) ;
  assign n5867 = n1992 | n5840 ;
  assign n5868 = n5862 | n5867 ;
  assign n5869 = ( ~n209 & n1095 ) | ( ~n209 & n5868 ) | ( n1095 & n5868 ) ;
  assign n5870 = ( ~n987 & n2795 ) | ( ~n987 & n5858 ) | ( n2795 & n5858 ) ;
  assign n5871 = n987 | n5870 ;
  assign n5872 = n1740 | n5866 ;
  assign n5873 = ( n532 & ~n1630 ) | ( n532 & n4932 ) | ( ~n1630 & n4932 ) ;
  assign n5874 = ( ~n182 & n426 ) | ( ~n182 & n4592 ) | ( n426 & n4592 ) ;
  assign n5875 = n182 | n5874 ;
  assign n5876 = ( n832 & ~n872 ) | ( n832 & n5875 ) | ( ~n872 & n5875 ) ;
  assign n5877 = ( n561 & ~n2663 ) | ( n561 & n5343 ) | ( ~n2663 & n5343 ) ;
  assign n5878 = ~n561 & n5688 ;
  assign n5879 = n872 | n5876 ;
  assign n5880 = n5702 & ~n5768 ;
  assign n5881 = n1577 | n5812 ;
  assign n5882 = ( n312 & ~n5879 ) | ( n312 & n5880 ) | ( ~n5879 & n5880 ) ;
  assign n5883 = ( ~n578 & n955 ) | ( ~n578 & n5593 ) | ( n955 & n5593 ) ;
  assign n5884 = ( ~n1318 & n2909 ) | ( ~n1318 & n4329 ) | ( n2909 & n4329 ) ;
  assign n5885 = ( n213 & ~n1630 ) | ( n213 & n5069 ) | ( ~n1630 & n5069 ) ;
  assign n5886 = ~n1246 & n5732 ;
  assign n5887 = ( ~n302 & n313 ) | ( ~n302 & n5886 ) | ( n313 & n5886 ) ;
  assign n5888 = ~n313 & n5887 ;
  assign n5889 = ( n1338 & ~n1630 ) | ( n1338 & n5708 ) | ( ~n1630 & n5708 ) ;
  assign n5890 = ~n381 & n583 ;
  assign n5891 = ~n1512 & n5890 ;
  assign n5892 = n1630 | n5339 ;
  assign n5893 = n1630 | n5497 ;
  assign n5894 = ~n312 & n5882 ;
  assign n5895 = n938 | n5879 ;
  assign n5896 = n5675 | n5879 ;
  assign n5897 = n371 | n5881 ;
  assign n5898 = n2191 | n5897 ;
  assign n5899 = n5057 | n5898 ;
  assign n5900 = n3748 | n5899 ;
  assign n5901 = ( n938 & n5768 ) | ( n938 & ~n5900 ) | ( n5768 & ~n5900 ) ;
  assign n5902 = ( n1051 & ~n3568 ) | ( n1051 & n5408 ) | ( ~n3568 & n5408 ) ;
  assign n5903 = n5900 | n5901 ;
  assign n5904 = n3568 | n5902 ;
  assign n5905 = ( n1338 & ~n2266 ) | ( n1338 & n5125 ) | ( ~n2266 & n5125 ) ;
  assign n5906 = ( ~n91 & n561 ) | ( ~n91 & n5892 ) | ( n561 & n5892 ) ;
  assign n5907 = ~n955 & n5883 ;
  assign n5908 = ~n1390 & n5891 ;
  assign n5909 = n717 | n963 ;
  assign n5910 = n5686 | n5909 ;
  assign n5911 = ~n1338 & n5889 ;
  assign n5912 = n777 | n1195 ;
  assign n5913 = n5896 | n5910 ;
  assign n5914 = n5908 & ~n5912 ;
  assign n5915 = ( ~n86 & n2657 ) | ( ~n86 & n5904 ) | ( n2657 & n5904 ) ;
  assign n5916 = ( ~n1837 & n2657 ) | ( ~n1837 & n5893 ) | ( n2657 & n5893 ) ;
  assign n5917 = ( ~n279 & n2098 ) | ( ~n279 & n5903 ) | ( n2098 & n5903 ) ;
  assign n5918 = n4282 | n5913 ;
  assign n5919 = n213 | n1663 ;
  assign n5920 = ~n1663 & n5891 ;
  assign n5921 = ~n5898 & n5920 ;
  assign n5922 = n2191 | n5293 ;
  assign n5923 = n1159 | n4967 ;
  assign n5924 = n1318 | n5884 ;
  assign n5925 = n1837 | n5916 ;
  assign n5926 = ( n125 & ~n228 ) | ( n125 & n5577 ) | ( ~n228 & n5577 ) ;
  assign n5927 = ~n125 & n5926 ;
  assign n5928 = n1318 | n5881 ;
  assign n5929 = n5014 | n5919 ;
  assign n5930 = ~n4056 & n5914 ;
  assign n5931 = ~n1159 & n5930 ;
  assign n5932 = n381 | n1512 ;
  assign n5933 = n1338 | n5034 ;
  assign n5934 = ( ~n82 & n4999 ) | ( ~n82 & n5924 ) | ( n4999 & n5924 ) ;
  assign n5935 = ( n423 & ~n534 ) | ( n423 & n5927 ) | ( ~n534 & n5927 ) ;
  assign n5936 = ~n2098 & n5931 ;
  assign n5937 = ( n701 & ~n759 ) | ( n701 & n5907 ) | ( ~n759 & n5907 ) ;
  assign n5938 = n5928 | n5929 ;
  assign n5939 = n1630 | n5885 ;
  assign n5940 = n5922 | n5932 ;
  assign n5941 = ~n5918 & n5921 ;
  assign n5942 = ( n213 & ~n4999 ) | ( n213 & n5911 ) | ( ~n4999 & n5911 ) ;
  assign n5943 = ( ~n82 & n341 ) | ( ~n82 & n5925 ) | ( n341 & n5925 ) ;
  assign n5944 = ( ~n91 & n165 ) | ( ~n91 & n5446 ) | ( n165 & n5446 ) ;
  assign n5945 = n2663 | n5877 ;
  assign n5946 = n235 | n5827 ;
  assign n5947 = n2549 | n4935 ;
  assign n5948 = ( ~n167 & n593 ) | ( ~n167 & n5347 ) | ( n593 & n5347 ) ;
  assign n5949 = ~n165 & n5944 ;
  assign n5950 = ( n345 & ~n461 ) | ( n345 & n5949 ) | ( ~n461 & n5949 ) ;
  assign n5951 = ~n345 & n5950 ;
  assign n5952 = ( n497 & ~n715 ) | ( n497 & n5951 ) | ( ~n715 & n5951 ) ;
  assign n5953 = ~n497 & n5952 ;
  assign n5954 = ~n165 & n5785 ;
  assign n5955 = ~n2549 & n4808 ;
  assign n5956 = ( ~n165 & n300 ) | ( ~n165 & n5619 ) | ( n300 & n5619 ) ;
  assign n5957 = ( ~n501 & n832 ) | ( ~n501 & n5953 ) | ( n832 & n5953 ) ;
  assign n5958 = ( n2446 & ~n2663 ) | ( n2446 & n5936 ) | ( ~n2663 & n5936 ) ;
  assign n5959 = ( n229 & ~n2663 ) | ( n229 & n5894 ) | ( ~n2663 & n5894 ) ;
  assign n5960 = ~n832 & n5957 ;
  assign n5961 = ~n147 & n5660 ;
  assign n5962 = n340 | n744 ;
  assign n5963 = ~n5206 & n5961 ;
  assign n5964 = ~n5962 & n5963 ;
  assign n5965 = ~n102 & n5964 ;
  assign n5966 = ( ~n522 & n602 ) | ( ~n522 & n5833 ) | ( n602 & n5833 ) ;
  assign n5967 = n228 | n5812 ;
  assign n5968 = n1051 | n4765 ;
  assign n5969 = ( ~n287 & n1485 ) | ( ~n287 & n5939 ) | ( n1485 & n5939 ) ;
  assign n5970 = n5965 & ~n5967 ;
  assign n5971 = n1974 | n5293 ;
  assign n5972 = n433 | n522 ;
  assign n5973 = n209 | n5869 ;
  assign n5974 = n448 | n5972 ;
  assign n5975 = n522 | n5966 ;
  assign n5976 = n1195 | n5973 ;
  assign n5977 = n612 | n658 ;
  assign n5978 = n5970 & ~n5971 ;
  assign n5979 = n287 | n5969 ;
  assign n5980 = ( n653 & ~n849 ) | ( n653 & n5979 ) | ( ~n849 & n5979 ) ;
  assign n5981 = n5974 | n5977 ;
  assign n5982 = n960 | n5981 ;
  assign n5983 = n849 | n5980 ;
  assign n5984 = ~n1354 & n5330 ;
  assign n5985 = n5973 | n5981 ;
  assign n5986 = n1349 | n4302 ;
  assign n5987 = ( ~n343 & n3428 ) | ( ~n343 & n5983 ) | ( n3428 & n5983 ) ;
  assign n5988 = n343 | n5987 ;
  assign n5989 = n5940 | n5982 ;
  assign n5990 = n4670 | n5989 ;
  assign n5991 = n2871 | n5990 ;
  assign n5992 = ( ~n1354 & n4654 ) | ( ~n1354 & n5988 ) | ( n4654 & n5988 ) ;
  assign n5993 = n343 | n5983 ;
  assign n5994 = ( ~n777 & n5991 ) | ( ~n777 & n5993 ) | ( n5991 & n5993 ) ;
  assign n5995 = n777 | n5994 ;
  assign n5996 = ( n948 & ~n2613 ) | ( n948 & n5995 ) | ( ~n2613 & n5995 ) ;
  assign n5997 = n2613 | n5996 ;
  assign n5998 = ~n1349 & n5964 ;
  assign n5999 = ( n1136 & ~n2549 ) | ( n1136 & n5997 ) | ( ~n2549 & n5997 ) ;
  assign n6000 = n1354 | n5992 ;
  assign n6001 = ( ~n1051 & n2663 ) | ( ~n1051 & n6000 ) | ( n2663 & n6000 ) ;
  assign n6002 = n2549 | n5999 ;
  assign n6003 = ~n5946 & n5998 ;
  assign n6004 = ~n5985 & n6003 ;
  assign n6005 = ( n2329 & ~n3568 ) | ( n2329 & n6002 ) | ( ~n3568 & n6002 ) ;
  assign n6006 = n3568 | n6005 ;
  assign n6007 = n1051 | n6001 ;
  assign n6008 = ( ~n154 & n497 ) | ( ~n154 & n6006 ) | ( n497 & n6006 ) ;
  assign n6009 = ( n367 & ~n655 ) | ( n367 & n5512 ) | ( ~n655 & n5512 ) ;
  assign n6010 = ( ~n585 & n1056 ) | ( ~n585 & n5968 ) | ( n1056 & n5968 ) ;
  assign n6011 = n585 | n6010 ;
  assign n6012 = ( n235 & ~n643 ) | ( n235 & n6011 ) | ( ~n643 & n6011 ) ;
  assign n6013 = n91 | n5906 ;
  assign n6014 = ( n214 & ~n228 ) | ( n214 & n6013 ) | ( ~n228 & n6013 ) ;
  assign n6015 = ~n1056 & n5650 ;
  assign n6016 = ( n345 & ~n731 ) | ( n345 & n5571 ) | ( ~n731 & n5571 ) ;
  assign n6017 = n125 | n3248 ;
  assign n6018 = ~n1679 & n5810 ;
  assign n6019 = ~n2329 & n6018 ;
  assign n6020 = n82 | n5934 ;
  assign n6021 = ( n149 & ~n702 ) | ( n149 & n6020 ) | ( ~n702 & n6020 ) ;
  assign n6022 = n702 | n6021 ;
  assign n6023 = ( n358 & ~n378 ) | ( n358 & n6022 ) | ( ~n378 & n6022 ) ;
  assign n6024 = ( ~n91 & n2795 ) | ( ~n91 & n4540 ) | ( n2795 & n4540 ) ;
  assign n6025 = n91 | n6024 ;
  assign n6026 = ( ~n318 & n415 ) | ( ~n318 & n6025 ) | ( n415 & n6025 ) ;
  assign n6027 = n318 | n6026 ;
  assign n6028 = ( ~n89 & n5016 ) | ( ~n89 & n6027 ) | ( n5016 & n6027 ) ;
  assign n6029 = ( n101 & ~n125 ) | ( n101 & n5954 ) | ( ~n125 & n5954 ) ;
  assign n6030 = ( ~n916 & n1056 ) | ( ~n916 & n5700 ) | ( n1056 & n5700 ) ;
  assign n6031 = ~n1056 & n6030 ;
  assign n6032 = ( ~n82 & n602 ) | ( ~n82 & n6031 ) | ( n602 & n6031 ) ;
  assign n6033 = ~n602 & n6032 ;
  assign n6034 = ( n583 & n744 ) | ( n583 & ~n5938 ) | ( n744 & ~n5938 ) ;
  assign n6035 = ~n744 & n6034 ;
  assign n6036 = ( n235 & ~n754 ) | ( n235 & n5814 ) | ( ~n754 & n5814 ) ;
  assign n6037 = n2329 | n3509 ;
  assign n6038 = n417 | n5359 ;
  assign n6039 = ( ~n102 & n345 ) | ( ~n102 & n6038 ) | ( n345 & n6038 ) ;
  assign n6040 = ( n247 & ~n422 ) | ( n247 & n5280 ) | ( ~n422 & n5280 ) ;
  assign n6041 = n422 | n6040 ;
  assign n6042 = n222 | n6041 ;
  assign n6043 = ( n2266 & ~n2446 ) | ( n2266 & n4915 ) | ( ~n2446 & n4915 ) ;
  assign n6044 = n2446 | n6043 ;
  assign n6045 = ( ~n91 & n2246 ) | ( ~n91 & n6044 ) | ( n2246 & n6044 ) ;
  assign n6046 = n91 | n6045 ;
  assign n6047 = ( ~n367 & n578 ) | ( ~n367 & n5783 ) | ( n578 & n5783 ) ;
  assign n6048 = n82 | n5943 ;
  assign n6049 = n82 | n5722 ;
  assign n6050 = ( ~n367 & n422 ) | ( ~n367 & n6049 ) | ( n422 & n6049 ) ;
  assign n6051 = n367 | n6050 ;
  assign n6052 = n302 | n5739 ;
  assign n6053 = ( ~n162 & n214 ) | ( ~n162 & n6052 ) | ( n214 & n6052 ) ;
  assign n6054 = ( n3963 & ~n5344 ) | ( n3963 & n5854 ) | ( ~n5344 & n5854 ) ;
  assign n6055 = ~n3963 & n6054 ;
  assign n6056 = ( ~n283 & n1837 ) | ( ~n283 & n4761 ) | ( n1837 & n4761 ) ;
  assign n6057 = n283 | n6056 ;
  assign n6058 = ( n290 & ~n415 ) | ( n290 & n6057 ) | ( ~n415 & n6057 ) ;
  assign n6059 = n415 | n6058 ;
  assign n6060 = ( ~n145 & n222 ) | ( ~n145 & n6059 ) | ( n222 & n6059 ) ;
  assign n6061 = ~n1056 & n5744 ;
  assign n6062 = n1974 | n5989 ;
  assign n6063 = ~n5672 & n6035 ;
  assign n6064 = ~n5895 & n6063 ;
  assign n6065 = ~n6062 & n6064 ;
  assign n6066 = ~n2246 & n4219 ;
  assign n6067 = ( ~n296 & n879 ) | ( ~n296 & n5955 ) | ( n879 & n5955 ) ;
  assign n6068 = ~n879 & n6067 ;
  assign n6069 = n2446 | n5281 ;
  assign n6070 = ( n81 & ~n286 ) | ( n81 & n6069 ) | ( ~n286 & n6069 ) ;
  assign n6071 = n286 | n6070 ;
  assign n6072 = n1246 | n5682 ;
  assign n6073 = ( ~n693 & n1384 ) | ( ~n693 & n6072 ) | ( n1384 & n6072 ) ;
  assign n6074 = ( n303 & ~n503 ) | ( n303 & n5871 ) | ( ~n503 & n5871 ) ;
  assign n6075 = ~n2942 & n4588 ;
  assign n6076 = ~n1246 & n6075 ;
  assign n6077 = ( n303 & ~n605 ) | ( n303 & n6076 ) | ( ~n605 & n6076 ) ;
  assign n6078 = ~n303 & n6077 ;
  assign n6079 = n286 | n4858 ;
  assign n6080 = ( n169 & ~n592 ) | ( n169 & n5863 ) | ( ~n592 & n5863 ) ;
  assign n6081 = n592 | n6080 ;
  assign n6082 = ( n172 & ~n420 ) | ( n172 & n6081 ) | ( ~n420 & n6081 ) ;
  assign n6083 = n420 | n6082 ;
  assign n6084 = ( n148 & ~n559 ) | ( n148 & n6083 ) | ( ~n559 & n6083 ) ;
  assign n6085 = n559 | n6084 ;
  assign n6086 = ( ~n161 & n1837 ) | ( ~n161 & n2737 ) | ( n1837 & n2737 ) ;
  assign n6087 = n161 | n6086 ;
  assign n6088 = ( n786 & ~n829 ) | ( n786 & n6087 ) | ( ~n829 & n6087 ) ;
  assign n6089 = n829 | n6088 ;
  assign n6090 = ( ~n168 & n188 ) | ( ~n168 & n6089 ) | ( n188 & n6089 ) ;
  assign n6091 = n168 | n6090 ;
  assign n6092 = ( n219 & ~n655 ) | ( n219 & n6091 ) | ( ~n655 & n6091 ) ;
  assign n6093 = n655 | n6092 ;
  assign n6094 = ( n5540 & n6085 ) | ( n5540 & ~n6093 ) | ( n6085 & ~n6093 ) ;
  assign n6095 = ~n6085 & n6094 ;
  assign n6096 = ( n879 & ~n1384 ) | ( n879 & n6095 ) | ( ~n1384 & n6095 ) ;
  assign n6097 = ~n879 & n6096 ;
  assign n6098 = ( n2246 & ~n2942 ) | ( n2246 & n6097 ) | ( ~n2942 & n6097 ) ;
  assign n6099 = ~n2246 & n6098 ;
  assign n6100 = ~n5153 & n6099 ;
  assign n6101 = ~n5095 & n6100 ;
  assign n6102 = ( ~n650 & n955 ) | ( ~n650 & n6101 ) | ( n955 & n6101 ) ;
  assign n6103 = ( ~n2909 & n5984 ) | ( ~n2909 & n6093 ) | ( n5984 & n6093 ) ;
  assign n6104 = ~n6093 & n6103 ;
  assign n6105 = ( ~n1246 & n2909 ) | ( ~n1246 & n5258 ) | ( n2909 & n5258 ) ;
  assign n6106 = ~n2909 & n6105 ;
  assign n6107 = ( ~n693 & n6007 ) | ( ~n693 & n6093 ) | ( n6007 & n6093 ) ;
  assign n6108 = ( ~n81 & n2246 ) | ( ~n81 & n3315 ) | ( n2246 & n3315 ) ;
  assign n6109 = n81 | n6108 ;
  assign n6110 = ( ~n302 & n879 ) | ( ~n302 & n5986 ) | ( n879 & n5986 ) ;
  assign n6111 = ( ~n1246 & n2232 ) | ( ~n1246 & n4353 ) | ( n2232 & n4353 ) ;
  assign n6112 = ( ~n2795 & n5725 ) | ( ~n2795 & n6085 ) | ( n5725 & n6085 ) ;
  assign n6113 = n2942 | n5754 ;
  assign n6114 = ( n81 & ~n86 ) | ( n81 & n6113 ) | ( ~n86 & n6113 ) ;
  assign n6115 = n5344 | n5784 ;
  assign n6116 = ~n5344 & n5591 ;
  assign n6117 = ( ~n294 & n296 ) | ( ~n294 & n6116 ) | ( n296 & n6116 ) ;
  assign n6118 = ~n296 & n6117 ;
  assign n6119 = ( ~n420 & n960 ) | ( ~n420 & n6118 ) | ( n960 & n6118 ) ;
  assign n6120 = ( ~n296 & n2446 ) | ( ~n296 & n4443 ) | ( n2446 & n4443 ) ;
  assign n6121 = ~n2232 & n5460 ;
  assign n6122 = ( ~n287 & n2266 ) | ( ~n287 & n6121 ) | ( n2266 & n6121 ) ;
  assign n6123 = ~n2266 & n6122 ;
  assign n6124 = ( ~n318 & n923 ) | ( ~n318 & n6123 ) | ( n923 & n6123 ) ;
  assign n6125 = ~n923 & n6124 ;
  assign n6126 = ( n103 & ~n461 ) | ( n103 & n6125 ) | ( ~n461 & n6125 ) ;
  assign n6127 = n693 | n6073 ;
  assign n6128 = ( ~n693 & n943 ) | ( ~n693 & n4809 ) | ( n943 & n4809 ) ;
  assign n6129 = ( ~n98 & n490 ) | ( ~n98 & n5366 ) | ( n490 & n5366 ) ;
  assign n6130 = n98 | n6129 ;
  assign n6131 = ( n96 & ~n294 ) | ( n96 & n6130 ) | ( ~n294 & n6130 ) ;
  assign n6132 = n294 | n6131 ;
  assign n6133 = ( n585 & ~n846 ) | ( n585 & n6132 ) | ( ~n846 & n6132 ) ;
  assign n6134 = n846 | n6133 ;
  assign n6135 = ( n139 & ~n694 ) | ( n139 & n6134 ) | ( ~n694 & n6134 ) ;
  assign n6136 = ( n585 & ~n887 ) | ( n585 & n6079 ) | ( ~n887 & n6079 ) ;
  assign n6137 = ( n139 & ~n173 ) | ( n139 & n5651 ) | ( ~n173 & n5651 ) ;
  assign n6138 = ( ~n98 & n109 ) | ( ~n98 & n5414 ) | ( n109 & n5414 ) ;
  assign n6139 = n2232 | n5705 ;
  assign n6140 = ( ~n731 & n5344 ) | ( ~n731 & n6139 ) | ( n5344 & n6139 ) ;
  assign n6141 = ( n154 & ~n294 ) | ( n154 & n6104 ) | ( ~n294 & n6104 ) ;
  assign n6142 = ~n154 & n6141 ;
  assign n6143 = ( ~n98 & n290 ) | ( ~n98 & n6106 ) | ( n290 & n6106 ) ;
  assign n6144 = ( ~n362 & n2795 ) | ( ~n362 & n5941 ) | ( n2795 & n5941 ) ;
  assign n6145 = ~n2795 & n6144 ;
  assign n6146 = n693 | n6107 ;
  assign n6147 = n2266 | n5905 ;
  assign n6148 = ( n149 & ~n420 ) | ( n149 & n5837 ) | ( ~n420 & n5837 ) ;
  assign n6149 = ~n149 & n6148 ;
  assign n6150 = ~n2232 & n6111 ;
  assign n6151 = n2795 | n6112 ;
  assign n6152 = ( ~n86 & n294 ) | ( ~n86 & n6151 ) | ( n294 & n6151 ) ;
  assign n6153 = ( ~n103 & n139 ) | ( ~n103 & n5333 ) | ( n139 & n5333 ) ;
  assign n6154 = ( n229 & ~n461 ) | ( n229 & n6061 ) | ( ~n461 & n6061 ) ;
  assign n6155 = ( ~n296 & n304 ) | ( ~n296 & n4881 ) | ( n304 & n4881 ) ;
  assign n6156 = ~n304 & n6155 ;
  assign n6157 = ( n149 & ~n923 ) | ( n149 & n6156 ) | ( ~n923 & n6156 ) ;
  assign n6158 = ~n149 & n6157 ;
  assign n6159 = ( n101 & ~n294 ) | ( n101 & n5590 ) | ( ~n294 & n5590 ) ;
  assign n6160 = ( n154 & ~n296 ) | ( n154 & n5746 ) | ( ~n296 & n5746 ) ;
  assign n6161 = ~n154 & n6160 ;
  assign n6162 = n154 | n6008 ;
  assign n6163 = n86 | n5836 ;
  assign n6164 = ( ~n447 & n965 ) | ( ~n447 & n6163 ) | ( n965 & n6163 ) ;
  assign n6165 = ( n287 & ~n965 ) | ( n287 & n6066 ) | ( ~n965 & n6066 ) ;
  assign n6166 = ( n332 & ~n592 ) | ( n332 & n6068 ) | ( ~n592 & n6068 ) ;
  assign n6167 = ~n332 & n6166 ;
  assign n6168 = ( n503 & ~n605 ) | ( n503 & n6167 ) | ( ~n605 & n6167 ) ;
  assign n6169 = ~n503 & n6168 ;
  assign n6170 = ~n778 & n6169 ;
  assign n6171 = ( ~n779 & n2227 ) | ( ~n779 & n5933 ) | ( n2227 & n5933 ) ;
  assign n6172 = ~n2446 & n6120 ;
  assign n6173 = ~n2446 & n5753 ;
  assign n6174 = ( ~n916 & n2227 ) | ( ~n916 & n3371 ) | ( n2227 & n3371 ) ;
  assign n6175 = ~n2227 & n6174 ;
  assign n6176 = ( ~n109 & n150 ) | ( ~n109 & n6175 ) | ( n150 & n6175 ) ;
  assign n6177 = ~n150 & n6176 ;
  assign n6178 = ( ~n145 & n643 ) | ( ~n145 & n6033 ) | ( n643 & n6033 ) ;
  assign n6179 = ~n643 & n6178 ;
  assign n6180 = ( n89 & ~n841 ) | ( n89 & n6179 ) | ( ~n841 & n6179 ) ;
  assign n6181 = n503 | n6074 ;
  assign n6182 = ~n2446 & n5958 ;
  assign n6183 = ( n172 & ~n283 ) | ( n172 & n6182 ) | ( ~n283 & n6182 ) ;
  assign n6184 = ( n255 & ~n503 ) | ( n255 & n6037 ) | ( ~n503 & n6037 ) ;
  assign n6185 = n503 | n6184 ;
  assign n6186 = ( ~n96 & n150 ) | ( ~n96 & n4827 ) | ( n150 & n4827 ) ;
  assign n6187 = ~n109 & n6138 ;
  assign n6188 = ( n124 & ~n255 ) | ( n124 & n6187 ) | ( ~n255 & n6187 ) ;
  assign n6189 = ( ~n592 & n2227 ) | ( ~n592 & n5838 ) | ( n2227 & n5838 ) ;
  assign n6190 = n592 | n6189 ;
  assign n6191 = ( ~n592 & n1679 ) | ( ~n592 & n6147 ) | ( n1679 & n6147 ) ;
  assign n6192 = n592 | n6191 ;
  assign n6193 = ( ~n168 & n520 ) | ( ~n168 & n6192 ) | ( n520 & n6192 ) ;
  assign n6194 = n168 | n6193 ;
  assign n6195 = ( n109 & ~n714 ) | ( n109 & n5782 ) | ( ~n714 & n5782 ) ;
  assign n6196 = ~n109 & n6195 ;
  assign n6197 = ( ~n255 & n349 ) | ( ~n255 & n2703 ) | ( n349 & n2703 ) ;
  assign n6198 = n255 | n6197 ;
  assign n6199 = ~n2446 & n5498 ;
  assign n6200 = ~n213 & n5942 ;
  assign n6201 = ( ~n283 & n332 ) | ( ~n283 & n6200 ) | ( n332 & n6200 ) ;
  assign n6202 = ~n332 & n6201 ;
  assign n6203 = ( ~n644 & n969 ) | ( ~n644 & n1803 ) | ( n969 & n1803 ) ;
  assign n6204 = n644 | n6203 ;
  assign n6205 = ( n101 & ~n825 ) | ( n101 & n6172 ) | ( ~n825 & n6172 ) ;
  assign n6206 = ~n101 & n6205 ;
  assign n6207 = ( ~n887 & n4444 ) | ( ~n887 & n6206 ) | ( n4444 & n6206 ) ;
  assign n6208 = ~n4444 & n6207 ;
  assign n6209 = ~n103 & n6126 ;
  assign n6210 = n372 | n5264 ;
  assign n6211 = ( ~n173 & n502 ) | ( ~n173 & n6017 ) | ( n502 & n6017 ) ;
  assign n6212 = n173 | n6211 ;
  assign n6213 = ( ~n605 & n887 ) | ( ~n605 & n6212 ) | ( n887 & n6212 ) ;
  assign n6214 = n605 | n6213 ;
  assign n6215 = ( n89 & ~n715 ) | ( n89 & n6214 ) | ( ~n715 & n6214 ) ;
  assign n6216 = n715 | n6215 ;
  assign n6217 = ( n578 & ~n872 ) | ( n578 & n6216 ) | ( ~n872 & n6216 ) ;
  assign n6218 = n872 | n6217 ;
  assign n6219 = n5338 & ~n6218 ;
  assign n6220 = ~n6210 & n6219 ;
  assign n6221 = ( ~n499 & n731 ) | ( ~n499 & n6220 ) | ( n731 & n6220 ) ;
  assign n6222 = ~n731 & n6221 ;
  assign n6223 = n103 | n862 ;
  assign n6224 = n6222 & ~n6223 ;
  assign n6225 = ~n5367 & n6224 ;
  assign n6226 = n520 | n5755 ;
  assign n6227 = ~n101 & n6029 ;
  assign n6228 = ( ~n302 & n731 ) | ( ~n302 & n5923 ) | ( n731 & n5923 ) ;
  assign n6229 = n302 | n6228 ;
  assign n6230 = ( ~n207 & n644 ) | ( ~n207 & n6229 ) | ( n644 & n6229 ) ;
  assign n6231 = ( ~n499 & n1485 ) | ( ~n499 & n4644 ) | ( n1485 & n4644 ) ;
  assign n6232 = ( n101 & ~n304 ) | ( n101 & n4149 ) | ( ~n304 & n4149 ) ;
  assign n6233 = ~n101 & n6232 ;
  assign n6234 = n103 | n6153 ;
  assign n6235 = n916 | n5170 ;
  assign n6236 = ( n304 & ~n872 ) | ( n304 & n6235 ) | ( ~n872 & n6235 ) ;
  assign n6237 = n872 | n6236 ;
  assign n6238 = ~n578 & n6047 ;
  assign n6239 = ( ~n96 & n1679 ) | ( ~n96 & n5878 ) | ( n1679 & n5878 ) ;
  assign n6240 = ~n1679 & n6239 ;
  assign n6241 = ( ~n605 & n943 ) | ( ~n605 & n6227 ) | ( n943 & n6227 ) ;
  assign n6242 = ( ~n1837 & n5945 ) | ( ~n1837 & n6218 ) | ( n5945 & n6218 ) ;
  assign n6243 = n1837 | n6242 ;
  assign n6244 = ( ~n1679 & n5358 ) | ( ~n1679 & n6218 ) | ( n5358 & n6218 ) ;
  assign n6245 = n1679 | n6244 ;
  assign n6246 = n86 | n6114 ;
  assign n6247 = ( n304 & ~n520 ) | ( n304 & n6246 ) | ( ~n520 & n6246 ) ;
  assign n6248 = n520 | n6247 ;
  assign n6249 = ~n101 & n6159 ;
  assign n6250 = ( ~n499 & n593 ) | ( ~n499 & n6199 ) | ( n593 & n6199 ) ;
  assign n6251 = ( ~n318 & n731 ) | ( ~n318 & n4523 ) | ( n731 & n4523 ) ;
  assign n6252 = ~n731 & n6251 ;
  assign n6253 = ( n349 & ~n375 ) | ( n349 & n6252 ) | ( ~n375 & n6252 ) ;
  assign n6254 = ~n349 & n6253 ;
  assign n6255 = ( ~n433 & n713 ) | ( ~n433 & n6254 ) | ( n713 & n6254 ) ;
  assign n6256 = n731 | n6016 ;
  assign n6257 = ( n164 & ~n887 ) | ( n164 & n6226 ) | ( ~n887 & n6226 ) ;
  assign n6258 = n887 | n6257 ;
  assign n6259 = ( n608 & ~n827 ) | ( n608 & n6258 ) | ( ~n827 & n6258 ) ;
  assign n6260 = n827 | n6259 ;
  assign n6261 = n651 | n6260 ;
  assign n6262 = n6173 & ~n6261 ;
  assign n6263 = ~n211 & n6262 ;
  assign n6264 = ( n502 & ~n829 ) | ( n502 & n6263 ) | ( ~n829 & n6263 ) ;
  assign n6265 = ~n502 & n6264 ;
  assign n6266 = ( ~n397 & n941 ) | ( ~n397 & n6265 ) | ( n941 & n6265 ) ;
  assign n6267 = ~n941 & n6266 ;
  assign n6268 = ( n349 & ~n591 ) | ( n349 & n6127 ) | ( ~n591 & n6127 ) ;
  assign n6269 = n207 | n6230 ;
  assign n6270 = ~n490 & n2419 ;
  assign n6271 = ( ~n433 & n502 ) | ( ~n433 & n6270 ) | ( n502 & n6270 ) ;
  assign n6272 = ~n502 & n6271 ;
  assign n6273 = n887 | n6136 ;
  assign n6274 = ( ~n397 & n643 ) | ( ~n397 & n5521 ) | ( n643 & n5521 ) ;
  assign n6275 = n397 | n6274 ;
  assign n6276 = n731 | n6140 ;
  assign n6277 = ( n302 & ~n318 ) | ( n302 & n5947 ) | ( ~n318 & n5947 ) ;
  assign n6278 = n302 | n6110 ;
  assign n6279 = ( ~n941 & n943 ) | ( ~n941 & n6278 ) | ( n943 & n6278 ) ;
  assign n6280 = n941 | n6279 ;
  assign n6281 = ( ~n601 & n4594 ) | ( ~n601 & n6280 ) | ( n4594 & n6280 ) ;
  assign n6282 = ( ~n207 & n362 ) | ( ~n207 & n2107 ) | ( n362 & n2107 ) ;
  assign n6283 = ( ~n5206 & n6055 ) | ( ~n5206 & n6261 ) | ( n6055 & n6261 ) ;
  assign n6284 = ~n6261 & n6283 ;
  assign n6285 = ( ~n302 & n916 ) | ( ~n302 & n6284 ) | ( n916 & n6284 ) ;
  assign n6286 = ~n916 & n6285 ;
  assign n6287 = ( n211 & ~n747 ) | ( n211 & n6161 ) | ( ~n747 & n6161 ) ;
  assign n6288 = ~n211 & n6287 ;
  assign n6289 = ( ~n147 & n5206 ) | ( ~n147 & n6065 ) | ( n5206 & n6065 ) ;
  assign n6290 = ~n5206 & n6289 ;
  assign n6291 = ~n713 & n6255 ;
  assign n6292 = ( n416 & ~n643 ) | ( n416 & n6209 ) | ( ~n643 & n6209 ) ;
  assign n6293 = ~n416 & n6292 ;
  assign n6294 = ( ~n209 & n717 ) | ( ~n209 & n6293 ) | ( n717 & n6293 ) ;
  assign n6295 = ~n532 & n5873 ;
  assign n6296 = ( n89 & ~n375 ) | ( n89 & n6295 ) | ( ~n375 & n6295 ) ;
  assign n6297 = ~n825 & n5797 ;
  assign n6298 = ~n417 & n6019 ;
  assign n6299 = ~n943 & n6241 ;
  assign n6300 = n591 | n6268 ;
  assign n6301 = ~n943 & n6128 ;
  assign n6302 = ( ~n100 & n147 ) | ( ~n100 & n6301 ) | ( n147 & n6301 ) ;
  assign n6303 = n96 | n6186 ;
  assign n6304 = ~n423 & n5935 ;
  assign n6305 = ( n248 & ~n900 ) | ( n248 & n6304 ) | ( ~n900 & n6304 ) ;
  assign n6306 = n295 | n3648 ;
  assign n6307 = ~n1485 & n6231 ;
  assign n6308 = ~n810 & n6233 ;
  assign n6309 = ( n250 & ~n352 ) | ( n250 & n2071 ) | ( ~n352 & n2071 ) ;
  assign n6310 = n352 | n6309 ;
  assign n6311 = ( ~n825 & n1485 ) | ( ~n825 & n5859 ) | ( n1485 & n5859 ) ;
  assign n6312 = n825 | n6311 ;
  assign n6313 = ( ~n100 & n660 ) | ( ~n100 & n6312 ) | ( n660 & n6312 ) ;
  assign n6314 = n100 | n6313 ;
  assign n6315 = ( ~n825 & n943 ) | ( ~n825 & n5888 ) | ( n943 & n5888 ) ;
  assign n6316 = ~n943 & n6315 ;
  assign n6317 = ~n290 & n6143 ;
  assign n6318 = n213 | n660 ;
  assign n6319 = n5014 | n6237 ;
  assign n6320 = n6318 | n6319 ;
  assign n6321 = ( n122 & ~n210 ) | ( n122 & n5761 ) | ( ~n210 & n5761 ) ;
  assign n6322 = ( n96 & ~n747 ) | ( n96 & n5092 ) | ( ~n747 & n5092 ) ;
  assign n6323 = ~n295 & n4709 ;
  assign n6324 = ( n173 & ~n352 ) | ( n173 & n6323 ) | ( ~n352 & n6323 ) ;
  assign n6325 = n86 | n5915 ;
  assign n6326 = ( n167 & ~n829 ) | ( n167 & n6325 ) | ( ~n829 & n6325 ) ;
  assign n6327 = n829 | n6326 ;
  assign n6328 = ( n371 & ~n489 ) | ( n371 & n6327 ) | ( ~n489 & n6327 ) ;
  assign n6329 = n489 | n6328 ;
  assign n6330 = ( n96 & ~n900 ) | ( n96 & n6109 ) | ( ~n900 & n6109 ) ;
  assign n6331 = n900 | n6330 ;
  assign n6332 = ( n583 & n702 ) | ( n583 & ~n6331 ) | ( n702 & ~n6331 ) ;
  assign n6333 = ( n167 & ~n723 ) | ( n167 & n6048 ) | ( ~n723 & n6048 ) ;
  assign n6334 = n723 | n6333 ;
  assign n6335 = ( ~n658 & n659 ) | ( ~n658 & n6334 ) | ( n659 & n6334 ) ;
  assign n6336 = n658 | n6335 ;
  assign n6337 = ( n122 & ~n827 ) | ( n122 & n6336 ) | ( ~n827 & n6336 ) ;
  assign n6338 = ( ~n279 & n375 ) | ( ~n279 & n5804 ) | ( n375 & n5804 ) ;
  assign n6339 = ~n250 & n4251 ;
  assign n6340 = ~n300 & n5956 ;
  assign n6341 = ( n417 & ~n423 ) | ( n417 & n6340 ) | ( ~n423 & n6340 ) ;
  assign n6342 = ~n417 & n6341 ;
  assign n6343 = ( ~n489 & n717 ) | ( ~n489 & n5861 ) | ( n717 & n5861 ) ;
  assign n6344 = ( n290 & ~n300 ) | ( n290 & n6243 ) | ( ~n300 & n6243 ) ;
  assign n6345 = n300 | n6344 ;
  assign n6346 = ( n583 & n960 ) | ( n583 & ~n6345 ) | ( n960 & ~n6345 ) ;
  assign n6347 = ( n348 & ~n591 ) | ( n348 & n5175 ) | ( ~n591 & n5175 ) ;
  assign n6348 = n591 | n6347 ;
  assign n6349 = ~n100 & n5703 ;
  assign n6350 = ( ~n300 & n1485 ) | ( ~n300 & n6150 ) | ( n1485 & n6150 ) ;
  assign n6351 = ~n1485 & n6350 ;
  assign n6352 = ( n250 & ~n442 ) | ( n250 & n6245 ) | ( ~n442 & n6245 ) ;
  assign n6353 = n442 | n6352 ;
  assign n6354 = ( n122 & n583 ) | ( n122 & ~n6353 ) | ( n583 & ~n6353 ) ;
  assign n6355 = ~n122 & n6354 ;
  assign n6356 = ( ~n555 & n559 ) | ( ~n555 & n6355 ) | ( n559 & n6355 ) ;
  assign n6357 = ( ~n219 & n295 ) | ( ~n219 & n5835 ) | ( n295 & n5835 ) ;
  assign n6358 = ( n229 & ~n295 ) | ( n229 & n5364 ) | ( ~n295 & n5364 ) ;
  assign n6359 = ( n589 & ~n810 ) | ( n589 & n5747 ) | ( ~n810 & n5747 ) ;
  assign n6360 = n810 | n6359 ;
  assign n6361 = ( ~n96 & n713 ) | ( ~n96 & n4721 ) | ( n713 & n4721 ) ;
  assign n6362 = ~n713 & n6361 ;
  assign n6363 = ( ~n161 & n290 ) | ( ~n161 & n5417 ) | ( n290 & n5417 ) ;
  assign n6364 = n721 | n6314 ;
  assign n6365 = n318 | n6277 ;
  assign n6366 = ~n229 & n5849 ;
  assign n6367 = ~n786 & n5396 ;
  assign n6368 = ( n169 & ~n643 ) | ( n169 & n5779 ) | ( ~n643 & n5779 ) ;
  assign n6369 = ( ~n318 & n643 ) | ( ~n318 & n6115 ) | ( n643 & n6115 ) ;
  assign n6370 = n447 | n6164 ;
  assign n6371 = n643 | n6012 ;
  assign n6372 = ~n546 & n5796 ;
  assign n6373 = ( ~n643 & n660 ) | ( ~n643 & n5626 ) | ( n660 & n5626 ) ;
  assign n6374 = ~n229 & n5959 ;
  assign n6375 = n643 | n6368 ;
  assign n6376 = ( n173 & ~n714 ) | ( n173 & n6365 ) | ( ~n714 & n6365 ) ;
  assign n6377 = n161 | n6363 ;
  assign n6378 = ( ~n442 & n546 ) | ( ~n442 & n6366 ) | ( n546 & n6366 ) ;
  assign n6379 = ~n546 & n6378 ;
  assign n6380 = ( ~n351 & n5033 ) | ( ~n351 & n6379 ) | ( n5033 & n6379 ) ;
  assign n6381 = ~n5033 & n6380 ;
  assign n6382 = ( n247 & ~n702 ) | ( n247 & n6377 ) | ( ~n702 & n6377 ) ;
  assign n6383 = ~n247 & n5420 ;
  assign n6384 = ( n448 & ~n834 ) | ( n448 & n6367 ) | ( ~n834 & n6367 ) ;
  assign n6385 = ~n448 & n6384 ;
  assign n6386 = ( n371 & ~n735 ) | ( n371 & n6385 ) | ( ~n735 & n6385 ) ;
  assign n6387 = ( n448 & ~n659 ) | ( n448 & n6339 ) | ( ~n659 & n6339 ) ;
  assign n6388 = ( ~n447 & n490 ) | ( ~n447 & n6015 ) | ( n490 & n6015 ) ;
  assign n6389 = ~n490 & n6388 ;
  assign n6390 = ( n124 & ~n735 ) | ( n124 & n6389 ) | ( ~n735 & n6389 ) ;
  assign n6391 = ( n447 & ~n714 ) | ( n447 & n5629 ) | ( ~n714 & n5629 ) ;
  assign n6392 = ~n447 & n6391 ;
  assign n6393 = ~n247 & n6392 ;
  assign n6394 = ( n161 & ~n447 ) | ( n161 & n6317 ) | ( ~n447 & n6317 ) ;
  assign n6395 = ~n229 & n6358 ;
  assign n6396 = ( ~n318 & n546 ) | ( ~n318 & n6146 ) | ( n546 & n6146 ) ;
  assign n6397 = ~n229 & n6154 ;
  assign n6398 = ~n248 & n6305 ;
  assign n6399 = ( ~n161 & n348 ) | ( ~n161 & n6351 ) | ( n348 & n6351 ) ;
  assign n6400 = ( n490 & ~n834 ) | ( n490 & n5617 ) | ( ~n834 & n5617 ) ;
  assign n6401 = n318 | n6396 ;
  assign n6402 = n318 | n6369 ;
  assign n6403 = ~n490 & n6400 ;
  assign n6404 = ~n371 & n6386 ;
  assign n6405 = ( n448 & ~n827 ) | ( n448 & n6370 ) | ( ~n827 & n6370 ) ;
  assign n6406 = ~n448 & n6387 ;
  assign n6407 = ~n124 & n6390 ;
  assign n6408 = ( ~n184 & n786 ) | ( ~n184 & n4244 ) | ( n786 & n4244 ) ;
  assign n6409 = ( n248 & ~n788 ) | ( n248 & n6375 ) | ( ~n788 & n6375 ) ;
  assign n6410 = ~n161 & n6394 ;
  assign n6411 = n714 | n6376 ;
  assign n6412 = ~n287 & n6165 ;
  assign n6413 = n228 | n6014 ;
  assign n6414 = ( ~n221 & n719 ) | ( ~n221 & n6413 ) | ( n719 & n6413 ) ;
  assign n6415 = n221 | n6414 ;
  assign n6416 = ( ~n232 & n501 ) | ( ~n232 & n6407 ) | ( n501 & n6407 ) ;
  assign n6417 = ( ~n182 & n786 ) | ( ~n182 & n5300 ) | ( n786 & n5300 ) ;
  assign n6418 = n786 | n4457 ;
  assign n6419 = ( ~n348 & n593 ) | ( ~n348 & n6177 ) | ( n593 & n6177 ) ;
  assign n6420 = ~n593 & n6419 ;
  assign n6421 = ( n172 & ~n287 ) | ( n172 & n6071 ) | ( ~n287 & n6071 ) ;
  assign n6422 = n287 | n6421 ;
  assign n6423 = ( ~n754 & n955 ) | ( ~n754 & n6297 ) | ( n955 & n6297 ) ;
  assign n6424 = ( n232 & ~n834 ) | ( n232 & n6300 ) | ( ~n834 & n6300 ) ;
  assign n6425 = n754 | n6036 ;
  assign n6426 = ~n86 & n3566 ;
  assign n6427 = ( n167 & ~n423 ) | ( n167 & n6426 ) | ( ~n423 & n6426 ) ;
  assign n6428 = ~n788 & n6272 ;
  assign n6429 = n788 | n6409 ;
  assign n6430 = ( ~n423 & n754 ) | ( ~n423 & n6316 ) | ( n754 & n6316 ) ;
  assign n6431 = ~n754 & n6430 ;
  assign n6432 = ~n287 & n6374 ;
  assign n6433 = ( ~n410 & n593 ) | ( ~n410 & n6046 ) | ( n593 & n6046 ) ;
  assign n6434 = ~n221 & n5270 ;
  assign n6435 = ( n169 & ~n723 ) | ( n169 & n6434 ) | ( ~n723 & n6434 ) ;
  assign n6436 = ( ~n86 & n960 ) | ( ~n86 & n5872 ) | ( n960 & n5872 ) ;
  assign n6437 = n86 | n6436 ;
  assign n6438 = ( ~n197 & n362 ) | ( ~n197 & n6437 ) | ( n362 & n6437 ) ;
  assign n6439 = n197 | n6438 ;
  assign n6440 = n739 | n6439 ;
  assign n6441 = ( ~n357 & n719 ) | ( ~n357 & n6240 ) | ( n719 & n6240 ) ;
  assign n6442 = ~n719 & n6441 ;
  assign n6443 = ~n107 & n6442 ;
  assign n6444 = ~n559 & n6356 ;
  assign n6445 = ( ~n107 & n645 ) | ( ~n107 & n6444 ) | ( n645 & n6444 ) ;
  assign n6446 = n86 | n6152 ;
  assign n6447 = n423 | n5326 ;
  assign n6448 = ( ~n184 & n719 ) | ( ~n184 & n6447 ) | ( n719 & n6447 ) ;
  assign n6449 = ~n593 & n6250 ;
  assign n6450 = ( ~n723 & n788 ) | ( ~n723 & n6449 ) | ( n788 & n6449 ) ;
  assign n6451 = ~n788 & n6450 ;
  assign n6452 = ( ~n476 & n559 ) | ( ~n476 & n6291 ) | ( n559 & n6291 ) ;
  assign n6453 = ~n559 & n6452 ;
  assign n6454 = ( n162 & ~n834 ) | ( n162 & n6402 ) | ( ~n834 & n6402 ) ;
  assign n6455 = n834 | n6454 ;
  assign n6456 = ~n960 & n6119 ;
  assign n6457 = ( ~n612 & n779 ) | ( ~n612 & n6456 ) | ( n779 & n6456 ) ;
  assign n6458 = ( ~n124 & n148 ) | ( ~n124 & n6267 ) | ( n148 & n6267 ) ;
  assign n6459 = ~n148 & n6458 ;
  assign n6460 = ~n89 & n6296 ;
  assign n6461 = ~n414 & n6460 ;
  assign n6462 = ~n442 & n6299 ;
  assign n6463 = n834 | n6424 ;
  assign n6464 = n468 | n6463 ;
  assign n6465 = ( n148 & ~n442 ) | ( n148 & n6190 ) | ( ~n442 & n6190 ) ;
  assign n6466 = n442 | n6465 ;
  assign n6467 = ( ~n182 & n645 ) | ( ~n182 & n6466 ) | ( n645 & n6466 ) ;
  assign n6468 = n182 | n6467 ;
  assign n6469 = n381 | n6468 ;
  assign n6470 = ( ~n442 & n955 ) | ( ~n442 & n6269 ) | ( n955 & n6269 ) ;
  assign n6471 = n442 | n6470 ;
  assign n6472 = ( ~n400 & n468 ) | ( ~n400 & n6471 ) | ( n468 & n6471 ) ;
  assign n6473 = ~n172 & n6183 ;
  assign n6474 = ( ~n102 & n660 ) | ( ~n102 & n6473 ) | ( n660 & n6473 ) ;
  assign n6475 = ~n660 & n6474 ;
  assign n6476 = ( ~n164 & n188 ) | ( ~n164 & n6475 ) | ( n188 & n6475 ) ;
  assign n6477 = ~n188 & n6476 ;
  assign n6478 = n145 | n5642 ;
  assign n6479 = ( n124 & ~n197 ) | ( n124 & n6478 ) | ( ~n197 & n6478 ) ;
  assign n6480 = n197 | n6479 ;
  assign n6481 = ~n167 & n6427 ;
  assign n6482 = ( ~n197 & n378 ) | ( ~n197 & n6481 ) | ( n378 & n6481 ) ;
  assign n6483 = ( n124 & ~n747 ) | ( n124 & n6306 ) | ( ~n747 & n6306 ) ;
  assign n6484 = ( n162 & ~n649 ) | ( n162 & n5597 ) | ( ~n649 & n5597 ) ;
  assign n6485 = n649 | n6484 ;
  assign n6486 = n173 | n6137 ;
  assign n6487 = n102 | n6039 ;
  assign n6488 = ~n124 & n6188 ;
  assign n6489 = ( n649 & ~n827 ) | ( n649 & n6307 ) | ( ~n827 & n6307 ) ;
  assign n6490 = ~n649 & n6489 ;
  assign n6491 = ( ~n169 & n172 ) | ( ~n169 & n6142 ) | ( n172 & n6142 ) ;
  assign n6492 = ~n172 & n6491 ;
  assign n6493 = n173 | n1708 ;
  assign n6494 = ~n173 & n6324 ;
  assign n6495 = ( ~n162 & n348 ) | ( ~n162 & n6494 ) | ( n348 & n6494 ) ;
  assign n6496 = ~n348 & n6495 ;
  assign n6497 = ~n173 & n5335 ;
  assign n6498 = ( ~n210 & n612 ) | ( ~n210 & n6196 ) | ( n612 & n6196 ) ;
  assign n6499 = ~n612 & n6498 ;
  assign n6500 = ~n169 & n6435 ;
  assign n6501 = n279 | n6338 ;
  assign n6502 = ( n559 & ~n694 ) | ( n559 & n6501 ) | ( ~n694 & n6501 ) ;
  assign n6503 = n162 | n6053 ;
  assign n6504 = ( n124 & ~n416 ) | ( n124 & n6503 ) | ( ~n416 & n6503 ) ;
  assign n6505 = n416 | n6504 ;
  assign n6506 = ( n111 & ~n162 ) | ( n111 & n6348 ) | ( ~n162 & n6348 ) ;
  assign n6507 = n162 | n6506 ;
  assign n6508 = ~n348 & n6399 ;
  assign n6509 = ( n111 & ~n530 ) | ( n111 & n6508 ) | ( ~n530 & n6508 ) ;
  assign n6510 = ~n111 & n6509 ;
  assign n6511 = ( ~n362 & n532 ) | ( ~n362 & n6286 ) | ( n532 & n6286 ) ;
  assign n6512 = ~n532 & n6511 ;
  assign n6513 = ~n416 & n5715 ;
  assign n6514 = ( n148 & ~n184 ) | ( n148 & n6493 ) | ( ~n184 & n6493 ) ;
  assign n6515 = ( ~n145 & n162 ) | ( ~n145 & n6395 ) | ( n162 & n6395 ) ;
  assign n6516 = ~n162 & n6515 ;
  assign n6517 = ( n172 & ~n414 ) | ( n172 & n6516 ) | ( ~n414 & n6516 ) ;
  assign n6518 = ~n172 & n6517 ;
  assign n6519 = ( ~n102 & n532 ) | ( ~n102 & n6249 ) | ( n532 & n6249 ) ;
  assign n6520 = ~n532 & n6519 ;
  assign n6521 = ( ~n147 & n169 ) | ( ~n147 & n6202 ) | ( n169 & n6202 ) ;
  assign n6522 = ~n169 & n6521 ;
  assign n6523 = ( n833 & ~n834 ) | ( n833 & n6522 ) | ( ~n834 & n6522 ) ;
  assign n6524 = n655 | n6009 ;
  assign n6525 = ( n89 & ~n362 ) | ( n89 & n6412 ) | ( ~n362 & n6412 ) ;
  assign n6526 = ~n89 & n6525 ;
  assign n6527 = ( ~n476 & n756 ) | ( ~n476 & n6415 ) | ( n756 & n6415 ) ;
  assign n6528 = n476 | n6527 ;
  assign n6529 = n177 | n6528 ;
  assign n6530 = n779 | n6171 ;
  assign n6531 = ( n552 & ~n715 ) | ( n552 & n6530 ) | ( ~n715 & n6530 ) ;
  assign n6532 = ~n501 & n6416 ;
  assign n6533 = ~n444 & n6532 ;
  assign n6534 = ~n779 & n6457 ;
  assign n6535 = ( ~n184 & n779 ) | ( ~n184 & n6208 ) | ( n779 & n6208 ) ;
  assign n6536 = ~n779 & n6535 ;
  assign n6537 = ~n717 & n6294 ;
  assign n6538 = ( ~n717 & n747 ) | ( ~n717 & n6420 ) | ( n747 & n6420 ) ;
  assign n6539 = ~n955 & n6423 ;
  assign n6540 = n89 | n6028 ;
  assign n6541 = ~n89 & n6180 ;
  assign n6542 = n476 | n6425 ;
  assign n6543 = n362 | n6542 ;
  assign n6544 = ( ~n164 & n362 ) | ( ~n164 & n6480 ) | ( n362 & n6480 ) ;
  assign n6545 = n164 | n6544 ;
  assign n6546 = n747 | n6483 ;
  assign n6547 = n476 | n6546 ;
  assign n6548 = ( ~n88 & n779 ) | ( ~n88 & n6485 ) | ( n779 & n6485 ) ;
  assign n6549 = n88 | n6548 ;
  assign n6550 = ( ~n372 & n945 ) | ( ~n372 & n6549 ) | ( n945 & n6549 ) ;
  assign n6551 = ( n164 & ~n600 ) | ( n164 & n6487 ) | ( ~n600 & n6487 ) ;
  assign n6552 = ( ~n343 & n827 ) | ( ~n343 & n6276 ) | ( n827 & n6276 ) ;
  assign n6553 = n343 | n6552 ;
  assign n6554 = n655 | n6553 ;
  assign n6555 = ( ~n145 & n953 ) | ( ~n145 & n6310 ) | ( n953 & n6310 ) ;
  assign n6556 = n145 | n6555 ;
  assign n6557 = ( n717 & ~n942 ) | ( n717 & n6556 ) | ( ~n942 & n6556 ) ;
  assign n6558 = n942 | n6557 ;
  assign n6559 = n184 | n6408 ;
  assign n6560 = ~n955 & n6102 ;
  assign n6561 = ~n177 & n6560 ;
  assign n6562 = n184 | n6514 ;
  assign n6563 = ( ~n589 & n955 ) | ( ~n589 & n6403 ) | ( n955 & n6403 ) ;
  assign n6564 = ( ~n351 & n701 ) | ( ~n351 & n6401 ) | ( n701 & n6401 ) ;
  assign n6565 = n351 | n6564 ;
  assign n6566 = ~n357 & n6499 ;
  assign n6567 = ( n600 & ~n942 ) | ( n600 & n6149 ) | ( ~n942 & n6149 ) ;
  assign n6568 = ~n717 & n6343 ;
  assign n6569 = ( n231 & ~n444 ) | ( n231 & n6568 ) | ( ~n444 & n6568 ) ;
  assign n6570 = n228 | n5989 ;
  assign n6571 = ~n362 & n5660 ;
  assign n6572 = ~n6570 & n6571 ;
  assign n6573 = ~n5976 & n6572 ;
  assign n6574 = n340 | n6542 ;
  assign n6575 = n6570 | n6574 ;
  assign n6576 = ~n960 & n6346 ;
  assign n6577 = ( n88 & ~n231 ) | ( n88 & n6576 ) | ( ~n231 & n6576 ) ;
  assign n6578 = ~n88 & n6577 ;
  assign n6579 = ~n955 & n6563 ;
  assign n6580 = ~n945 & n6349 ;
  assign n6581 = ~n362 & n6282 ;
  assign n6582 = ( n351 & ~n357 ) | ( n351 & n6581 ) | ( ~n357 & n6581 ) ;
  assign n6583 = ~n351 & n6582 ;
  assign n6584 = ( ~n164 & n973 ) | ( ~n164 & n5294 ) | ( n973 & n5294 ) ;
  assign n6585 = n164 | n6584 ;
  assign n6586 = n967 | n6585 ;
  assign n6587 = ( ~n343 & n942 ) | ( ~n343 & n6446 ) | ( n942 & n6446 ) ;
  assign n6588 = n343 | n6587 ;
  assign n6589 = n145 | n6060 ;
  assign n6590 = ( n357 & ~n651 ) | ( n357 & n6589 ) | ( ~n651 & n6589 ) ;
  assign n6591 = n184 | n6448 ;
  assign n6592 = ( n146 & ~n967 ) | ( n146 & n6397 ) | ( ~n967 & n6397 ) ;
  assign n6593 = ( ~n145 & n552 ) | ( ~n145 & n6158 ) | ( n552 & n6158 ) ;
  assign n6594 = ~n552 & n6593 ;
  assign n6595 = ( n87 & ~n343 ) | ( n87 & n5773 ) | ( ~n343 & n5773 ) ;
  assign n6596 = n827 | n6405 ;
  assign n6597 = n862 | n5975 ;
  assign n6598 = n715 | n6531 ;
  assign n6599 = ( ~n87 & n530 ) | ( ~n87 & n6598 ) | ( n530 & n6598 ) ;
  assign n6600 = n87 | n6599 ;
  assign n6601 = ( ~n279 & n701 ) | ( ~n279 & n6455 ) | ( n701 & n6455 ) ;
  assign n6602 = ~n187 & n5451 ;
  assign n6603 = n182 | n6417 ;
  assign n6604 = ( n501 & ~n862 ) | ( n501 & n6418 ) | ( ~n862 & n6418 ) ;
  assign n6605 = n862 | n6604 ;
  assign n6606 = ( n146 & ~n973 ) | ( n146 & n6225 ) | ( ~n973 & n6225 ) ;
  assign n6607 = ~n701 & n5937 ;
  assign n6608 = ( ~n651 & n969 ) | ( ~n651 & n6607 ) | ( n969 & n6607 ) ;
  assign n6609 = ~n147 & n6302 ;
  assign n6610 = ( n378 & ~n589 ) | ( n378 & n6609 ) | ( ~n589 & n6609 ) ;
  assign n6611 = ( n833 & ~n849 ) | ( n833 & n4259 ) | ( ~n849 & n4259 ) ;
  assign n6612 = ~n833 & n6611 ;
  assign n6613 = n167 | n5948 ;
  assign n6614 = ( n589 & ~n694 ) | ( n589 & n6078 ) | ( ~n694 & n6078 ) ;
  assign n6615 = ~n589 & n6614 ;
  assign n6616 = ( n219 & ~n833 ) | ( n219 & n6615 ) | ( ~n833 & n6615 ) ;
  assign n6617 = ~n651 & n6537 ;
  assign n6618 = ( ~n659 & n973 ) | ( ~n659 & n6383 ) | ( n973 & n6383 ) ;
  assign n6619 = ~n973 & n6618 ;
  assign n6620 = ( ~n147 & n960 ) | ( ~n147 & n6185 ) | ( n960 & n6185 ) ;
  assign n6621 = n147 | n6620 ;
  assign n6622 = ( ~n167 & n530 ) | ( ~n167 & n6621 ) | ( n530 & n6621 ) ;
  assign n6623 = n167 | n6622 ;
  assign n6624 = ( ~n147 & n653 ) | ( ~n147 & n6273 ) | ( n653 & n6273 ) ;
  assign n6625 = n147 | n6624 ;
  assign n6626 = ( ~n501 & n715 ) | ( ~n501 & n6625 ) | ( n715 & n6625 ) ;
  assign n6627 = n501 | n6626 ;
  assign n6628 = ( ~n694 & n973 ) | ( ~n694 & n6429 ) | ( n973 & n6429 ) ;
  assign n6629 = ~n701 & n4706 ;
  assign n6630 = n589 | n6562 ;
  assign n6631 = ( ~n167 & n715 ) | ( ~n167 & n6410 ) | ( n715 & n6410 ) ;
  assign n6632 = ~n715 & n6631 ;
  assign n6633 = ~n182 & n6496 ;
  assign n6634 = ~n702 & n6332 ;
  assign n6635 = ( n701 & ~n862 ) | ( n701 & n6634 ) | ( ~n862 & n6634 ) ;
  assign n6636 = ~n701 & n6635 ;
  assign n6637 = ( ~n182 & n219 ) | ( ~n182 & n6636 ) | ( n219 & n6636 ) ;
  assign n6638 = n827 | n6337 ;
  assign n6639 = ( n219 & ~n702 ) | ( n219 & n6500 ) | ( ~n702 & n6500 ) ;
  assign n6640 = ~n219 & n6639 ;
  assign n6641 = ~n849 & n6640 ;
  assign n6642 = ( ~n87 & n187 ) | ( ~n87 & n6583 ) | ( n187 & n6583 ) ;
  assign n6643 = ~n187 & n6642 ;
  assign n6644 = ( ~n827 & n961 ) | ( ~n827 & n6643 ) | ( n961 & n6643 ) ;
  assign n6645 = ( n715 & ~n862 ) | ( n715 & n6512 ) | ( ~n862 & n6512 ) ;
  assign n6646 = ~n715 & n6645 ;
  assign n6647 = ~n756 & n6646 ;
  assign n6648 = n651 | n6590 ;
  assign n6649 = n756 | n6591 ;
  assign n6650 = ~n87 & n6595 ;
  assign n6651 = n702 | n6382 ;
  assign n6652 = ~n833 & n6523 ;
  assign n6653 = ( n187 & ~n702 ) | ( n187 & n6162 ) | ( ~n702 & n6162 ) ;
  assign n6654 = n702 | n6653 ;
  assign n6655 = ( n628 & ~n963 ) | ( n628 & n6406 ) | ( ~n963 & n6406 ) ;
  assign n6656 = ( ~n425 & n653 ) | ( ~n425 & n5769 ) | ( n653 & n5769 ) ;
  assign n6657 = n279 | n6601 ;
  assign n6658 = ( ~n628 & n969 ) | ( ~n628 & n6536 ) | ( n969 & n6536 ) ;
  assign n6659 = n425 | n6656 ;
  assign n6660 = n694 | n6502 ;
  assign n6661 = ( ~n659 & n660 ) | ( ~n659 & n6288 ) | ( n660 & n6288 ) ;
  assign n6662 = n5913 | n5940 ;
  assign n6663 = n228 | n6662 ;
  assign n6664 = ~n969 & n6608 ;
  assign n6665 = ( n378 & ~n400 ) | ( n378 & n6594 ) | ( ~n400 & n6594 ) ;
  assign n6666 = ( ~n378 & n747 ) | ( ~n378 & n6398 ) | ( n747 & n6398 ) ;
  assign n6667 = ~n747 & n6666 ;
  assign n6668 = ~n747 & n6538 ;
  assign n6669 = n747 | n6322 ;
  assign n6670 = ~n378 & n6665 ;
  assign n6671 = ~n378 & n6482 ;
  assign n6672 = ~n378 & n6610 ;
  assign n6673 = n378 | n6023 ;
  assign n6674 = ( ~n279 & n653 ) | ( ~n279 & n6492 ) | ( n653 & n6492 ) ;
  assign n6675 = ~n210 & n6404 ;
  assign n6676 = ( ~n372 & n645 ) | ( ~n372 & n6329 ) | ( n645 & n6329 ) ;
  assign n6677 = ~n210 & n6632 ;
  assign n6678 = n210 | n6321 ;
  assign n6679 = ( ~n659 & n969 ) | ( ~n659 & n6303 ) | ( n969 & n6303 ) ;
  assign n6680 = ( ~n600 & n744 ) | ( ~n600 & n6194 ) | ( n744 & n6194 ) ;
  assign n6681 = n600 | n6551 ;
  assign n6682 = ~n653 & n6674 ;
  assign n6683 = ~n146 & n6592 ;
  assign n6684 = ~n146 & n6497 ;
  assign n6685 = ~n146 & n6606 ;
  assign n6686 = ~n600 & n6567 ;
  assign n6687 = n5982 | n6543 ;
  assign n6688 = n659 | n5325 ;
  assign n6689 = ( n425 & ~n600 ) | ( n425 & n6381 ) | ( ~n600 & n6381 ) ;
  assign n6690 = ~n960 & n6372 ;
  assign n6691 = n659 | n6275 ;
  assign n6692 = ~n960 & n6035 ;
  assign n6693 = n694 | n6628 ;
  assign n6694 = ( ~n400 & n963 ) | ( ~n400 & n6298 ) | ( n963 & n6298 ) ;
  assign n6695 = n279 | n5917 ;
  assign n6696 = n400 | n6472 ;
  assign n6697 = ~n660 & n6373 ;
  assign n6698 = n628 | n6248 ;
  assign n6699 = ~n961 & n6644 ;
  assign n6700 = n660 | n6411 ;
  assign n6701 = n580 | n5534 ;
  assign n6702 = n961 | n6651 ;
  assign n6703 = n600 | n6680 ;
  assign n6704 = ( ~n600 & n659 ) | ( ~n600 & n5778 ) | ( n659 & n5778 ) ;
  assign n6705 = ~n410 & n6362 ;
  assign n6706 = n372 | n6550 ;
  assign n6707 = ~n6663 & n6692 ;
  assign n6708 = ~n400 & n6612 ;
  assign n6709 = ~n279 & n5978 ;
  assign n6710 = n372 | n6676 ;
  assign n6711 = ~n659 & n6704 ;
  assign n6712 = ~n961 & n6667 ;
  assign n6713 = ~n628 & n6655 ;
  assign n6714 = n410 | n6433 ;
  assign n6715 = ~n660 & n6661 ;
  assign n6716 = n580 | n6681 ;
  assign n6717 = n410 | n6659 ;
  assign n6718 = ~n969 & n6658 ;
  assign n6719 = ( n653 & ~n744 ) | ( n653 & n6145 ) | ( ~n744 & n6145 ) ;
  assign n6720 = ( ~n372 & n530 ) | ( ~n372 & n6619 ) | ( n530 & n6619 ) ;
  assign n6721 = n659 | n6679 ;
  assign n6722 = n628 | n6507 ;
  assign n6723 = n694 | n6135 ;
  assign n6724 = n580 | n6657 ;
  assign n6725 = ~n653 & n6719 ;
  assign n6726 = n6543 | n6662 ;
  assign n6727 = ( ~n203 & n245 ) | ( ~n203 & n6453 ) | ( n245 & n6453 ) ;
  assign n6728 = ~n245 & n6727 ;
  assign n6729 = ~n219 & n6526 ;
  assign n6730 = ( ~n427 & n601 ) | ( ~n427 & n6534 ) | ( n601 & n6534 ) ;
  assign n6731 = ~n601 & n6730 ;
  assign n6732 = ( n271 & ~n645 ) | ( n271 & n6605 ) | ( ~n645 & n6605 ) ;
  assign n6733 = n645 | n6732 ;
  assign n6734 = ( n219 & ~n427 ) | ( n219 & n6459 ) | ( ~n427 & n6459 ) ;
  assign n6735 = ~n219 & n6734 ;
  assign n6736 = ( ~n425 & n426 ) | ( ~n425 & n6422 ) | ( n426 & n6422 ) ;
  assign n6737 = n425 | n6736 ;
  assign n6738 = ( n245 & ~n953 ) | ( n245 & n6737 ) | ( ~n953 & n6737 ) ;
  assign n6739 = n953 | n6738 ;
  assign n6740 = n271 | n6739 ;
  assign n6741 = ~n963 & n6694 ;
  assign n6742 = ( n203 & ~n425 ) | ( n203 & n6688 ) | ( ~n425 & n6688 ) ;
  assign n6743 = n425 | n6742 ;
  assign n6744 = n645 | n6743 ;
  assign n6745 = n271 | n6696 ;
  assign n6746 = ~n953 & n6541 ;
  assign n6747 = n953 | n6613 ;
  assign n6748 = ( n203 & ~n963 ) | ( n203 & n6723 ) | ( ~n963 & n6723 ) ;
  assign n6749 = n963 | n6748 ;
  assign n6750 = ( n426 & ~n427 ) | ( n426 & n6181 ) | ( ~n427 & n6181 ) ;
  assign n6751 = n427 | n6750 ;
  assign n6752 = ~n219 & n6616 ;
  assign n6753 = ~n530 & n6720 ;
  assign n6754 = n530 | n6706 ;
  assign n6755 = ( n426 & ~n434 ) | ( n426 & n6486 ) | ( ~n434 & n6486 ) ;
  assign n6756 = n434 | n6755 ;
  assign n6757 = ( n245 & ~n963 ) | ( n245 & n6756 ) | ( ~n963 & n6756 ) ;
  assign n6758 = n963 | n6757 ;
  assign n6759 = ~n203 & n6488 ;
  assign n6760 = ( ~n231 & n645 ) | ( ~n231 & n6693 ) | ( n645 & n6693 ) ;
  assign n6761 = n530 | n6558 ;
  assign n6762 = ( ~n426 & n601 ) | ( ~n426 & n6559 ) | ( n601 & n6559 ) ;
  assign n6763 = n426 | n6762 ;
  assign n6764 = ( ~n434 & n608 ) | ( ~n434 & n6431 ) | ( n608 & n6431 ) ;
  assign n6765 = ~n608 & n6764 ;
  assign n6766 = ( ~n427 & n608 ) | ( ~n427 & n6695 ) | ( n608 & n6695 ) ;
  assign n6767 = n427 | n6766 ;
  assign n6768 = n953 | n6565 ;
  assign n6769 = ( n426 & ~n744 ) | ( n426 & n6234 ) | ( ~n744 & n6234 ) ;
  assign n6770 = n744 | n6769 ;
  assign n6771 = ( ~n744 & n963 ) | ( ~n744 & n6669 ) | ( n963 & n6669 ) ;
  assign n6772 = n744 | n6771 ;
  assign n6773 = n530 | n6772 ;
  assign n6774 = ~n219 & n6637 ;
  assign n6775 = ~n608 & n6774 ;
  assign n6776 = ( n434 & ~n953 ) | ( n434 & n6238 ) | ( ~n953 & n6238 ) ;
  assign n6777 = ~n434 & n6776 ;
  assign n6778 = n601 | n6051 ;
  assign n6779 = ~n425 & n6689 ;
  assign n6780 = n601 | n6281 ;
  assign n6781 = ~n645 & n6445 ;
  assign n6782 = n219 | n6357 ;
  assign n6783 = ~n601 & n6518 ;
  assign n6784 = ( n203 & ~n608 ) | ( n203 & n6360 ) | ( ~n608 & n6360 ) ;
  assign n6785 = n608 | n6784 ;
  assign n6786 = ( ~n231 & n608 ) | ( ~n231 & n6198 ) | ( n608 & n6198 ) ;
  assign n6787 = x30 ^ x29 ^ 1'b0 ;
  assign n6788 = ~x31 & n6787 ;
  assign n6789 = x31 & n6787 ;
  assign n6790 = x31 & n36 ;
  assign n6791 = n6789 ^ n36 ^ x31 ;
  assign n6792 = n6740 & n6791 ;
  assign n6793 = ( ~n6461 & n6790 ) | ( ~n6461 & n6792 ) | ( n6790 & n6792 ) ;
  assign n6794 = ( ~n6668 & n6788 ) | ( ~n6668 & n6792 ) | ( n6788 & n6792 ) ;
  assign n6795 = n6792 | n6794 ;
  assign n6796 = n6793 | n6795 ;
  assign n6797 = ~n6461 & n6539 ;
  assign n6798 = n6797 ^ n6740 ^ 1'b0 ;
  assign n6799 = n6789 & n6798 ;
  assign n6800 = ( ~n6539 & n6790 ) | ( ~n6539 & n6799 ) | ( n6790 & n6799 ) ;
  assign n6801 = n6740 & ~n6788 ;
  assign n6802 = ( n6461 & n6539 ) | ( n6461 & ~n6740 ) | ( n6539 & ~n6740 ) ;
  assign n6803 = n6461 | n6802 ;
  assign n6804 = ( ~n6461 & n6791 ) | ( ~n6461 & n6799 ) | ( n6791 & n6799 ) ;
  assign n6805 = n6799 | n6804 ;
  assign n6806 = ( n6668 & ~n6740 ) | ( n6668 & n6803 ) | ( ~n6740 & n6803 ) ;
  assign n6807 = n6800 | n6805 ;
  assign n6808 = n6803 ^ n6740 ^ n6668 ;
  assign n6809 = ( n6740 & ~n6801 ) | ( n6740 & n6807 ) | ( ~n6801 & n6807 ) ;
  assign n6810 = n6789 & ~n6808 ;
  assign n6811 = n6806 ^ n6735 ^ n6668 ;
  assign n6812 = ( n6789 & n6796 ) | ( n6789 & ~n6810 ) | ( n6796 & ~n6810 ) ;
  assign n6813 = ~n6462 & n6809 ;
  assign n6814 = ( n6668 & n6735 ) | ( n6668 & n6806 ) | ( n6735 & n6806 ) ;
  assign n6815 = n6809 ^ n6462 ^ 1'b0 ;
  assign n6816 = n6813 ^ n6812 ^ n6664 ;
  assign n6817 = ( ~n6664 & n6812 ) | ( ~n6664 & n6813 ) | ( n6812 & n6813 ) ;
  assign n6818 = n6789 & ~n6811 ;
  assign n6819 = n231 | n6760 ;
  assign n6820 = ( ~n6668 & n6791 ) | ( ~n6668 & n6818 ) | ( n6791 & n6818 ) ;
  assign n6821 = n6818 | n6820 ;
  assign n6822 = ( n6740 & n6790 ) | ( n6740 & n6818 ) | ( n6790 & n6818 ) ;
  assign n6823 = n231 | n6749 ;
  assign n6824 = n231 | n6678 ;
  assign n6825 = n231 | n6786 ;
  assign n6826 = n6821 | n6822 ;
  assign n6827 = ~n231 & n6569 ;
  assign n6828 = n6814 ^ n6735 ^ n6685 ;
  assign n6829 = n6735 & n6788 ;
  assign n6830 = ( n6685 & n6735 ) | ( n6685 & n6814 ) | ( n6735 & n6814 ) ;
  assign n6831 = ( n6788 & n6826 ) | ( n6788 & ~n6829 ) | ( n6826 & ~n6829 ) ;
  assign n6832 = n6831 ^ n6817 ^ n6464 ;
  assign n6833 = ( n6464 & n6817 ) | ( n6464 & n6831 ) | ( n6817 & n6831 ) ;
  assign n6834 = n6789 & ~n6828 ;
  assign n6835 = ( ~n6735 & n6791 ) | ( ~n6735 & n6834 ) | ( n6791 & n6834 ) ;
  assign n6836 = n6834 | n6835 ;
  assign n6837 = ( ~n6668 & n6790 ) | ( ~n6668 & n6834 ) | ( n6790 & n6834 ) ;
  assign n6838 = n6836 | n6837 ;
  assign n6839 = n6685 & n6788 ;
  assign n6840 = ( n6788 & n6838 ) | ( n6788 & ~n6839 ) | ( n6838 & ~n6839 ) ;
  assign n6841 = n6840 ^ n6833 ^ n6672 ;
  assign n6842 = ( ~n6672 & n6833 ) | ( ~n6672 & n6840 ) | ( n6833 & n6840 ) ;
  assign n6843 = n6830 ^ n6733 ^ n6685 ;
  assign n6844 = n6789 & n6843 ;
  assign n6845 = ( ~n6685 & n6791 ) | ( ~n6685 & n6844 ) | ( n6791 & n6844 ) ;
  assign n6846 = n6844 | n6845 ;
  assign n6847 = ( ~n6735 & n6790 ) | ( ~n6735 & n6844 ) | ( n6790 & n6844 ) ;
  assign n6848 = n6846 | n6847 ;
  assign n6849 = n5851 & n6791 ;
  assign n6850 = ( n6685 & ~n6733 ) | ( n6685 & n6830 ) | ( ~n6733 & n6830 ) ;
  assign n6851 = ( n5851 & n6733 ) | ( n5851 & ~n6850 ) | ( n6733 & ~n6850 ) ;
  assign n6852 = n6733 & ~n6788 ;
  assign n6853 = ( n6256 & n6788 ) | ( n6256 & n6849 ) | ( n6788 & n6849 ) ;
  assign n6854 = ( n6733 & n6848 ) | ( n6733 & ~n6852 ) | ( n6848 & ~n6852 ) ;
  assign n6855 = n6849 | n6853 ;
  assign n6856 = ( n6540 & n6842 ) | ( n6540 & n6854 ) | ( n6842 & n6854 ) ;
  assign n6857 = n6854 ^ n6842 ^ n6540 ;
  assign n6858 = n6851 ^ n6256 ^ n5851 ;
  assign n6859 = n6789 & ~n6858 ;
  assign n6860 = n5851 & ~n6788 ;
  assign n6861 = n6850 ^ n6733 ^ n5851 ;
  assign n6862 = n6789 & ~n6861 ;
  assign n6863 = ( ~n6685 & n6790 ) | ( ~n6685 & n6862 ) | ( n6790 & n6862 ) ;
  assign n6864 = ( n6733 & n6790 ) | ( n6733 & n6849 ) | ( n6790 & n6849 ) ;
  assign n6865 = n6855 | n6864 ;
  assign n6866 = ( n6733 & n6791 ) | ( n6733 & n6862 ) | ( n6791 & n6862 ) ;
  assign n6867 = n6862 | n6866 ;
  assign n6868 = n6863 | n6867 ;
  assign n6869 = ( n5851 & ~n6860 ) | ( n5851 & n6868 ) | ( ~n6860 & n6868 ) ;
  assign n6870 = n6869 ^ n6856 ^ n6673 ;
  assign n6871 = ( n6789 & ~n6859 ) | ( n6789 & n6865 ) | ( ~n6859 & n6865 ) ;
  assign n6872 = ( x2 & n6744 ) | ( x2 & n6871 ) | ( n6744 & n6871 ) ;
  assign n6873 = ( n5851 & n6256 ) | ( n5851 & n6851 ) | ( n6256 & n6851 ) ;
  assign n6874 = ( n6256 & ~n6617 ) | ( n6256 & n6873 ) | ( ~n6617 & n6873 ) ;
  assign n6875 = ( x2 & n6469 ) | ( x2 & n6872 ) | ( n6469 & n6872 ) ;
  assign n6876 = ( n6673 & n6856 ) | ( n6673 & n6869 ) | ( n6856 & n6869 ) ;
  assign n6877 = n6874 ^ n6718 ^ n6617 ;
  assign n6878 = n6789 & n6877 ;
  assign n6879 = n6872 ^ n6469 ^ x2 ;
  assign n6880 = ( ~n6617 & n6791 ) | ( ~n6617 & n6878 ) | ( n6791 & n6878 ) ;
  assign n6881 = n6878 | n6880 ;
  assign n6882 = ( n6256 & n6790 ) | ( n6256 & n6878 ) | ( n6790 & n6878 ) ;
  assign n6883 = n6881 | n6882 ;
  assign n6884 = ( x2 & ~n6708 ) | ( x2 & n6875 ) | ( ~n6708 & n6875 ) ;
  assign n6885 = n6873 ^ n6617 ^ n6256 ;
  assign n6886 = n6871 ^ n6744 ^ x2 ;
  assign n6887 = n6789 & ~n6885 ;
  assign n6888 = ( n6617 & n6718 ) | ( n6617 & ~n6874 ) | ( n6718 & ~n6874 ) ;
  assign n6889 = n6875 ^ n6708 ^ x2 ;
  assign n6890 = ( n6256 & n6791 ) | ( n6256 & n6887 ) | ( n6791 & n6887 ) ;
  assign n6891 = n6887 | n6890 ;
  assign n6892 = ( n5851 & n6790 ) | ( n5851 & n6887 ) | ( n6790 & n6887 ) ;
  assign n6893 = n6891 | n6892 ;
  assign n6894 = n6718 & n6788 ;
  assign n6895 = ( n6788 & n6883 ) | ( n6788 & ~n6894 ) | ( n6883 & ~n6894 ) ;
  assign n6896 = n6617 & n6788 ;
  assign n6897 = ( n6788 & n6893 ) | ( n6788 & ~n6896 ) | ( n6893 & ~n6896 ) ;
  assign n6898 = x27 ^ x26 ^ 1'b0 ;
  assign n6899 = x28 ^ x27 ^ 1'b0 ;
  assign n6900 = x29 ^ x28 ^ 1'b0 ;
  assign n6901 = ~n6898 & n6899 ;
  assign n6902 = n6898 | n6900 ;
  assign n6903 = n6899 | n6902 ;
  assign n6904 = ~n6718 & n6901 ;
  assign n6905 = ( n6718 & n6731 ) | ( n6718 & n6888 ) | ( n6731 & n6888 ) ;
  assign n6906 = n6903 ^ n6901 ^ n6898 ;
  assign n6907 = n6898 & ~n6900 ;
  assign n6908 = ( ~n6617 & n6904 ) | ( ~n6617 & n6906 ) | ( n6904 & n6906 ) ;
  assign n6909 = n6904 | n6908 ;
  assign n6910 = ( ~n6731 & n6904 ) | ( ~n6731 & n6907 ) | ( n6904 & n6907 ) ;
  assign n6911 = n6256 & n6907 ;
  assign n6912 = n6909 | n6910 ;
  assign n6913 = ( n6733 & n6906 ) | ( n6733 & n6911 ) | ( n6906 & n6911 ) ;
  assign n6914 = ( n5851 & n6901 ) | ( n5851 & n6911 ) | ( n6901 & n6911 ) ;
  assign n6915 = n6911 | n6914 ;
  assign n6916 = n6913 | n6915 ;
  assign n6917 = n6888 ^ n6731 ^ n6718 ;
  assign n6918 = n6898 & n6900 ;
  assign n6919 = ~n6917 & n6918 ;
  assign n6920 = n6912 & ~n6919 ;
  assign n6921 = n6920 ^ n6919 ^ x29 ;
  assign n6922 = ( n6876 & n6886 ) | ( n6876 & n6921 ) | ( n6886 & n6921 ) ;
  assign n6923 = ( n6879 & n6897 ) | ( n6879 & n6922 ) | ( n6897 & n6922 ) ;
  assign n6924 = n6922 ^ n6897 ^ n6879 ;
  assign n6925 = n6923 ^ n6895 ^ n6889 ;
  assign n6926 = ( ~n6889 & n6895 ) | ( ~n6889 & n6923 ) | ( n6895 & n6923 ) ;
  assign n6927 = n6733 & n6907 ;
  assign n6928 = n6843 & n6918 ;
  assign n6929 = n6921 ^ n6886 ^ n6876 ;
  assign n6930 = ( ~n6685 & n6901 ) | ( ~n6685 & n6927 ) | ( n6901 & n6927 ) ;
  assign n6931 = n6927 | n6930 ;
  assign n6932 = ~n6461 & n6901 ;
  assign n6933 = ( ~n6735 & n6906 ) | ( ~n6735 & n6927 ) | ( n6906 & n6927 ) ;
  assign n6934 = n6808 & n6918 ;
  assign n6935 = n6931 | n6933 ;
  assign n6936 = n6928 | n6935 ;
  assign n6937 = n6740 & n6901 ;
  assign n6938 = ( ~n6539 & n6906 ) | ( ~n6539 & n6932 ) | ( n6906 & n6932 ) ;
  assign n6939 = n6932 | n6938 ;
  assign n6940 = ( n6740 & n6907 ) | ( n6740 & n6939 ) | ( n6907 & n6939 ) ;
  assign n6941 = n6939 | n6940 ;
  assign n6942 = ( n6798 & n6918 ) | ( n6798 & n6939 ) | ( n6918 & n6939 ) ;
  assign n6943 = n6936 ^ x29 ^ 1'b0 ;
  assign n6944 = n6941 | n6942 ;
  assign n6945 = ( ~n6461 & n6906 ) | ( ~n6461 & n6937 ) | ( n6906 & n6937 ) ;
  assign n6946 = n6937 | n6945 ;
  assign n6947 = ( ~n6668 & n6907 ) | ( ~n6668 & n6937 ) | ( n6907 & n6937 ) ;
  assign n6948 = n6946 | n6947 ;
  assign n6949 = n6934 | n6948 ;
  assign n6950 = ~n6735 & n6901 ;
  assign n6951 = n6858 & n6918 ;
  assign n6952 = n6916 | n6951 ;
  assign n6953 = n6949 ^ x29 ^ 1'b0 ;
  assign n6954 = n6944 ^ x29 ^ 1'b0 ;
  assign n6955 = ( ~n6668 & n6906 ) | ( ~n6668 & n6950 ) | ( n6906 & n6950 ) ;
  assign n6956 = n6950 | n6955 ;
  assign n6957 = ( ~n6685 & n6907 ) | ( ~n6685 & n6950 ) | ( n6907 & n6950 ) ;
  assign n6958 = n6956 | n6957 ;
  assign n6959 = ~n6828 & n6918 ;
  assign n6960 = n6958 | n6959 ;
  assign n6961 = n6960 ^ x29 ^ 1'b0 ;
  assign n6962 = n6539 ^ n6461 ^ 1'b0 ;
  assign n6963 = n6918 & n6962 ;
  assign n6964 = ( ~n6461 & n6907 ) | ( ~n6461 & n6963 ) | ( n6907 & n6963 ) ;
  assign n6965 = ( ~n6539 & n6901 ) | ( ~n6539 & n6963 ) | ( n6901 & n6963 ) ;
  assign n6966 = ~n6539 & n6898 ;
  assign n6967 = x29 & ~n6966 ;
  assign n6968 = n6963 | n6965 ;
  assign n6969 = n6964 | n6968 ;
  assign n6970 = n6969 ^ x29 ^ 1'b0 ;
  assign n6971 = n6967 & n6970 ;
  assign n6972 = n6954 & n6971 ;
  assign n6973 = n6970 ^ n6967 ^ 1'b0 ;
  assign n6974 = ~n6539 & n6787 ;
  assign n6975 = n6974 ^ n6972 ^ n6953 ;
  assign n6976 = ( n6953 & n6972 ) | ( n6953 & n6974 ) | ( n6972 & n6974 ) ;
  assign n6977 = n6789 & n6962 ;
  assign n6978 = ( ~n6539 & n6791 ) | ( ~n6539 & n6977 ) | ( n6791 & n6977 ) ;
  assign n6979 = n6977 | n6978 ;
  assign n6980 = ( ~n6461 & n6788 ) | ( ~n6461 & n6977 ) | ( n6788 & n6977 ) ;
  assign n6981 = n6979 | n6980 ;
  assign n6982 = n6740 & n6906 ;
  assign n6983 = n6971 ^ n6954 ^ 1'b0 ;
  assign n6984 = ( ~n6668 & n6901 ) | ( ~n6668 & n6982 ) | ( n6901 & n6982 ) ;
  assign n6985 = n6982 | n6984 ;
  assign n6986 = ( ~n6735 & n6907 ) | ( ~n6735 & n6982 ) | ( n6907 & n6982 ) ;
  assign n6987 = n6985 | n6986 ;
  assign n6988 = ~n6811 & n6918 ;
  assign n6989 = n6987 | n6988 ;
  assign n6990 = n6989 ^ x29 ^ 1'b0 ;
  assign n6991 = ( n6976 & n6981 ) | ( n6976 & n6990 ) | ( n6981 & n6990 ) ;
  assign n6992 = n6990 ^ n6981 ^ n6976 ;
  assign n6993 = ( ~n6815 & n6961 ) | ( ~n6815 & n6991 ) | ( n6961 & n6991 ) ;
  assign n6994 = ( ~n6816 & n6943 ) | ( ~n6816 & n6993 ) | ( n6943 & n6993 ) ;
  assign n6995 = n6993 ^ n6943 ^ n6816 ;
  assign n6996 = n6256 & n6906 ;
  assign n6997 = ( ~n6617 & n6901 ) | ( ~n6617 & n6996 ) | ( n6901 & n6996 ) ;
  assign n6998 = n6996 | n6997 ;
  assign n6999 = ( ~n6718 & n6907 ) | ( ~n6718 & n6996 ) | ( n6907 & n6996 ) ;
  assign n7000 = n6998 | n6999 ;
  assign n7001 = ~n6861 & n6918 ;
  assign n7002 = n6991 ^ n6961 ^ n6815 ;
  assign n7003 = n5851 & n6907 ;
  assign n7004 = ( n6733 & n6901 ) | ( n6733 & n7003 ) | ( n6901 & n7003 ) ;
  assign n7005 = n7003 | n7004 ;
  assign n7006 = ( ~n6685 & n6906 ) | ( ~n6685 & n7003 ) | ( n6906 & n7003 ) ;
  assign n7007 = n7005 | n7006 ;
  assign n7008 = n6256 & n6901 ;
  assign n7009 = n7001 | n7007 ;
  assign n7010 = ( n5851 & n6906 ) | ( n5851 & n7008 ) | ( n6906 & n7008 ) ;
  assign n7011 = n7008 | n7010 ;
  assign n7012 = n7009 ^ x29 ^ 1'b0 ;
  assign n7013 = ( ~n6617 & n6907 ) | ( ~n6617 & n7008 ) | ( n6907 & n7008 ) ;
  assign n7014 = n7011 | n7013 ;
  assign n7015 = n7012 ^ n6994 ^ n6832 ;
  assign n7016 = ( n6832 & n6994 ) | ( n6832 & n7012 ) | ( n6994 & n7012 ) ;
  assign n7017 = ( n6877 & n6918 ) | ( n6877 & n7000 ) | ( n6918 & n7000 ) ;
  assign n7018 = n6952 ^ x29 ^ 1'b0 ;
  assign n7019 = n7000 | n7017 ;
  assign n7020 = ~n6885 & n6918 ;
  assign n7021 = n7014 & ~n7020 ;
  assign n7022 = ( ~n6841 & n7016 ) | ( ~n6841 & n7018 ) | ( n7016 & n7018 ) ;
  assign n7023 = n7021 ^ n7020 ^ x29 ;
  assign n7024 = ( n6857 & n7022 ) | ( n6857 & n7023 ) | ( n7022 & n7023 ) ;
  assign n7025 = n7019 ^ x29 ^ 1'b0 ;
  assign n7026 = n7023 ^ n7022 ^ n6857 ;
  assign n7027 = n7018 ^ n7016 ^ n6841 ;
  assign n7028 = ( n6870 & n7024 ) | ( n6870 & n7025 ) | ( n7024 & n7025 ) ;
  assign n7029 = n7025 ^ n7024 ^ n6870 ;
  assign n7030 = x24 ^ x23 ^ 1'b0 ;
  assign n7031 = x26 ^ x25 ^ 1'b0 ;
  assign n7032 = n7030 | n7031 ;
  assign n7033 = x25 ^ x24 ^ 1'b0 ;
  assign n7034 = n7032 | n7033 ;
  assign n7035 = n7030 & n7031 ;
  assign n7036 = ~n7030 & n7033 ;
  assign n7037 = n7030 & ~n7031 ;
  assign n7038 = n6740 & n7036 ;
  assign n7039 = ~n6461 & n7037 ;
  assign n7040 = ( ~n6539 & n7036 ) | ( ~n6539 & n7039 ) | ( n7036 & n7039 ) ;
  assign n7041 = ~n6539 & n7030 ;
  assign n7042 = x26 & ~n7041 ;
  assign n7043 = ( n6962 & n7035 ) | ( n6962 & n7039 ) | ( n7035 & n7039 ) ;
  assign n7044 = ( ~n6668 & n7037 ) | ( ~n6668 & n7038 ) | ( n7037 & n7038 ) ;
  assign n7045 = n7039 | n7040 ;
  assign n7046 = n7043 | n7045 ;
  assign n7047 = n7046 ^ x26 ^ 1'b0 ;
  assign n7048 = n7047 ^ n7042 ^ 1'b0 ;
  assign n7049 = n7042 & n7047 ;
  assign n7050 = n6808 & n7035 ;
  assign n7051 = n7038 | n7044 ;
  assign n7052 = n7036 ^ n7034 ^ n7030 ;
  assign n7053 = ( ~n6461 & n7038 ) | ( ~n6461 & n7052 ) | ( n7038 & n7052 ) ;
  assign n7054 = n7051 | n7053 ;
  assign n7055 = n7050 | n7054 ;
  assign n7056 = ~n6461 & n7036 ;
  assign n7057 = ( ~n6539 & n7052 ) | ( ~n6539 & n7056 ) | ( n7052 & n7056 ) ;
  assign n7058 = n7056 | n7057 ;
  assign n7059 = ( n6740 & n7037 ) | ( n6740 & n7058 ) | ( n7037 & n7058 ) ;
  assign n7060 = n7058 | n7059 ;
  assign n7061 = ( n6798 & n7035 ) | ( n6798 & n7058 ) | ( n7035 & n7058 ) ;
  assign n7062 = n7060 | n7061 ;
  assign n7063 = n7062 ^ x26 ^ 1'b0 ;
  assign n7064 = n7055 ^ x26 ^ 1'b0 ;
  assign n7065 = n7049 & n7063 ;
  assign n7066 = n7063 ^ n7049 ^ 1'b0 ;
  assign n7067 = ( n6966 & n7064 ) | ( n6966 & n7065 ) | ( n7064 & n7065 ) ;
  assign n7068 = n7065 ^ n7064 ^ n6966 ;
  assign n7069 = n6740 & n7052 ;
  assign n7070 = ( ~n6735 & n7037 ) | ( ~n6735 & n7069 ) | ( n7037 & n7069 ) ;
  assign n7071 = n7069 | n7070 ;
  assign n7072 = ( ~n6668 & n7036 ) | ( ~n6668 & n7069 ) | ( n7036 & n7069 ) ;
  assign n7073 = n7071 | n7072 ;
  assign n7074 = ~n6811 & n7035 ;
  assign n7075 = n7073 & ~n7074 ;
  assign n7076 = n7075 ^ n7074 ^ x26 ;
  assign n7077 = n7076 ^ n7067 ^ n6973 ;
  assign n7078 = ( n6973 & n7067 ) | ( n6973 & n7076 ) | ( n7067 & n7076 ) ;
  assign n7079 = ~n6685 & n7037 ;
  assign n7080 = ( ~n6735 & n7036 ) | ( ~n6735 & n7079 ) | ( n7036 & n7079 ) ;
  assign n7081 = n7079 | n7080 ;
  assign n7082 = ( ~n6668 & n7052 ) | ( ~n6668 & n7079 ) | ( n7052 & n7079 ) ;
  assign n7083 = n7081 | n7082 ;
  assign n7084 = ~n6828 & n7035 ;
  assign n7085 = n7083 | n7084 ;
  assign n7086 = n7085 ^ x26 ^ 1'b0 ;
  assign n7087 = ( n6983 & n7078 ) | ( n6983 & n7086 ) | ( n7078 & n7086 ) ;
  assign n7088 = n7086 ^ n7078 ^ n6983 ;
  assign n7089 = n6733 & n7037 ;
  assign n7090 = ( ~n6685 & n7036 ) | ( ~n6685 & n7089 ) | ( n7036 & n7089 ) ;
  assign n7091 = n7089 | n7090 ;
  assign n7092 = ( ~n6735 & n7052 ) | ( ~n6735 & n7089 ) | ( n7052 & n7089 ) ;
  assign n7093 = n7091 | n7092 ;
  assign n7094 = n6843 & n7035 ;
  assign n7095 = n7093 | n7094 ;
  assign n7096 = n7095 ^ x26 ^ 1'b0 ;
  assign n7097 = ( n6975 & n7087 ) | ( n6975 & n7096 ) | ( n7087 & n7096 ) ;
  assign n7098 = n7096 ^ n7087 ^ n6975 ;
  assign n7099 = n5851 & n7037 ;
  assign n7100 = ( n6733 & n7036 ) | ( n6733 & n7099 ) | ( n7036 & n7099 ) ;
  assign n7101 = n7099 | n7100 ;
  assign n7102 = ( ~n6685 & n7052 ) | ( ~n6685 & n7099 ) | ( n7052 & n7099 ) ;
  assign n7103 = n7101 | n7102 ;
  assign n7104 = ~n6861 & n7035 ;
  assign n7105 = n7103 & ~n7104 ;
  assign n7106 = n7105 ^ n7104 ^ x26 ;
  assign n7107 = ( n6992 & n7097 ) | ( n6992 & n7106 ) | ( n7097 & n7106 ) ;
  assign n7108 = n7106 ^ n7097 ^ n6992 ;
  assign n7109 = n6256 & n7036 ;
  assign n7110 = ( n5851 & n7052 ) | ( n5851 & n7109 ) | ( n7052 & n7109 ) ;
  assign n7111 = n7109 | n7110 ;
  assign n7112 = n6256 & n7037 ;
  assign n7113 = ( ~n6617 & n7037 ) | ( ~n6617 & n7109 ) | ( n7037 & n7109 ) ;
  assign n7114 = ( n6733 & n7052 ) | ( n6733 & n7112 ) | ( n7052 & n7112 ) ;
  assign n7115 = ( n5851 & n7036 ) | ( n5851 & n7112 ) | ( n7036 & n7112 ) ;
  assign n7116 = n7112 | n7115 ;
  assign n7117 = ~n6885 & n7035 ;
  assign n7118 = n7111 | n7113 ;
  assign n7119 = ~n7117 & n7118 ;
  assign n7120 = n7114 | n7116 ;
  assign n7121 = ( ~n6603 & n6731 ) | ( ~n6603 & n6905 ) | ( n6731 & n6905 ) ;
  assign n7122 = ( n6858 & n7035 ) | ( n6858 & n7120 ) | ( n7035 & n7120 ) ;
  assign n7123 = n7119 ^ n7117 ^ x26 ;
  assign n7124 = n7120 | n7122 ;
  assign n7125 = n7121 ^ n6603 ^ n6602 ;
  assign n7126 = n7124 ^ x26 ^ 1'b0 ;
  assign n7127 = ( ~n7002 & n7107 ) | ( ~n7002 & n7126 ) | ( n7107 & n7126 ) ;
  assign n7128 = n7126 ^ n7107 ^ n7002 ;
  assign n7129 = n7127 ^ n7123 ^ n6995 ;
  assign n7130 = ( ~n6995 & n7123 ) | ( ~n6995 & n7127 ) | ( n7123 & n7127 ) ;
  assign n7131 = n6603 & n7052 ;
  assign n7132 = ( ~n6533 & n7037 ) | ( ~n6533 & n7131 ) | ( n7037 & n7131 ) ;
  assign n7133 = n7131 | n7132 ;
  assign n7134 = ( n6602 & ~n6603 ) | ( n6602 & n7121 ) | ( ~n6603 & n7121 ) ;
  assign n7135 = n7134 ^ n6602 ^ n6533 ;
  assign n7136 = ( ~n6602 & n7036 ) | ( ~n6602 & n7131 ) | ( n7036 & n7131 ) ;
  assign n7137 = n7133 | n7136 ;
  assign n7138 = n7035 & ~n7135 ;
  assign n7139 = n7137 | n7138 ;
  assign n7140 = n7139 ^ x26 ^ 1'b0 ;
  assign n7141 = ( n6929 & n7028 ) | ( n6929 & n7140 ) | ( n7028 & n7140 ) ;
  assign n7142 = n7140 ^ n7028 ^ n6929 ;
  assign n7143 = n6256 & n7052 ;
  assign n7144 = ( ~n6718 & n7037 ) | ( ~n6718 & n7143 ) | ( n7037 & n7143 ) ;
  assign n7145 = n7143 | n7144 ;
  assign n7146 = ( n6533 & n6602 ) | ( n6533 & n7134 ) | ( n6602 & n7134 ) ;
  assign n7147 = n6905 ^ n6731 ^ n6603 ;
  assign n7148 = ( ~n6617 & n7036 ) | ( ~n6617 & n7143 ) | ( n7036 & n7143 ) ;
  assign n7149 = n7145 | n7148 ;
  assign n7150 = ( n6877 & n7035 ) | ( n6877 & n7149 ) | ( n7035 & n7149 ) ;
  assign n7151 = n7149 | n7150 ;
  assign n7152 = n7151 ^ x26 ^ 1'b0 ;
  assign n7153 = n7152 ^ n7130 ^ n7015 ;
  assign n7154 = ( n7015 & n7130 ) | ( n7015 & n7152 ) | ( n7130 & n7152 ) ;
  assign n7155 = ~n6731 & n7037 ;
  assign n7156 = ( ~n6718 & n7036 ) | ( ~n6718 & n7155 ) | ( n7036 & n7155 ) ;
  assign n7157 = n7155 | n7156 ;
  assign n7158 = ( ~n6617 & n7052 ) | ( ~n6617 & n7155 ) | ( n7052 & n7155 ) ;
  assign n7159 = n7157 | n7158 ;
  assign n7160 = ~n6917 & n7035 ;
  assign n7161 = n7159 & ~n7160 ;
  assign n7162 = n7161 ^ n7160 ^ x26 ;
  assign n7163 = ( ~n7027 & n7154 ) | ( ~n7027 & n7162 ) | ( n7154 & n7162 ) ;
  assign n7164 = n7162 ^ n7154 ^ n7027 ;
  assign n7165 = n6603 & n7037 ;
  assign n7166 = ( ~n6731 & n7036 ) | ( ~n6731 & n7165 ) | ( n7036 & n7165 ) ;
  assign n7167 = n7165 | n7166 ;
  assign n7168 = ( ~n6718 & n7052 ) | ( ~n6718 & n7165 ) | ( n7052 & n7165 ) ;
  assign n7169 = n7167 | n7168 ;
  assign n7170 = ( n7035 & n7147 ) | ( n7035 & n7169 ) | ( n7147 & n7169 ) ;
  assign n7171 = n7169 | n7170 ;
  assign n7172 = n7171 ^ x26 ^ 1'b0 ;
  assign n7173 = ( n7026 & n7163 ) | ( n7026 & n7172 ) | ( n7163 & n7172 ) ;
  assign n7174 = n7172 ^ n7163 ^ n7026 ;
  assign n7175 = n6603 & n7036 ;
  assign n7176 = ( ~n6602 & n7037 ) | ( ~n6602 & n7175 ) | ( n7037 & n7175 ) ;
  assign n7177 = n7175 | n7176 ;
  assign n7178 = ( ~n6731 & n7052 ) | ( ~n6731 & n7175 ) | ( n7052 & n7175 ) ;
  assign n7179 = n7177 | n7178 ;
  assign n7180 = ( n7035 & n7125 ) | ( n7035 & n7179 ) | ( n7125 & n7179 ) ;
  assign n7181 = n7179 | n7180 ;
  assign n7182 = n7181 ^ x26 ^ 1'b0 ;
  assign n7183 = n7182 ^ n7173 ^ n7029 ;
  assign n7184 = ( n7029 & n7173 ) | ( n7029 & n7182 ) | ( n7173 & n7182 ) ;
  assign n7185 = x23 ^ x22 ^ 1'b0 ;
  assign n7186 = x22 ^ x21 ^ 1'b0 ;
  assign n7187 = x21 ^ x20 ^ 1'b0 ;
  assign n7188 = ~n7185 & n7187 ;
  assign n7189 = n7186 | n7187 ;
  assign n7190 = ( n7185 & n7188 ) | ( n7185 & ~n7189 ) | ( n7188 & ~n7189 ) ;
  assign n7191 = ~n6539 & n7187 ;
  assign n7192 = n7186 & ~n7187 ;
  assign n7193 = ~n6539 & n7190 ;
  assign n7194 = x23 & ~n7191 ;
  assign n7195 = ( ~n6461 & n7192 ) | ( ~n6461 & n7193 ) | ( n7192 & n7193 ) ;
  assign n7196 = n7185 & n7187 ;
  assign n7197 = n7193 | n7195 ;
  assign n7198 = ( n6798 & n7196 ) | ( n6798 & n7197 ) | ( n7196 & n7197 ) ;
  assign n7199 = ( n6740 & n7188 ) | ( n6740 & n7197 ) | ( n7188 & n7197 ) ;
  assign n7200 = n7197 | n7199 ;
  assign n7201 = n7198 | n7200 ;
  assign n7202 = n7201 ^ x23 ^ 1'b0 ;
  assign n7203 = n6740 & n7192 ;
  assign n7204 = ~n6461 & n7188 ;
  assign n7205 = ( n6962 & n7196 ) | ( n6962 & n7204 ) | ( n7196 & n7204 ) ;
  assign n7206 = n7204 | n7205 ;
  assign n7207 = ( ~n6539 & n7192 ) | ( ~n6539 & n7204 ) | ( n7192 & n7204 ) ;
  assign n7208 = n7206 | n7207 ;
  assign n7209 = n7208 ^ x23 ^ 1'b0 ;
  assign n7210 = n7209 ^ n7194 ^ 1'b0 ;
  assign n7211 = n7194 & n7209 ;
  assign n7212 = n7202 & n7211 ;
  assign n7213 = n7211 ^ n7202 ^ 1'b0 ;
  assign n7214 = ( ~n6668 & n7188 ) | ( ~n6668 & n7203 ) | ( n7188 & n7203 ) ;
  assign n7215 = n7203 | n7214 ;
  assign n7216 = ( ~n6461 & n7190 ) | ( ~n6461 & n7203 ) | ( n7190 & n7203 ) ;
  assign n7217 = n7215 | n7216 ;
  assign n7218 = n6808 & n7196 ;
  assign n7219 = n7217 | n7218 ;
  assign n7220 = n7219 ^ x23 ^ 1'b0 ;
  assign n7221 = n7220 ^ n7212 ^ n7041 ;
  assign n7222 = ( n7041 & n7212 ) | ( n7041 & n7220 ) | ( n7212 & n7220 ) ;
  assign n7223 = n6740 & n7190 ;
  assign n7224 = ( ~n6735 & n7188 ) | ( ~n6735 & n7223 ) | ( n7188 & n7223 ) ;
  assign n7225 = n7223 | n7224 ;
  assign n7226 = ( ~n6668 & n7192 ) | ( ~n6668 & n7223 ) | ( n7192 & n7223 ) ;
  assign n7227 = n7225 | n7226 ;
  assign n7228 = ~n6811 & n7196 ;
  assign n7229 = n7227 & ~n7228 ;
  assign n7230 = n7229 ^ n7228 ^ x23 ;
  assign n7231 = ( n7048 & n7222 ) | ( n7048 & n7230 ) | ( n7222 & n7230 ) ;
  assign n7232 = n7230 ^ n7222 ^ n7048 ;
  assign n7233 = ~n6685 & n7188 ;
  assign n7234 = ( ~n6668 & n7190 ) | ( ~n6668 & n7233 ) | ( n7190 & n7233 ) ;
  assign n7235 = n7233 | n7234 ;
  assign n7236 = ( ~n6735 & n7192 ) | ( ~n6735 & n7233 ) | ( n7192 & n7233 ) ;
  assign n7237 = n7235 | n7236 ;
  assign n7238 = ~n6828 & n7196 ;
  assign n7239 = n7237 | n7238 ;
  assign n7240 = n7239 ^ x23 ^ 1'b0 ;
  assign n7241 = ( n7066 & n7231 ) | ( n7066 & n7240 ) | ( n7231 & n7240 ) ;
  assign n7242 = n7240 ^ n7231 ^ n7066 ;
  assign n7243 = n6733 & n7188 ;
  assign n7244 = ( ~n6735 & n7190 ) | ( ~n6735 & n7243 ) | ( n7190 & n7243 ) ;
  assign n7245 = n7243 | n7244 ;
  assign n7246 = ( ~n6685 & n7192 ) | ( ~n6685 & n7243 ) | ( n7192 & n7243 ) ;
  assign n7247 = n7245 | n7246 ;
  assign n7248 = ( n6843 & n7196 ) | ( n6843 & n7247 ) | ( n7196 & n7247 ) ;
  assign n7249 = n7247 | n7248 ;
  assign n7250 = n7249 ^ x23 ^ 1'b0 ;
  assign n7251 = ( n7068 & n7241 ) | ( n7068 & n7250 ) | ( n7241 & n7250 ) ;
  assign n7252 = n7250 ^ n7241 ^ n7068 ;
  assign n7253 = n5851 & n7188 ;
  assign n7254 = ( n6733 & n7192 ) | ( n6733 & n7253 ) | ( n7192 & n7253 ) ;
  assign n7255 = n7253 | n7254 ;
  assign n7256 = ( ~n6685 & n7190 ) | ( ~n6685 & n7253 ) | ( n7190 & n7253 ) ;
  assign n7257 = n7255 | n7256 ;
  assign n7258 = ~n6861 & n7196 ;
  assign n7259 = n7257 | n7258 ;
  assign n7260 = n7259 ^ x23 ^ 1'b0 ;
  assign n7261 = ( n7077 & n7251 ) | ( n7077 & n7260 ) | ( n7251 & n7260 ) ;
  assign n7262 = n7260 ^ n7251 ^ n7077 ;
  assign n7263 = n6256 & n7188 ;
  assign n7264 = n6256 & n7192 ;
  assign n7265 = ( n5851 & n7190 ) | ( n5851 & n7264 ) | ( n7190 & n7264 ) ;
  assign n7266 = ( ~n6617 & n7188 ) | ( ~n6617 & n7264 ) | ( n7188 & n7264 ) ;
  assign n7267 = n7264 | n7265 ;
  assign n7268 = n7266 | n7267 ;
  assign n7269 = ~n6885 & n7196 ;
  assign n7270 = ( n5851 & n7192 ) | ( n5851 & n7263 ) | ( n7192 & n7263 ) ;
  assign n7271 = n7263 | n7270 ;
  assign n7272 = ( n6733 & n7190 ) | ( n6733 & n7263 ) | ( n7190 & n7263 ) ;
  assign n7273 = n7271 | n7272 ;
  assign n7274 = ( n6858 & n7196 ) | ( n6858 & n7273 ) | ( n7196 & n7273 ) ;
  assign n7275 = ~n6917 & n7196 ;
  assign n7276 = n7273 | n7274 ;
  assign n7277 = n7276 ^ x23 ^ 1'b0 ;
  assign n7278 = n7268 & ~n7269 ;
  assign n7279 = n7278 ^ n7269 ^ x23 ;
  assign n7280 = ( n7088 & n7261 ) | ( n7088 & n7277 ) | ( n7261 & n7277 ) ;
  assign n7281 = ( n7098 & n7279 ) | ( n7098 & n7280 ) | ( n7279 & n7280 ) ;
  assign n7282 = n7280 ^ n7279 ^ n7098 ;
  assign n7283 = n6603 & n7188 ;
  assign n7284 = ( ~n6718 & n7190 ) | ( ~n6718 & n7283 ) | ( n7190 & n7283 ) ;
  assign n7285 = n7283 | n7284 ;
  assign n7286 = ( ~n6731 & n7192 ) | ( ~n6731 & n7283 ) | ( n7192 & n7283 ) ;
  assign n7287 = n7277 ^ n7261 ^ n7088 ;
  assign n7288 = ~n6731 & n7188 ;
  assign n7289 = ( ~n6617 & n7190 ) | ( ~n6617 & n7288 ) | ( n7190 & n7288 ) ;
  assign n7290 = n7285 | n7286 ;
  assign n7291 = ( ~n6718 & n7192 ) | ( ~n6718 & n7288 ) | ( n7192 & n7288 ) ;
  assign n7292 = n7288 | n7289 ;
  assign n7293 = n7291 | n7292 ;
  assign n7294 = n7275 | n7293 ;
  assign n7295 = n6256 & n7190 ;
  assign n7296 = ( ~n6718 & n7188 ) | ( ~n6718 & n7295 ) | ( n7188 & n7295 ) ;
  assign n7297 = n7295 | n7296 ;
  assign n7298 = ( ~n6617 & n7192 ) | ( ~n6617 & n7295 ) | ( n7192 & n7295 ) ;
  assign n7299 = n7297 | n7298 ;
  assign n7300 = n6877 & n7196 ;
  assign n7301 = n7299 | n7300 ;
  assign n7302 = n7301 ^ x23 ^ 1'b0 ;
  assign n7303 = n7302 ^ n7281 ^ n7108 ;
  assign n7304 = n6603 & n7192 ;
  assign n7305 = ( n7108 & n7281 ) | ( n7108 & n7302 ) | ( n7281 & n7302 ) ;
  assign n7306 = ( ~n6602 & n7188 ) | ( ~n6602 & n7304 ) | ( n7188 & n7304 ) ;
  assign n7307 = n7304 | n7306 ;
  assign n7308 = ( ~n6731 & n7190 ) | ( ~n6731 & n7304 ) | ( n7190 & n7304 ) ;
  assign n7309 = n7294 ^ x23 ^ 1'b0 ;
  assign n7310 = n7147 & n7196 ;
  assign n7311 = n7290 | n7310 ;
  assign n7312 = n7309 ^ n7305 ^ n7128 ;
  assign n7313 = ( ~n7128 & n7305 ) | ( ~n7128 & n7309 ) | ( n7305 & n7309 ) ;
  assign n7314 = n7311 ^ x23 ^ 1'b0 ;
  assign n7315 = n7314 ^ n7313 ^ n7129 ;
  assign n7316 = n7125 & n7196 ;
  assign n7317 = n7307 | n7308 ;
  assign n7318 = ~n7135 & n7196 ;
  assign n7319 = n7316 | n7317 ;
  assign n7320 = ( ~n7129 & n7313 ) | ( ~n7129 & n7314 ) | ( n7313 & n7314 ) ;
  assign n7321 = n6603 & n7190 ;
  assign n7322 = ( ~n6602 & n7192 ) | ( ~n6602 & n7321 ) | ( n7192 & n7321 ) ;
  assign n7323 = n7319 ^ x23 ^ 1'b0 ;
  assign n7324 = ( ~n6533 & n7188 ) | ( ~n6533 & n7321 ) | ( n7188 & n7321 ) ;
  assign n7325 = n7321 | n7324 ;
  assign n7326 = n7322 | n7325 ;
  assign n7327 = n7323 ^ n7320 ^ n7153 ;
  assign n7328 = ( n7153 & n7320 ) | ( n7153 & n7323 ) | ( n7320 & n7323 ) ;
  assign n7329 = n7318 | n7326 ;
  assign n7330 = n7329 ^ x23 ^ 1'b0 ;
  assign n7331 = n7330 ^ n7328 ^ n7164 ;
  assign n7332 = ( ~n7164 & n7328 ) | ( ~n7164 & n7330 ) | ( n7328 & n7330 ) ;
  assign n7333 = x18 ^ x17 ^ 1'b0 ;
  assign n7334 = x19 ^ x18 ^ 1'b0 ;
  assign n7335 = x20 ^ x19 ^ 1'b0 ;
  assign n7336 = ~n7334 & n7335 ;
  assign n7337 = n7333 & ~n7335 ;
  assign n7338 = ~n7333 & n7336 ;
  assign n7339 = ~n7333 & n7334 ;
  assign n7340 = n7333 & n7335 ;
  assign n7341 = n6962 & n7340 ;
  assign n7342 = ( ~n6539 & n7339 ) | ( ~n6539 & n7341 ) | ( n7339 & n7341 ) ;
  assign n7343 = ( ~n6461 & n7337 ) | ( ~n6461 & n7341 ) | ( n7337 & n7341 ) ;
  assign n7344 = n7341 | n7342 ;
  assign n7345 = n7343 | n7344 ;
  assign n7346 = n7345 ^ x20 ^ 1'b0 ;
  assign n7347 = n6740 & n7339 ;
  assign n7348 = ~n6461 & n7339 ;
  assign n7349 = ( ~n6539 & n7338 ) | ( ~n6539 & n7348 ) | ( n7338 & n7348 ) ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = ( n6740 & n7337 ) | ( n6740 & n7350 ) | ( n7337 & n7350 ) ;
  assign n7352 = n7350 | n7351 ;
  assign n7353 = ~n6539 & n7333 ;
  assign n7354 = x20 & ~n7353 ;
  assign n7355 = ( n6798 & n7340 ) | ( n6798 & n7350 ) | ( n7340 & n7350 ) ;
  assign n7356 = n7352 | n7355 ;
  assign n7357 = n7354 ^ n7346 ^ 1'b0 ;
  assign n7358 = n7356 ^ x20 ^ 1'b0 ;
  assign n7359 = n7346 & n7354 ;
  assign n7360 = n7359 ^ n7358 ^ 1'b0 ;
  assign n7361 = n7358 & n7359 ;
  assign n7362 = ( ~n6668 & n7337 ) | ( ~n6668 & n7347 ) | ( n7337 & n7347 ) ;
  assign n7363 = n7347 | n7362 ;
  assign n7364 = ( ~n6461 & n7338 ) | ( ~n6461 & n7347 ) | ( n7338 & n7347 ) ;
  assign n7365 = n7363 | n7364 ;
  assign n7366 = n6808 & n7340 ;
  assign n7367 = n7365 | n7366 ;
  assign n7368 = n7367 ^ x20 ^ 1'b0 ;
  assign n7369 = ( n7191 & n7361 ) | ( n7191 & n7368 ) | ( n7361 & n7368 ) ;
  assign n7370 = n7368 ^ n7361 ^ n7191 ;
  assign n7371 = n6740 & n7338 ;
  assign n7372 = ( ~n6668 & n7339 ) | ( ~n6668 & n7371 ) | ( n7339 & n7371 ) ;
  assign n7373 = n7371 | n7372 ;
  assign n7374 = ( ~n6735 & n7337 ) | ( ~n6735 & n7371 ) | ( n7337 & n7371 ) ;
  assign n7375 = n7373 | n7374 ;
  assign n7376 = ~n6811 & n7340 ;
  assign n7377 = n7375 & ~n7376 ;
  assign n7378 = n7377 ^ n7376 ^ x20 ;
  assign n7379 = ( n7210 & n7369 ) | ( n7210 & n7378 ) | ( n7369 & n7378 ) ;
  assign n7380 = n7378 ^ n7369 ^ n7210 ;
  assign n7381 = ~n6735 & n7339 ;
  assign n7382 = ( ~n6685 & n7337 ) | ( ~n6685 & n7381 ) | ( n7337 & n7381 ) ;
  assign n7383 = n7381 | n7382 ;
  assign n7384 = ( ~n6668 & n7338 ) | ( ~n6668 & n7381 ) | ( n7338 & n7381 ) ;
  assign n7385 = n7383 | n7384 ;
  assign n7386 = ~n6828 & n7340 ;
  assign n7387 = n7385 | n7386 ;
  assign n7388 = n7387 ^ x20 ^ 1'b0 ;
  assign n7389 = n7388 ^ n7379 ^ n7213 ;
  assign n7390 = ( n7213 & n7379 ) | ( n7213 & n7388 ) | ( n7379 & n7388 ) ;
  assign n7391 = n6733 & n7337 ;
  assign n7392 = ( ~n6685 & n7339 ) | ( ~n6685 & n7391 ) | ( n7339 & n7391 ) ;
  assign n7393 = n7391 | n7392 ;
  assign n7394 = ( ~n6735 & n7338 ) | ( ~n6735 & n7391 ) | ( n7338 & n7391 ) ;
  assign n7395 = n7393 | n7394 ;
  assign n7396 = ( n6843 & n7340 ) | ( n6843 & n7395 ) | ( n7340 & n7395 ) ;
  assign n7397 = n7395 | n7396 ;
  assign n7398 = n7397 ^ x20 ^ 1'b0 ;
  assign n7399 = n7398 ^ n7390 ^ n7221 ;
  assign n7400 = ( n7221 & n7390 ) | ( n7221 & n7398 ) | ( n7390 & n7398 ) ;
  assign n7401 = n5851 & n7337 ;
  assign n7402 = ( n6733 & n7339 ) | ( n6733 & n7401 ) | ( n7339 & n7401 ) ;
  assign n7403 = n7401 | n7402 ;
  assign n7404 = ( ~n6685 & n7338 ) | ( ~n6685 & n7401 ) | ( n7338 & n7401 ) ;
  assign n7405 = n7403 | n7404 ;
  assign n7406 = ~n6861 & n7340 ;
  assign n7407 = n7405 | n7406 ;
  assign n7408 = n7407 ^ x20 ^ 1'b0 ;
  assign n7409 = n7408 ^ n7400 ^ n7232 ;
  assign n7410 = ( n7232 & n7400 ) | ( n7232 & n7408 ) | ( n7400 & n7408 ) ;
  assign n7411 = n6256 & n7337 ;
  assign n7412 = ( n5851 & n7339 ) | ( n5851 & n7411 ) | ( n7339 & n7411 ) ;
  assign n7413 = n7411 | n7412 ;
  assign n7414 = ( n6733 & n7338 ) | ( n6733 & n7411 ) | ( n7338 & n7411 ) ;
  assign n7415 = n7413 | n7414 ;
  assign n7416 = ( n6858 & n7340 ) | ( n6858 & n7415 ) | ( n7340 & n7415 ) ;
  assign n7417 = n7415 | n7416 ;
  assign n7418 = n7417 ^ x20 ^ 1'b0 ;
  assign n7419 = ( n7242 & n7410 ) | ( n7242 & n7418 ) | ( n7410 & n7418 ) ;
  assign n7420 = n7418 ^ n7410 ^ n7242 ;
  assign n7421 = n6256 & n7339 ;
  assign n7422 = ( n5851 & n7338 ) | ( n5851 & n7421 ) | ( n7338 & n7421 ) ;
  assign n7423 = n7421 | n7422 ;
  assign n7424 = ( ~n6617 & n7337 ) | ( ~n6617 & n7421 ) | ( n7337 & n7421 ) ;
  assign n7425 = n7423 | n7424 ;
  assign n7426 = ~n6885 & n7340 ;
  assign n7427 = n7425 & ~n7426 ;
  assign n7428 = n7427 ^ n7426 ^ x20 ;
  assign n7429 = ( n7252 & n7419 ) | ( n7252 & n7428 ) | ( n7419 & n7428 ) ;
  assign n7430 = n7428 ^ n7419 ^ n7252 ;
  assign n7431 = n6256 & n7338 ;
  assign n7432 = ( ~n6617 & n7339 ) | ( ~n6617 & n7431 ) | ( n7339 & n7431 ) ;
  assign n7433 = n7431 | n7432 ;
  assign n7434 = ( ~n6718 & n7337 ) | ( ~n6718 & n7431 ) | ( n7337 & n7431 ) ;
  assign n7435 = n7433 | n7434 ;
  assign n7436 = ( n6877 & n7340 ) | ( n6877 & n7435 ) | ( n7340 & n7435 ) ;
  assign n7437 = n7435 | n7436 ;
  assign n7438 = n7437 ^ x20 ^ 1'b0 ;
  assign n7439 = ( n7262 & n7429 ) | ( n7262 & n7438 ) | ( n7429 & n7438 ) ;
  assign n7440 = n7438 ^ n7429 ^ n7262 ;
  assign n7441 = ~n6718 & n7339 ;
  assign n7442 = ( ~n6731 & n7337 ) | ( ~n6731 & n7441 ) | ( n7337 & n7441 ) ;
  assign n7443 = n7441 | n7442 ;
  assign n7444 = ( ~n6617 & n7338 ) | ( ~n6617 & n7441 ) | ( n7338 & n7441 ) ;
  assign n7445 = n7443 | n7444 ;
  assign n7446 = ~n6917 & n7340 ;
  assign n7447 = n7445 | n7446 ;
  assign n7448 = n7447 ^ x20 ^ 1'b0 ;
  assign n7449 = ( n7287 & n7439 ) | ( n7287 & n7448 ) | ( n7439 & n7448 ) ;
  assign n7450 = n7448 ^ n7439 ^ n7287 ;
  assign n7451 = n6603 & n7337 ;
  assign n7452 = ( ~n6731 & n7339 ) | ( ~n6731 & n7451 ) | ( n7339 & n7451 ) ;
  assign n7453 = n7451 | n7452 ;
  assign n7454 = ( ~n6718 & n7338 ) | ( ~n6718 & n7451 ) | ( n7338 & n7451 ) ;
  assign n7455 = n7453 | n7454 ;
  assign n7456 = n7147 & n7340 ;
  assign n7457 = n7455 | n7456 ;
  assign n7458 = n7457 ^ x20 ^ 1'b0 ;
  assign n7459 = ( n7282 & n7449 ) | ( n7282 & n7458 ) | ( n7449 & n7458 ) ;
  assign n7460 = n7458 ^ n7449 ^ n7282 ;
  assign n7461 = n6603 & n7339 ;
  assign n7462 = ( ~n6602 & n7337 ) | ( ~n6602 & n7461 ) | ( n7337 & n7461 ) ;
  assign n7463 = n7461 | n7462 ;
  assign n7464 = ( ~n6731 & n7338 ) | ( ~n6731 & n7461 ) | ( n7338 & n7461 ) ;
  assign n7465 = n7463 | n7464 ;
  assign n7466 = ( n7125 & n7340 ) | ( n7125 & n7465 ) | ( n7340 & n7465 ) ;
  assign n7467 = n7465 | n7466 ;
  assign n7468 = n7467 ^ x20 ^ 1'b0 ;
  assign n7469 = n7468 ^ n7459 ^ n7303 ;
  assign n7470 = ( n7303 & n7459 ) | ( n7303 & n7468 ) | ( n7459 & n7468 ) ;
  assign n7471 = n6603 & n7338 ;
  assign n7472 = ( ~n6602 & n7339 ) | ( ~n6602 & n7471 ) | ( n7339 & n7471 ) ;
  assign n7473 = n7471 | n7472 ;
  assign n7474 = ( ~n6533 & n7337 ) | ( ~n6533 & n7471 ) | ( n7337 & n7471 ) ;
  assign n7475 = n7473 | n7474 ;
  assign n7476 = ~n7135 & n7340 ;
  assign n7477 = n7475 & ~n7476 ;
  assign n7478 = n7477 ^ n7476 ^ x20 ;
  assign n7479 = ( ~n7312 & n7470 ) | ( ~n7312 & n7478 ) | ( n7470 & n7478 ) ;
  assign n7480 = n7478 ^ n7470 ^ n7312 ;
  assign n7481 = x16 ^ x15 ^ 1'b0 ;
  assign n7482 = x17 ^ x16 ^ 1'b0 ;
  assign n7483 = x15 ^ x14 ^ 1'b0 ;
  assign n7484 = ~n6539 & n7483 ;
  assign n7485 = n7481 & ~n7483 ;
  assign n7486 = ~n7482 & n7483 ;
  assign n7487 = n7482 & n7483 ;
  assign n7488 = n6740 & n7485 ;
  assign n7489 = n6808 & n7487 ;
  assign n7490 = ( ~n6668 & n7486 ) | ( ~n6668 & n7488 ) | ( n7486 & n7488 ) ;
  assign n7491 = n7488 | n7490 ;
  assign n7492 = n7481 | n7483 ;
  assign n7493 = ( n7482 & n7486 ) | ( n7482 & ~n7492 ) | ( n7486 & ~n7492 ) ;
  assign n7494 = ~n6461 & n7485 ;
  assign n7495 = ( ~n6539 & n7493 ) | ( ~n6539 & n7494 ) | ( n7493 & n7494 ) ;
  assign n7496 = n7494 | n7495 ;
  assign n7497 = ( n6740 & n7486 ) | ( n6740 & n7496 ) | ( n7486 & n7496 ) ;
  assign n7498 = n7496 | n7497 ;
  assign n7499 = ( n6798 & n7487 ) | ( n6798 & n7496 ) | ( n7487 & n7496 ) ;
  assign n7500 = n7498 | n7499 ;
  assign n7501 = n7500 ^ x17 ^ 1'b0 ;
  assign n7502 = ( ~n6461 & n7488 ) | ( ~n6461 & n7493 ) | ( n7488 & n7493 ) ;
  assign n7503 = ~n6539 & n7485 ;
  assign n7504 = n7491 | n7502 ;
  assign n7505 = ( ~n6461 & n7486 ) | ( ~n6461 & n7503 ) | ( n7486 & n7503 ) ;
  assign n7506 = n7489 | n7504 ;
  assign n7507 = n7506 ^ x17 ^ 1'b0 ;
  assign n7508 = ( n6962 & n7487 ) | ( n6962 & n7503 ) | ( n7487 & n7503 ) ;
  assign n7509 = n7503 | n7508 ;
  assign n7510 = x17 & ~n7484 ;
  assign n7511 = n7505 | n7509 ;
  assign n7512 = n7511 ^ x17 ^ 1'b0 ;
  assign n7513 = n7512 ^ n7510 ^ 1'b0 ;
  assign n7514 = n7510 & n7512 ;
  assign n7515 = n7514 ^ n7501 ^ 1'b0 ;
  assign n7516 = n7501 & n7514 ;
  assign n7517 = ( n7353 & n7507 ) | ( n7353 & n7516 ) | ( n7507 & n7516 ) ;
  assign n7518 = n7516 ^ n7507 ^ n7353 ;
  assign n7519 = n6740 & n7493 ;
  assign n7520 = ( ~n6668 & n7485 ) | ( ~n6668 & n7519 ) | ( n7485 & n7519 ) ;
  assign n7521 = n7519 | n7520 ;
  assign n7522 = ( ~n6735 & n7486 ) | ( ~n6735 & n7519 ) | ( n7486 & n7519 ) ;
  assign n7523 = n7521 | n7522 ;
  assign n7524 = ~n6811 & n7487 ;
  assign n7525 = n7523 & ~n7524 ;
  assign n7526 = n7525 ^ n7524 ^ x17 ;
  assign n7527 = ( n7357 & n7517 ) | ( n7357 & n7526 ) | ( n7517 & n7526 ) ;
  assign n7528 = n7526 ^ n7517 ^ n7357 ;
  assign n7529 = ~n6735 & n7485 ;
  assign n7530 = ( ~n6685 & n7486 ) | ( ~n6685 & n7529 ) | ( n7486 & n7529 ) ;
  assign n7531 = n7529 | n7530 ;
  assign n7532 = ( ~n6668 & n7493 ) | ( ~n6668 & n7529 ) | ( n7493 & n7529 ) ;
  assign n7533 = n7531 | n7532 ;
  assign n7534 = ~n6828 & n7487 ;
  assign n7535 = n7533 | n7534 ;
  assign n7536 = n7535 ^ x17 ^ 1'b0 ;
  assign n7537 = ( n7360 & n7527 ) | ( n7360 & n7536 ) | ( n7527 & n7536 ) ;
  assign n7538 = n7536 ^ n7527 ^ n7360 ;
  assign n7539 = n6733 & n7486 ;
  assign n7540 = ( ~n6685 & n7485 ) | ( ~n6685 & n7539 ) | ( n7485 & n7539 ) ;
  assign n7541 = n7539 | n7540 ;
  assign n7542 = ( ~n6735 & n7493 ) | ( ~n6735 & n7539 ) | ( n7493 & n7539 ) ;
  assign n7543 = n7541 | n7542 ;
  assign n7544 = ( n6843 & n7487 ) | ( n6843 & n7543 ) | ( n7487 & n7543 ) ;
  assign n7545 = n7543 | n7544 ;
  assign n7546 = n7545 ^ x17 ^ 1'b0 ;
  assign n7547 = ( n7370 & n7537 ) | ( n7370 & n7546 ) | ( n7537 & n7546 ) ;
  assign n7548 = n7546 ^ n7537 ^ n7370 ;
  assign n7549 = n5851 & n7486 ;
  assign n7550 = ( n6733 & n7485 ) | ( n6733 & n7549 ) | ( n7485 & n7549 ) ;
  assign n7551 = n7549 | n7550 ;
  assign n7552 = ( ~n6685 & n7493 ) | ( ~n6685 & n7549 ) | ( n7493 & n7549 ) ;
  assign n7553 = n7551 | n7552 ;
  assign n7554 = ~n6861 & n7487 ;
  assign n7555 = n7553 | n7554 ;
  assign n7556 = n7555 ^ x17 ^ 1'b0 ;
  assign n7557 = ( n7380 & n7547 ) | ( n7380 & n7556 ) | ( n7547 & n7556 ) ;
  assign n7558 = n7556 ^ n7547 ^ n7380 ;
  assign n7559 = n6256 & n7486 ;
  assign n7560 = ( n5851 & n7485 ) | ( n5851 & n7559 ) | ( n7485 & n7559 ) ;
  assign n7561 = n7559 | n7560 ;
  assign n7562 = ( n6733 & n7493 ) | ( n6733 & n7559 ) | ( n7493 & n7559 ) ;
  assign n7563 = n7561 | n7562 ;
  assign n7564 = ( n6858 & n7487 ) | ( n6858 & n7563 ) | ( n7487 & n7563 ) ;
  assign n7565 = n7563 | n7564 ;
  assign n7566 = n7565 ^ x17 ^ 1'b0 ;
  assign n7567 = ( n7389 & n7557 ) | ( n7389 & n7566 ) | ( n7557 & n7566 ) ;
  assign n7568 = n7566 ^ n7557 ^ n7389 ;
  assign n7569 = n6256 & n7485 ;
  assign n7570 = ( n5851 & n7493 ) | ( n5851 & n7569 ) | ( n7493 & n7569 ) ;
  assign n7571 = n7569 | n7570 ;
  assign n7572 = ( ~n6617 & n7486 ) | ( ~n6617 & n7569 ) | ( n7486 & n7569 ) ;
  assign n7573 = n7571 | n7572 ;
  assign n7574 = ~n6885 & n7487 ;
  assign n7575 = n7573 & ~n7574 ;
  assign n7576 = n7575 ^ n7574 ^ x17 ;
  assign n7577 = n7576 ^ n7567 ^ n7399 ;
  assign n7578 = ( n7399 & n7567 ) | ( n7399 & n7576 ) | ( n7567 & n7576 ) ;
  assign n7579 = n6256 & n7493 ;
  assign n7580 = ( ~n6617 & n7485 ) | ( ~n6617 & n7579 ) | ( n7485 & n7579 ) ;
  assign n7581 = n7579 | n7580 ;
  assign n7582 = ( ~n6718 & n7486 ) | ( ~n6718 & n7579 ) | ( n7486 & n7579 ) ;
  assign n7583 = n7581 | n7582 ;
  assign n7584 = ( n6877 & n7487 ) | ( n6877 & n7583 ) | ( n7487 & n7583 ) ;
  assign n7585 = n7583 | n7584 ;
  assign n7586 = n7585 ^ x17 ^ 1'b0 ;
  assign n7587 = ( n7409 & n7578 ) | ( n7409 & n7586 ) | ( n7578 & n7586 ) ;
  assign n7588 = n7586 ^ n7578 ^ n7409 ;
  assign n7589 = ~n6718 & n7485 ;
  assign n7590 = ( ~n6731 & n7486 ) | ( ~n6731 & n7589 ) | ( n7486 & n7589 ) ;
  assign n7591 = n7589 | n7590 ;
  assign n7592 = ( ~n6617 & n7493 ) | ( ~n6617 & n7589 ) | ( n7493 & n7589 ) ;
  assign n7593 = n7591 | n7592 ;
  assign n7594 = ~n6917 & n7487 ;
  assign n7595 = n7593 | n7594 ;
  assign n7596 = n7595 ^ x17 ^ 1'b0 ;
  assign n7597 = ( n7420 & n7587 ) | ( n7420 & n7596 ) | ( n7587 & n7596 ) ;
  assign n7598 = n7596 ^ n7587 ^ n7420 ;
  assign n7599 = n6603 & n7486 ;
  assign n7600 = ( ~n6731 & n7485 ) | ( ~n6731 & n7599 ) | ( n7485 & n7599 ) ;
  assign n7601 = n7599 | n7600 ;
  assign n7602 = ( ~n6718 & n7493 ) | ( ~n6718 & n7599 ) | ( n7493 & n7599 ) ;
  assign n7603 = n7601 | n7602 ;
  assign n7604 = n7147 & n7487 ;
  assign n7605 = n7603 | n7604 ;
  assign n7606 = n7605 ^ x17 ^ 1'b0 ;
  assign n7607 = ( n7430 & n7597 ) | ( n7430 & n7606 ) | ( n7597 & n7606 ) ;
  assign n7608 = n7606 ^ n7597 ^ n7430 ;
  assign n7609 = n6603 & n7485 ;
  assign n7610 = ( ~n6602 & n7486 ) | ( ~n6602 & n7609 ) | ( n7486 & n7609 ) ;
  assign n7611 = n7609 | n7610 ;
  assign n7612 = ( ~n6731 & n7493 ) | ( ~n6731 & n7609 ) | ( n7493 & n7609 ) ;
  assign n7613 = n7611 | n7612 ;
  assign n7614 = n7125 & n7487 ;
  assign n7615 = n7613 | n7614 ;
  assign n7616 = n7615 ^ x17 ^ 1'b0 ;
  assign n7617 = ( n7440 & n7607 ) | ( n7440 & n7616 ) | ( n7607 & n7616 ) ;
  assign n7618 = n7616 ^ n7607 ^ n7440 ;
  assign n7619 = n6724 & n7188 ;
  assign n7620 = ( ~n6602 & n7190 ) | ( ~n6602 & n7619 ) | ( n7190 & n7619 ) ;
  assign n7621 = ( ~n6533 & n7192 ) | ( ~n6533 & n7619 ) | ( n7192 & n7619 ) ;
  assign n7622 = n7619 | n7620 ;
  assign n7623 = n7621 | n7622 ;
  assign n7624 = n7146 ^ n6724 ^ n6533 ;
  assign n7625 = n7196 & n7624 ;
  assign n7626 = n7623 | n7625 ;
  assign n7627 = n7626 ^ x23 ^ 1'b0 ;
  assign n7628 = n7627 ^ n7332 ^ n7174 ;
  assign n7629 = ( n7174 & n7332 ) | ( n7174 & n7627 ) | ( n7332 & n7627 ) ;
  assign n7630 = n6603 & n7493 ;
  assign n7631 = ( ~n6602 & n7485 ) | ( ~n6602 & n7630 ) | ( n7485 & n7630 ) ;
  assign n7632 = n7630 | n7631 ;
  assign n7633 = ( ~n6533 & n7486 ) | ( ~n6533 & n7630 ) | ( n7486 & n7630 ) ;
  assign n7634 = n7632 | n7633 ;
  assign n7635 = ~n7135 & n7487 ;
  assign n7636 = n7634 & ~n7635 ;
  assign n7637 = n7636 ^ n7635 ^ x17 ;
  assign n7638 = ( n7450 & n7617 ) | ( n7450 & n7637 ) | ( n7617 & n7637 ) ;
  assign n7639 = n7637 ^ n7617 ^ n7450 ;
  assign n7640 = n6724 & n7337 ;
  assign n7641 = ( ~n6533 & n7339 ) | ( ~n6533 & n7640 ) | ( n7339 & n7640 ) ;
  assign n7642 = n7640 | n7641 ;
  assign n7643 = ( ~n6602 & n7338 ) | ( ~n6602 & n7640 ) | ( n7338 & n7640 ) ;
  assign n7644 = n7642 | n7643 ;
  assign n7645 = ( n7340 & n7624 ) | ( n7340 & n7644 ) | ( n7624 & n7644 ) ;
  assign n7646 = n7644 | n7645 ;
  assign n7647 = n7646 ^ x20 ^ 1'b0 ;
  assign n7648 = n7647 ^ n7479 ^ n7315 ;
  assign n7649 = ( ~n7315 & n7479 ) | ( ~n7315 & n7647 ) | ( n7479 & n7647 ) ;
  assign n7650 = n6724 & n7486 ;
  assign n7651 = ( ~n6533 & n7485 ) | ( ~n6533 & n7650 ) | ( n7485 & n7650 ) ;
  assign n7652 = n7650 | n7651 ;
  assign n7653 = ( n6533 & ~n6724 ) | ( n6533 & n7146 ) | ( ~n6724 & n7146 ) ;
  assign n7654 = ( ~n6602 & n7493 ) | ( ~n6602 & n7650 ) | ( n7493 & n7650 ) ;
  assign n7655 = n7652 | n7654 ;
  assign n7656 = ( n7487 & n7624 ) | ( n7487 & n7655 ) | ( n7624 & n7655 ) ;
  assign n7657 = n7655 | n7656 ;
  assign n7658 = n7657 ^ x17 ^ 1'b0 ;
  assign n7659 = n7658 ^ n7638 ^ n7460 ;
  assign n7660 = ( n7460 & n7638 ) | ( n7460 & n7658 ) | ( n7638 & n7658 ) ;
  assign n7661 = x14 ^ x13 ^ 1'b0 ;
  assign n7662 = x13 ^ x12 ^ 1'b0 ;
  assign n7663 = x12 ^ x11 ^ 1'b0 ;
  assign n7664 = n7662 | n7663 ;
  assign n7665 = n7661 | n7664 ;
  assign n7666 = n7661 & n7663 ;
  assign n7667 = ~n7661 & n7663 ;
  assign n7668 = n6733 & n7667 ;
  assign n7669 = n7662 & ~n7663 ;
  assign n7670 = ( ~n6685 & n7668 ) | ( ~n6685 & n7669 ) | ( n7668 & n7669 ) ;
  assign n7671 = n7668 | n7670 ;
  assign n7672 = n6808 & n7666 ;
  assign n7673 = n6740 & n7669 ;
  assign n7674 = n7669 ^ n7665 ^ n7663 ;
  assign n7675 = ( ~n6461 & n7673 ) | ( ~n6461 & n7674 ) | ( n7673 & n7674 ) ;
  assign n7676 = n7673 | n7675 ;
  assign n7677 = ( ~n6668 & n7667 ) | ( ~n6668 & n7673 ) | ( n7667 & n7673 ) ;
  assign n7678 = n7676 | n7677 ;
  assign n7679 = n7672 | n7678 ;
  assign n7680 = n7679 ^ x14 ^ 1'b0 ;
  assign n7681 = ( ~n6735 & n7668 ) | ( ~n6735 & n7674 ) | ( n7668 & n7674 ) ;
  assign n7682 = n7671 | n7681 ;
  assign n7683 = ( n6843 & n7666 ) | ( n6843 & n7682 ) | ( n7666 & n7682 ) ;
  assign n7684 = n7682 | n7683 ;
  assign n7685 = n6740 & n7674 ;
  assign n7686 = ( ~n6668 & n7669 ) | ( ~n6668 & n7685 ) | ( n7669 & n7685 ) ;
  assign n7687 = n7685 | n7686 ;
  assign n7688 = ( ~n6735 & n7667 ) | ( ~n6735 & n7685 ) | ( n7667 & n7685 ) ;
  assign n7689 = n7684 ^ x14 ^ 1'b0 ;
  assign n7690 = ~n6461 & n7669 ;
  assign n7691 = n7687 | n7688 ;
  assign n7692 = ~n6811 & n7666 ;
  assign n7693 = n7691 & ~n7692 ;
  assign n7694 = n7693 ^ n7692 ^ x14 ;
  assign n7695 = ( ~n6539 & n7674 ) | ( ~n6539 & n7690 ) | ( n7674 & n7690 ) ;
  assign n7696 = n7690 | n7695 ;
  assign n7697 = ( n6740 & n7667 ) | ( n6740 & n7696 ) | ( n7667 & n7696 ) ;
  assign n7698 = n7696 | n7697 ;
  assign n7699 = ( n6798 & n7666 ) | ( n6798 & n7696 ) | ( n7666 & n7696 ) ;
  assign n7700 = n7698 | n7699 ;
  assign n7701 = n7700 ^ x14 ^ 1'b0 ;
  assign n7702 = ~n6539 & n7669 ;
  assign n7703 = ( ~n6461 & n7667 ) | ( ~n6461 & n7702 ) | ( n7667 & n7702 ) ;
  assign n7704 = ( n6962 & n7666 ) | ( n6962 & n7702 ) | ( n7666 & n7702 ) ;
  assign n7705 = n7702 | n7704 ;
  assign n7706 = n7703 | n7705 ;
  assign n7707 = n7706 ^ x14 ^ 1'b0 ;
  assign n7708 = ~n6539 & n7663 ;
  assign n7709 = x14 & ~n7708 ;
  assign n7710 = n7709 ^ n7707 ^ 1'b0 ;
  assign n7711 = n7707 & n7709 ;
  assign n7712 = n7701 & n7711 ;
  assign n7713 = n7711 ^ n7701 ^ 1'b0 ;
  assign n7714 = ( n7484 & n7680 ) | ( n7484 & n7712 ) | ( n7680 & n7712 ) ;
  assign n7715 = n7712 ^ n7680 ^ n7484 ;
  assign n7716 = ~n6735 & n7669 ;
  assign n7717 = ( ~n6668 & n7674 ) | ( ~n6668 & n7716 ) | ( n7674 & n7716 ) ;
  assign n7718 = n7716 | n7717 ;
  assign n7719 = ( ~n6685 & n7667 ) | ( ~n6685 & n7716 ) | ( n7667 & n7716 ) ;
  assign n7720 = n7718 | n7719 ;
  assign n7721 = ( n7513 & n7694 ) | ( n7513 & n7714 ) | ( n7694 & n7714 ) ;
  assign n7722 = n7714 ^ n7694 ^ n7513 ;
  assign n7723 = n5851 & n7667 ;
  assign n7724 = ( n6733 & n7669 ) | ( n6733 & n7723 ) | ( n7669 & n7723 ) ;
  assign n7725 = n7723 | n7724 ;
  assign n7726 = ( ~n6685 & n7674 ) | ( ~n6685 & n7723 ) | ( n7674 & n7723 ) ;
  assign n7727 = n7725 | n7726 ;
  assign n7728 = ~n6828 & n7666 ;
  assign n7729 = n7720 | n7728 ;
  assign n7730 = n7729 ^ x14 ^ 1'b0 ;
  assign n7731 = n7730 ^ n7721 ^ n7515 ;
  assign n7732 = ( n7515 & n7721 ) | ( n7515 & n7730 ) | ( n7721 & n7730 ) ;
  assign n7733 = n6256 & n7667 ;
  assign n7734 = ( n5851 & n7669 ) | ( n5851 & n7733 ) | ( n7669 & n7733 ) ;
  assign n7735 = n7733 | n7734 ;
  assign n7736 = ( n6733 & n7674 ) | ( n6733 & n7733 ) | ( n7674 & n7733 ) ;
  assign n7737 = n7735 | n7736 ;
  assign n7738 = ( n6858 & n7666 ) | ( n6858 & n7737 ) | ( n7666 & n7737 ) ;
  assign n7739 = n7737 | n7738 ;
  assign n7740 = n7739 ^ x14 ^ 1'b0 ;
  assign n7741 = ~n6861 & n7666 ;
  assign n7742 = n7727 | n7741 ;
  assign n7743 = n7732 ^ n7689 ^ n7518 ;
  assign n7744 = ( n7518 & n7689 ) | ( n7518 & n7732 ) | ( n7689 & n7732 ) ;
  assign n7745 = n7742 ^ x14 ^ 1'b0 ;
  assign n7746 = ( n7528 & n7744 ) | ( n7528 & n7745 ) | ( n7744 & n7745 ) ;
  assign n7747 = ( n7538 & n7740 ) | ( n7538 & n7746 ) | ( n7740 & n7746 ) ;
  assign n7748 = n7746 ^ n7740 ^ n7538 ;
  assign n7749 = n7745 ^ n7744 ^ n7528 ;
  assign n7750 = n6256 & n7669 ;
  assign n7751 = ( n5851 & n7674 ) | ( n5851 & n7750 ) | ( n7674 & n7750 ) ;
  assign n7752 = n7750 | n7751 ;
  assign n7753 = ( ~n6617 & n7667 ) | ( ~n6617 & n7750 ) | ( n7667 & n7750 ) ;
  assign n7754 = n7752 | n7753 ;
  assign n7755 = ~n6885 & n7666 ;
  assign n7756 = n7754 & ~n7755 ;
  assign n7757 = n7756 ^ n7755 ^ x14 ;
  assign n7758 = n7757 ^ n7747 ^ n7548 ;
  assign n7759 = ( n7548 & n7747 ) | ( n7548 & n7757 ) | ( n7747 & n7757 ) ;
  assign n7760 = n6256 & n7674 ;
  assign n7761 = ( ~n6617 & n7669 ) | ( ~n6617 & n7760 ) | ( n7669 & n7760 ) ;
  assign n7762 = n7760 | n7761 ;
  assign n7763 = ( ~n6718 & n7667 ) | ( ~n6718 & n7760 ) | ( n7667 & n7760 ) ;
  assign n7764 = n7762 | n7763 ;
  assign n7765 = ( n6877 & n7666 ) | ( n6877 & n7764 ) | ( n7666 & n7764 ) ;
  assign n7766 = n7764 | n7765 ;
  assign n7767 = n7766 ^ x14 ^ 1'b0 ;
  assign n7768 = n7767 ^ n7759 ^ n7558 ;
  assign n7769 = ( n7558 & n7759 ) | ( n7558 & n7767 ) | ( n7759 & n7767 ) ;
  assign n7770 = ~n6718 & n7669 ;
  assign n7771 = ( ~n6617 & n7674 ) | ( ~n6617 & n7770 ) | ( n7674 & n7770 ) ;
  assign n7772 = n7770 | n7771 ;
  assign n7773 = ( ~n6731 & n7667 ) | ( ~n6731 & n7770 ) | ( n7667 & n7770 ) ;
  assign n7774 = n7772 | n7773 ;
  assign n7775 = ~n6917 & n7666 ;
  assign n7776 = n7774 | n7775 ;
  assign n7777 = n7776 ^ x14 ^ 1'b0 ;
  assign n7778 = ( n7568 & n7769 ) | ( n7568 & n7777 ) | ( n7769 & n7777 ) ;
  assign n7779 = n7777 ^ n7769 ^ n7568 ;
  assign n7780 = n6603 & n7667 ;
  assign n7781 = ( ~n6731 & n7669 ) | ( ~n6731 & n7780 ) | ( n7669 & n7780 ) ;
  assign n7782 = n7780 | n7781 ;
  assign n7783 = ( ~n6718 & n7674 ) | ( ~n6718 & n7780 ) | ( n7674 & n7780 ) ;
  assign n7784 = n7782 | n7783 ;
  assign n7785 = n7147 & n7666 ;
  assign n7786 = n7784 | n7785 ;
  assign n7787 = n7786 ^ x14 ^ 1'b0 ;
  assign n7788 = ( n7577 & n7778 ) | ( n7577 & n7787 ) | ( n7778 & n7787 ) ;
  assign n7789 = n7787 ^ n7778 ^ n7577 ;
  assign n7790 = n6603 & n7669 ;
  assign n7791 = ( ~n6731 & n7674 ) | ( ~n6731 & n7790 ) | ( n7674 & n7790 ) ;
  assign n7792 = n7790 | n7791 ;
  assign n7793 = ( ~n6602 & n7667 ) | ( ~n6602 & n7790 ) | ( n7667 & n7790 ) ;
  assign n7794 = n7792 | n7793 ;
  assign n7795 = n7125 & n7666 ;
  assign n7796 = n7794 | n7795 ;
  assign n7797 = n7796 ^ x14 ^ 1'b0 ;
  assign n7798 = n7797 ^ n7788 ^ n7588 ;
  assign n7799 = ( n7588 & n7788 ) | ( n7588 & n7797 ) | ( n7788 & n7797 ) ;
  assign n7800 = n6603 & n7674 ;
  assign n7801 = ( ~n6602 & n7669 ) | ( ~n6602 & n7800 ) | ( n7669 & n7800 ) ;
  assign n7802 = n7800 | n7801 ;
  assign n7803 = ( ~n6533 & n7667 ) | ( ~n6533 & n7800 ) | ( n7667 & n7800 ) ;
  assign n7804 = n7802 | n7803 ;
  assign n7805 = ( ~n7135 & n7666 ) | ( ~n7135 & n7804 ) | ( n7666 & n7804 ) ;
  assign n7806 = n7804 | n7805 ;
  assign n7807 = n7806 ^ x14 ^ 1'b0 ;
  assign n7808 = n7807 ^ n7799 ^ n7598 ;
  assign n7809 = ( n7598 & n7799 ) | ( n7598 & n7807 ) | ( n7799 & n7807 ) ;
  assign n7810 = n6724 & n7667 ;
  assign n7811 = ( ~n6533 & n7669 ) | ( ~n6533 & n7810 ) | ( n7669 & n7810 ) ;
  assign n7812 = n7810 | n7811 ;
  assign n7813 = ( ~n6602 & n7674 ) | ( ~n6602 & n7810 ) | ( n7674 & n7810 ) ;
  assign n7814 = n7812 | n7813 ;
  assign n7815 = ( n7624 & n7666 ) | ( n7624 & n7814 ) | ( n7666 & n7814 ) ;
  assign n7816 = n7814 | n7815 ;
  assign n7817 = n7816 ^ x14 ^ 1'b0 ;
  assign n7818 = ( n7608 & n7809 ) | ( n7608 & n7817 ) | ( n7809 & n7817 ) ;
  assign n7819 = n7817 ^ n7809 ^ n7608 ;
  assign n7820 = n6789 & n7125 ;
  assign n7821 = ( n6603 & n6791 ) | ( n6603 & n7820 ) | ( n6791 & n7820 ) ;
  assign n7822 = n7820 | n7821 ;
  assign n7823 = ( ~n6731 & n6790 ) | ( ~n6731 & n7820 ) | ( n6790 & n7820 ) ;
  assign n7824 = n7822 | n7823 ;
  assign n7825 = n6602 & n6788 ;
  assign n7826 = ( n6788 & n7824 ) | ( n6788 & ~n7825 ) | ( n7824 & ~n7825 ) ;
  assign n7827 = x9 ^ x8 ^ 1'b0 ;
  assign n7828 = x10 ^ x9 ^ 1'b0 ;
  assign n7829 = ~n7827 & n7828 ;
  assign n7830 = n7827 | n7828 ;
  assign n7831 = x11 ^ x10 ^ 1'b0 ;
  assign n7832 = n7830 | n7831 ;
  assign n7833 = n7832 ^ n7829 ^ n7827 ;
  assign n7834 = n7827 & ~n7831 ;
  assign n7835 = ~n6461 & n7829 ;
  assign n7836 = ( ~n6539 & n7833 ) | ( ~n6539 & n7835 ) | ( n7833 & n7835 ) ;
  assign n7837 = n7835 | n7836 ;
  assign n7838 = n7827 & n7831 ;
  assign n7839 = ( n6798 & n7837 ) | ( n6798 & n7838 ) | ( n7837 & n7838 ) ;
  assign n7840 = n6962 & n7838 ;
  assign n7841 = ( ~n6539 & n7829 ) | ( ~n6539 & n7840 ) | ( n7829 & n7840 ) ;
  assign n7842 = n7840 | n7841 ;
  assign n7843 = ( n6740 & n7834 ) | ( n6740 & n7837 ) | ( n7834 & n7837 ) ;
  assign n7844 = n7837 | n7843 ;
  assign n7845 = n7839 | n7844 ;
  assign n7846 = n7845 ^ x11 ^ 1'b0 ;
  assign n7847 = ( ~n6461 & n7834 ) | ( ~n6461 & n7840 ) | ( n7834 & n7840 ) ;
  assign n7848 = n6740 & n7829 ;
  assign n7849 = ( ~n6461 & n7833 ) | ( ~n6461 & n7848 ) | ( n7833 & n7848 ) ;
  assign n7850 = n7842 | n7847 ;
  assign n7851 = n7850 ^ x11 ^ 1'b0 ;
  assign n7852 = ~n6539 & n7827 ;
  assign n7853 = n7848 | n7849 ;
  assign n7854 = x11 & ~n7852 ;
  assign n7855 = ( ~n6668 & n7834 ) | ( ~n6668 & n7848 ) | ( n7834 & n7848 ) ;
  assign n7856 = n7853 | n7855 ;
  assign n7857 = n6808 & n7838 ;
  assign n7858 = n7856 | n7857 ;
  assign n7859 = n7858 ^ x11 ^ 1'b0 ;
  assign n7860 = n7854 ^ n7851 ^ 1'b0 ;
  assign n7861 = n7851 & n7854 ;
  assign n7862 = n7846 & n7861 ;
  assign n7863 = n7861 ^ n7846 ^ 1'b0 ;
  assign n7864 = ( n7708 & n7859 ) | ( n7708 & n7862 ) | ( n7859 & n7862 ) ;
  assign n7865 = n7862 ^ n7859 ^ n7708 ;
  assign n7866 = n6740 & n7833 ;
  assign n7867 = ( ~n6668 & n7829 ) | ( ~n6668 & n7866 ) | ( n7829 & n7866 ) ;
  assign n7868 = n7866 | n7867 ;
  assign n7869 = ( ~n6735 & n7834 ) | ( ~n6735 & n7866 ) | ( n7834 & n7866 ) ;
  assign n7870 = n7868 | n7869 ;
  assign n7871 = ( ~n6811 & n7838 ) | ( ~n6811 & n7870 ) | ( n7838 & n7870 ) ;
  assign n7872 = n7870 | n7871 ;
  assign n7873 = n7872 ^ x11 ^ 1'b0 ;
  assign n7874 = n7873 ^ n7864 ^ n7710 ;
  assign n7875 = ( n7710 & n7864 ) | ( n7710 & n7873 ) | ( n7864 & n7873 ) ;
  assign n7876 = ~n6735 & n7829 ;
  assign n7877 = ( ~n6668 & n7833 ) | ( ~n6668 & n7876 ) | ( n7833 & n7876 ) ;
  assign n7878 = n7876 | n7877 ;
  assign n7879 = ( ~n6685 & n7834 ) | ( ~n6685 & n7876 ) | ( n7834 & n7876 ) ;
  assign n7880 = n7878 | n7879 ;
  assign n7881 = ~n6828 & n7838 ;
  assign n7882 = n7880 | n7881 ;
  assign n7883 = n7882 ^ x11 ^ 1'b0 ;
  assign n7884 = ( n7713 & n7875 ) | ( n7713 & n7883 ) | ( n7875 & n7883 ) ;
  assign n7885 = n7883 ^ n7875 ^ n7713 ;
  assign n7886 = n6733 & n7834 ;
  assign n7887 = ( ~n6685 & n7829 ) | ( ~n6685 & n7886 ) | ( n7829 & n7886 ) ;
  assign n7888 = n7886 | n7887 ;
  assign n7889 = ( ~n6735 & n7833 ) | ( ~n6735 & n7886 ) | ( n7833 & n7886 ) ;
  assign n7890 = n7888 | n7889 ;
  assign n7891 = ( n6843 & n7838 ) | ( n6843 & n7890 ) | ( n7838 & n7890 ) ;
  assign n7892 = n7890 | n7891 ;
  assign n7893 = n7892 ^ x11 ^ 1'b0 ;
  assign n7894 = ( n7715 & n7884 ) | ( n7715 & n7893 ) | ( n7884 & n7893 ) ;
  assign n7895 = n7893 ^ n7884 ^ n7715 ;
  assign n7896 = n5851 & n7834 ;
  assign n7897 = ( n6733 & n7829 ) | ( n6733 & n7896 ) | ( n7829 & n7896 ) ;
  assign n7898 = n7896 | n7897 ;
  assign n7899 = ( ~n6685 & n7833 ) | ( ~n6685 & n7896 ) | ( n7833 & n7896 ) ;
  assign n7900 = n7898 | n7899 ;
  assign n7901 = ~n6861 & n7838 ;
  assign n7902 = n7900 | n7901 ;
  assign n7903 = n7902 ^ x11 ^ 1'b0 ;
  assign n7904 = n7903 ^ n7894 ^ n7722 ;
  assign n7905 = ( n7722 & n7894 ) | ( n7722 & n7903 ) | ( n7894 & n7903 ) ;
  assign n7906 = n6256 & n7834 ;
  assign n7907 = ( n5851 & n7829 ) | ( n5851 & n7906 ) | ( n7829 & n7906 ) ;
  assign n7908 = n7906 | n7907 ;
  assign n7909 = ( n6733 & n7833 ) | ( n6733 & n7906 ) | ( n7833 & n7906 ) ;
  assign n7910 = n7908 | n7909 ;
  assign n7911 = ( n6858 & n7838 ) | ( n6858 & n7910 ) | ( n7838 & n7910 ) ;
  assign n7912 = n7910 | n7911 ;
  assign n7913 = n7912 ^ x11 ^ 1'b0 ;
  assign n7914 = n7913 ^ n7905 ^ n7731 ;
  assign n7915 = ( n7731 & n7905 ) | ( n7731 & n7913 ) | ( n7905 & n7913 ) ;
  assign n7916 = n6256 & n7829 ;
  assign n7917 = ( n5851 & n7833 ) | ( n5851 & n7916 ) | ( n7833 & n7916 ) ;
  assign n7918 = n7916 | n7917 ;
  assign n7919 = ( ~n6617 & n7834 ) | ( ~n6617 & n7916 ) | ( n7834 & n7916 ) ;
  assign n7920 = n7918 | n7919 ;
  assign n7921 = ( ~n6885 & n7838 ) | ( ~n6885 & n7920 ) | ( n7838 & n7920 ) ;
  assign n7922 = n7920 | n7921 ;
  assign n7923 = n7922 ^ x11 ^ 1'b0 ;
  assign n7924 = ( n7743 & n7915 ) | ( n7743 & n7923 ) | ( n7915 & n7923 ) ;
  assign n7925 = n7923 ^ n7915 ^ n7743 ;
  assign n7926 = x7 ^ x6 ^ 1'b0 ;
  assign n7927 = x6 ^ x5 ^ 1'b0 ;
  assign n7928 = x8 ^ x7 ^ 1'b0 ;
  assign n7929 = n7927 & ~n7928 ;
  assign n7930 = n7927 & n7928 ;
  assign n7931 = n6962 & n7930 ;
  assign n7932 = n7926 & ~n7927 ;
  assign n7933 = ( ~n6461 & n7929 ) | ( ~n6461 & n7931 ) | ( n7929 & n7931 ) ;
  assign n7934 = ( ~n6539 & n7931 ) | ( ~n6539 & n7932 ) | ( n7931 & n7932 ) ;
  assign n7935 = n7931 | n7934 ;
  assign n7936 = n7933 | n7935 ;
  assign n7937 = n7936 ^ x8 ^ 1'b0 ;
  assign n7938 = n6740 & n7932 ;
  assign n7939 = ~n6539 & n7927 ;
  assign n7940 = x8 & ~n7939 ;
  assign n7941 = n7926 | n7927 ;
  assign n7942 = n7928 | n7941 ;
  assign n7943 = n7942 ^ n7932 ^ n7927 ;
  assign n7944 = n7940 ^ n7937 ^ 1'b0 ;
  assign n7945 = ( ~n6461 & n7938 ) | ( ~n6461 & n7943 ) | ( n7938 & n7943 ) ;
  assign n7946 = n7938 | n7945 ;
  assign n7947 = ( ~n6668 & n7929 ) | ( ~n6668 & n7938 ) | ( n7929 & n7938 ) ;
  assign n7948 = n7946 | n7947 ;
  assign n7949 = n7937 & n7940 ;
  assign n7950 = ~n6461 & n7932 ;
  assign n7951 = ( ~n6539 & n7943 ) | ( ~n6539 & n7950 ) | ( n7943 & n7950 ) ;
  assign n7952 = n7950 | n7951 ;
  assign n7953 = ( n6740 & n7929 ) | ( n6740 & n7952 ) | ( n7929 & n7952 ) ;
  assign n7954 = n7952 | n7953 ;
  assign n7955 = ( n6798 & n7930 ) | ( n6798 & n7952 ) | ( n7930 & n7952 ) ;
  assign n7956 = n7954 | n7955 ;
  assign n7957 = n7956 ^ x8 ^ 1'b0 ;
  assign n7958 = n7957 ^ n7949 ^ 1'b0 ;
  assign n7959 = n7949 & n7957 ;
  assign n7960 = n6808 & n7930 ;
  assign n7961 = n7948 | n7960 ;
  assign n7962 = n7961 ^ x8 ^ 1'b0 ;
  assign n7963 = ( n7852 & n7959 ) | ( n7852 & n7962 ) | ( n7959 & n7962 ) ;
  assign n7964 = n7962 ^ n7959 ^ n7852 ;
  assign n7965 = n6740 & n7943 ;
  assign n7966 = ( ~n6668 & n7932 ) | ( ~n6668 & n7965 ) | ( n7932 & n7965 ) ;
  assign n7967 = n7965 | n7966 ;
  assign n7968 = ( ~n6735 & n7929 ) | ( ~n6735 & n7965 ) | ( n7929 & n7965 ) ;
  assign n7969 = n7967 | n7968 ;
  assign n7970 = ( ~n6811 & n7930 ) | ( ~n6811 & n7969 ) | ( n7930 & n7969 ) ;
  assign n7971 = n7969 | n7970 ;
  assign n7972 = n7971 ^ x8 ^ 1'b0 ;
  assign n7973 = n7972 ^ n7963 ^ n7860 ;
  assign n7974 = ( n7860 & n7963 ) | ( n7860 & n7972 ) | ( n7963 & n7972 ) ;
  assign n7975 = ~n6735 & n7932 ;
  assign n7976 = ( ~n6668 & n7943 ) | ( ~n6668 & n7975 ) | ( n7943 & n7975 ) ;
  assign n7977 = n7975 | n7976 ;
  assign n7978 = ( ~n6685 & n7929 ) | ( ~n6685 & n7975 ) | ( n7929 & n7975 ) ;
  assign n7979 = n7977 | n7978 ;
  assign n7980 = ~n6828 & n7930 ;
  assign n7981 = n7979 | n7980 ;
  assign n7982 = n7981 ^ x8 ^ 1'b0 ;
  assign n7983 = ( n7863 & n7974 ) | ( n7863 & n7982 ) | ( n7974 & n7982 ) ;
  assign n7984 = n7982 ^ n7974 ^ n7863 ;
  assign n7985 = n6733 & n7929 ;
  assign n7986 = ( ~n6685 & n7932 ) | ( ~n6685 & n7985 ) | ( n7932 & n7985 ) ;
  assign n7987 = n7985 | n7986 ;
  assign n7988 = ( ~n6735 & n7943 ) | ( ~n6735 & n7985 ) | ( n7943 & n7985 ) ;
  assign n7989 = n7987 | n7988 ;
  assign n7990 = ( n6843 & n7930 ) | ( n6843 & n7989 ) | ( n7930 & n7989 ) ;
  assign n7991 = n7989 | n7990 ;
  assign n7992 = n7991 ^ x8 ^ 1'b0 ;
  assign n7993 = ( n7865 & n7983 ) | ( n7865 & n7992 ) | ( n7983 & n7992 ) ;
  assign n7994 = n7992 ^ n7983 ^ n7865 ;
  assign n7995 = n5851 & n7929 ;
  assign n7996 = ( n6733 & n7932 ) | ( n6733 & n7995 ) | ( n7932 & n7995 ) ;
  assign n7997 = n7995 | n7996 ;
  assign n7998 = ( ~n6685 & n7943 ) | ( ~n6685 & n7995 ) | ( n7943 & n7995 ) ;
  assign n7999 = n7997 | n7998 ;
  assign n8000 = ~n6861 & n7930 ;
  assign n8001 = n7999 | n8000 ;
  assign n8002 = n8001 ^ x8 ^ 1'b0 ;
  assign n8003 = n8002 ^ n7993 ^ n7874 ;
  assign n8004 = ( n7874 & n7993 ) | ( n7874 & n8002 ) | ( n7993 & n8002 ) ;
  assign n8005 = n6256 & n7929 ;
  assign n8006 = ( n5851 & n7932 ) | ( n5851 & n8005 ) | ( n7932 & n8005 ) ;
  assign n8007 = n8005 | n8006 ;
  assign n8008 = ( n6733 & n7943 ) | ( n6733 & n8005 ) | ( n7943 & n8005 ) ;
  assign n8009 = n8007 | n8008 ;
  assign n8010 = ( n6858 & n7930 ) | ( n6858 & n8009 ) | ( n7930 & n8009 ) ;
  assign n8011 = n8009 | n8010 ;
  assign n8012 = n8011 ^ x8 ^ 1'b0 ;
  assign n8013 = n8012 ^ n8004 ^ n7885 ;
  assign n8014 = ( n7885 & n8004 ) | ( n7885 & n8012 ) | ( n8004 & n8012 ) ;
  assign n8015 = n6256 & n7932 ;
  assign n8016 = ( n5851 & n7943 ) | ( n5851 & n8015 ) | ( n7943 & n8015 ) ;
  assign n8017 = n8015 | n8016 ;
  assign n8018 = ( ~n6617 & n7929 ) | ( ~n6617 & n8015 ) | ( n7929 & n8015 ) ;
  assign n8019 = n8017 | n8018 ;
  assign n8020 = ( ~n6885 & n7930 ) | ( ~n6885 & n8019 ) | ( n7930 & n8019 ) ;
  assign n8021 = n8019 | n8020 ;
  assign n8022 = n8021 ^ x8 ^ 1'b0 ;
  assign n8023 = ( n7895 & n8014 ) | ( n7895 & n8022 ) | ( n8014 & n8022 ) ;
  assign n8024 = n8022 ^ n8014 ^ n7895 ;
  assign n8025 = x3 ^ x2 ^ 1'b0 ;
  assign n8026 = x5 ^ x4 ^ 1'b0 ;
  assign n8027 = n8025 | n8026 ;
  assign n8028 = x4 ^ x3 ^ 1'b0 ;
  assign n8029 = ~n8025 & n8028 ;
  assign n8030 = n8027 | n8028 ;
  assign n8031 = ~n6461 & n8029 ;
  assign n8032 = ~n6539 & n8025 ;
  assign n8033 = n8025 & ~n8026 ;
  assign n8034 = n8025 & n8026 ;
  assign n8035 = n6962 & n8034 ;
  assign n8036 = ( ~n6539 & n8029 ) | ( ~n6539 & n8035 ) | ( n8029 & n8035 ) ;
  assign n8037 = n8030 ^ n8029 ^ n8025 ;
  assign n8038 = n6740 & n8029 ;
  assign n8039 = n8035 | n8036 ;
  assign n8040 = ( ~n6539 & n8031 ) | ( ~n6539 & n8037 ) | ( n8031 & n8037 ) ;
  assign n8041 = n8031 | n8040 ;
  assign n8042 = ( ~n6461 & n8033 ) | ( ~n6461 & n8035 ) | ( n8033 & n8035 ) ;
  assign n8043 = n8039 | n8042 ;
  assign n8044 = x5 & ~n8032 ;
  assign n8045 = n8043 ^ x5 ^ 1'b0 ;
  assign n8046 = n8044 & n8045 ;
  assign n8047 = n8045 ^ n8044 ^ 1'b0 ;
  assign n8048 = ( ~n6461 & n8037 ) | ( ~n6461 & n8038 ) | ( n8037 & n8038 ) ;
  assign n8049 = n8038 | n8048 ;
  assign n8050 = ( ~n6668 & n8033 ) | ( ~n6668 & n8038 ) | ( n8033 & n8038 ) ;
  assign n8051 = n8049 | n8050 ;
  assign n8052 = ( n6740 & n8033 ) | ( n6740 & n8041 ) | ( n8033 & n8041 ) ;
  assign n8053 = n8041 | n8052 ;
  assign n8054 = ( n6798 & n8034 ) | ( n6798 & n8041 ) | ( n8034 & n8041 ) ;
  assign n8055 = n8053 | n8054 ;
  assign n8056 = n6808 & n8034 ;
  assign n8057 = n8051 | n8056 ;
  assign n8058 = n8055 ^ x5 ^ 1'b0 ;
  assign n8059 = n8046 & n8058 ;
  assign n8060 = n8058 ^ n8046 ^ 1'b0 ;
  assign n8061 = n8057 ^ x5 ^ 1'b0 ;
  assign n8062 = n8061 ^ n8059 ^ n7939 ;
  assign n8063 = ( n7939 & n8059 ) | ( n7939 & n8061 ) | ( n8059 & n8061 ) ;
  assign n8064 = n6740 & n8037 ;
  assign n8065 = ( ~n6668 & n8029 ) | ( ~n6668 & n8064 ) | ( n8029 & n8064 ) ;
  assign n8066 = n8064 | n8065 ;
  assign n8067 = ( ~n6735 & n8033 ) | ( ~n6735 & n8064 ) | ( n8033 & n8064 ) ;
  assign n8068 = n8066 | n8067 ;
  assign n8069 = ( ~n6811 & n8034 ) | ( ~n6811 & n8068 ) | ( n8034 & n8068 ) ;
  assign n8070 = n8068 | n8069 ;
  assign n8071 = n8070 ^ x5 ^ 1'b0 ;
  assign n8072 = ( n7944 & n8063 ) | ( n7944 & n8071 ) | ( n8063 & n8071 ) ;
  assign n8073 = n8071 ^ n8063 ^ n7944 ;
  assign n8074 = ~n6735 & n8029 ;
  assign n8075 = ( ~n6668 & n8037 ) | ( ~n6668 & n8074 ) | ( n8037 & n8074 ) ;
  assign n8076 = n8074 | n8075 ;
  assign n8077 = ( ~n6685 & n8033 ) | ( ~n6685 & n8074 ) | ( n8033 & n8074 ) ;
  assign n8078 = n8076 | n8077 ;
  assign n8079 = ~n6828 & n8034 ;
  assign n8080 = n8078 | n8079 ;
  assign n8081 = n8080 ^ x5 ^ 1'b0 ;
  assign n8082 = n8081 ^ n8072 ^ n7958 ;
  assign n8083 = ( n7958 & n8072 ) | ( n7958 & n8081 ) | ( n8072 & n8081 ) ;
  assign n8084 = x0 | x1 ;
  assign n8085 = x2 ^ x1 ^ 1'b0 ;
  assign n8086 = ~n8084 & n8085 ;
  assign n8087 = n6740 & n8086 ;
  assign n8088 = ~x0 & x1 ;
  assign n8089 = x0 & n8085 ;
  assign n8090 = x0 & ~n8085 ;
  assign n8091 = ( ~n6668 & n8087 ) | ( ~n6668 & n8088 ) | ( n8087 & n8088 ) ;
  assign n8092 = n8087 | n8091 ;
  assign n8093 = ( ~n6735 & n8087 ) | ( ~n6735 & n8090 ) | ( n8087 & n8090 ) ;
  assign n8094 = n8092 | n8093 ;
  assign n8095 = ( ~n6811 & n8089 ) | ( ~n6811 & n8094 ) | ( n8089 & n8094 ) ;
  assign n8096 = n8094 | n8095 ;
  assign n8097 = n6740 & n8088 ;
  assign n8098 = ( ~n6461 & n8086 ) | ( ~n6461 & n8097 ) | ( n8086 & n8097 ) ;
  assign n8099 = n8097 | n8098 ;
  assign n8100 = ( ~n6668 & n8090 ) | ( ~n6668 & n8097 ) | ( n8090 & n8097 ) ;
  assign n8101 = n8099 | n8100 ;
  assign n8102 = n6808 & n8089 ;
  assign n8103 = n8101 | n8102 ;
  assign n8104 = n6740 & n8090 ;
  assign n8105 = ~n6828 & n8089 ;
  assign n8106 = ~n6668 & n8086 ;
  assign n8107 = ( ~n6735 & n8088 ) | ( ~n6735 & n8106 ) | ( n8088 & n8106 ) ;
  assign n8108 = n8106 | n8107 ;
  assign n8109 = ( ~n6685 & n8090 ) | ( ~n6685 & n8106 ) | ( n8090 & n8106 ) ;
  assign n8110 = n8108 | n8109 ;
  assign n8111 = n8105 | n8110 ;
  assign n8112 = ( ~n6461 & n8088 ) | ( ~n6461 & n8104 ) | ( n8088 & n8104 ) ;
  assign n8113 = x2 & n8088 ;
  assign n8114 = ( ~n6539 & n8086 ) | ( ~n6539 & n8104 ) | ( n8086 & n8104 ) ;
  assign n8115 = n8104 | n8114 ;
  assign n8116 = ( x2 & n6539 ) | ( x2 & ~n8113 ) | ( n6539 & ~n8113 ) ;
  assign n8117 = x0 & ~n6539 ;
  assign n8118 = n8111 ^ x2 ^ 1'b0 ;
  assign n8119 = n8112 | n8115 ;
  assign n8120 = x2 & n8089 ;
  assign n8121 = n6798 & n8120 ;
  assign n8122 = ( x2 & n6461 ) | ( x2 & ~n8090 ) | ( n6461 & ~n8090 ) ;
  assign n8123 = x2 & n8122 ;
  assign n8124 = n8116 & n8123 ;
  assign n8125 = n6962 & n8120 ;
  assign n8126 = ( ~n8121 & n8124 ) | ( ~n8121 & n8125 ) | ( n8124 & n8125 ) ;
  assign n8127 = ( x2 & n8119 ) | ( x2 & n8121 ) | ( n8119 & n8121 ) ;
  assign n8128 = ~n8125 & n8126 ;
  assign n8129 = ( ~n8117 & n8127 ) | ( ~n8117 & n8128 ) | ( n8127 & n8128 ) ;
  assign n8130 = ~n8127 & n8129 ;
  assign n8131 = n8103 ^ x2 ^ 1'b0 ;
  assign n8132 = ( n8032 & n8130 ) | ( n8032 & n8131 ) | ( n8130 & n8131 ) ;
  assign n8133 = n8096 ^ x2 ^ 1'b0 ;
  assign n8134 = ( n8047 & n8132 ) | ( n8047 & n8133 ) | ( n8132 & n8133 ) ;
  assign n8135 = ( n8060 & n8118 ) | ( n8060 & n8134 ) | ( n8118 & n8134 ) ;
  assign n8136 = n6733 & n8090 ;
  assign n8137 = ( ~n6735 & n8086 ) | ( ~n6735 & n8136 ) | ( n8086 & n8136 ) ;
  assign n8138 = n8136 | n8137 ;
  assign n8139 = ( ~n6685 & n8088 ) | ( ~n6685 & n8136 ) | ( n8088 & n8136 ) ;
  assign n8140 = n8138 | n8139 ;
  assign n8141 = ( n6843 & n8089 ) | ( n6843 & n8140 ) | ( n8089 & n8140 ) ;
  assign n8142 = n8140 | n8141 ;
  assign n8143 = n8142 ^ x2 ^ 1'b0 ;
  assign n8144 = n5851 & n8033 ;
  assign n8145 = ( n8062 & n8135 ) | ( n8062 & n8143 ) | ( n8135 & n8143 ) ;
  assign n8146 = ( n6733 & n8029 ) | ( n6733 & n8144 ) | ( n8029 & n8144 ) ;
  assign n8147 = n8144 | n8146 ;
  assign n8148 = ~n6861 & n8034 ;
  assign n8149 = ( ~n6685 & n8037 ) | ( ~n6685 & n8144 ) | ( n8037 & n8144 ) ;
  assign n8150 = n8147 | n8149 ;
  assign n8151 = n8148 | n8150 ;
  assign n8152 = n5851 & n8090 ;
  assign n8153 = ( n6733 & n8088 ) | ( n6733 & n8152 ) | ( n8088 & n8152 ) ;
  assign n8154 = n8152 | n8153 ;
  assign n8155 = ( ~n6685 & n8086 ) | ( ~n6685 & n8152 ) | ( n8086 & n8152 ) ;
  assign n8156 = n8154 | n8155 ;
  assign n8157 = n6733 & n8033 ;
  assign n8158 = ~n6861 & n8089 ;
  assign n8159 = n8156 | n8158 ;
  assign n8160 = n8159 ^ x2 ^ 1'b0 ;
  assign n8161 = ( ~n6735 & n8037 ) | ( ~n6735 & n8157 ) | ( n8037 & n8157 ) ;
  assign n8162 = ( ~n6685 & n8029 ) | ( ~n6685 & n8157 ) | ( n8029 & n8157 ) ;
  assign n8163 = ( n8073 & n8145 ) | ( n8073 & n8160 ) | ( n8145 & n8160 ) ;
  assign n8164 = n6256 & n8090 ;
  assign n8165 = ( n5851 & n8088 ) | ( n5851 & n8164 ) | ( n8088 & n8164 ) ;
  assign n8166 = n8164 | n8165 ;
  assign n8167 = ( n6733 & n8086 ) | ( n6733 & n8164 ) | ( n8086 & n8164 ) ;
  assign n8168 = n6256 & n8033 ;
  assign n8169 = ( n6733 & n8037 ) | ( n6733 & n8168 ) | ( n8037 & n8168 ) ;
  assign n8170 = n8157 | n8162 ;
  assign n8171 = n8161 | n8170 ;
  assign n8172 = ( n6843 & n8034 ) | ( n6843 & n8171 ) | ( n8034 & n8171 ) ;
  assign n8173 = ( n5851 & n8029 ) | ( n5851 & n8168 ) | ( n8029 & n8168 ) ;
  assign n8174 = n8168 | n8173 ;
  assign n8175 = n8151 ^ x5 ^ 1'b0 ;
  assign n8176 = n8171 | n8172 ;
  assign n8177 = n8176 ^ x5 ^ 1'b0 ;
  assign n8178 = ( n7964 & n8083 ) | ( n7964 & n8177 ) | ( n8083 & n8177 ) ;
  assign n8179 = n8177 ^ n8083 ^ n7964 ;
  assign n8180 = ( n7973 & n8175 ) | ( n7973 & n8178 ) | ( n8175 & n8178 ) ;
  assign n8181 = n8166 | n8167 ;
  assign n8182 = ( n6858 & n8089 ) | ( n6858 & n8181 ) | ( n8089 & n8181 ) ;
  assign n8183 = n8181 | n8182 ;
  assign n8184 = n8183 ^ x2 ^ 1'b0 ;
  assign n8185 = n8178 ^ n8175 ^ n7973 ;
  assign n8186 = n8169 | n8174 ;
  assign n8187 = ( n6858 & n8034 ) | ( n6858 & n8186 ) | ( n8034 & n8186 ) ;
  assign n8188 = n8186 | n8187 ;
  assign n8189 = n8188 ^ x5 ^ 1'b0 ;
  assign n8190 = ( n8082 & n8163 ) | ( n8082 & n8184 ) | ( n8163 & n8184 ) ;
  assign n8191 = n8189 ^ n8180 ^ n7984 ;
  assign n8192 = ( n7984 & n8180 ) | ( n7984 & n8189 ) | ( n8180 & n8189 ) ;
  assign n8193 = n6256 & n8088 ;
  assign n8194 = ( n5851 & n8086 ) | ( n5851 & n8193 ) | ( n8086 & n8193 ) ;
  assign n8195 = n8193 | n8194 ;
  assign n8196 = ( ~n6617 & n8090 ) | ( ~n6617 & n8193 ) | ( n8090 & n8193 ) ;
  assign n8197 = n8195 | n8196 ;
  assign n8198 = ( ~n6885 & n8089 ) | ( ~n6885 & n8197 ) | ( n8089 & n8197 ) ;
  assign n8199 = n8197 | n8198 ;
  assign n8200 = n6256 & n8086 ;
  assign n8201 = n8199 ^ x2 ^ 1'b0 ;
  assign n8202 = ( n8179 & n8190 ) | ( n8179 & n8201 ) | ( n8190 & n8201 ) ;
  assign n8203 = ( ~n6617 & n8088 ) | ( ~n6617 & n8200 ) | ( n8088 & n8200 ) ;
  assign n8204 = ( ~n6718 & n8090 ) | ( ~n6718 & n8200 ) | ( n8090 & n8200 ) ;
  assign n8205 = n8200 | n8203 ;
  assign n8206 = n8204 | n8205 ;
  assign n8207 = ( n6877 & n8089 ) | ( n6877 & n8206 ) | ( n8089 & n8206 ) ;
  assign n8208 = n8206 | n8207 ;
  assign n8209 = ~n6617 & n8086 ;
  assign n8210 = ( ~n6718 & n8088 ) | ( ~n6718 & n8209 ) | ( n8088 & n8209 ) ;
  assign n8211 = n8209 | n8210 ;
  assign n8212 = ( ~n6731 & n8090 ) | ( ~n6731 & n8209 ) | ( n8090 & n8209 ) ;
  assign n8213 = n8208 ^ x2 ^ 1'b0 ;
  assign n8214 = ( n8185 & n8202 ) | ( n8185 & n8213 ) | ( n8202 & n8213 ) ;
  assign n8215 = n6256 & n8029 ;
  assign n8216 = n6603 & n8090 ;
  assign n8217 = n8211 | n8212 ;
  assign n8218 = ( n5851 & n8037 ) | ( n5851 & n8215 ) | ( n8037 & n8215 ) ;
  assign n8219 = ( ~n6617 & n8033 ) | ( ~n6617 & n8215 ) | ( n8033 & n8215 ) ;
  assign n8220 = n8215 | n8218 ;
  assign n8221 = ~n6917 & n8089 ;
  assign n8222 = n8217 | n8221 ;
  assign n8223 = n8222 ^ x2 ^ 1'b0 ;
  assign n8224 = n7147 & n8089 ;
  assign n8225 = ( n8191 & n8214 ) | ( n8191 & n8223 ) | ( n8214 & n8223 ) ;
  assign n8226 = ( ~n6718 & n8086 ) | ( ~n6718 & n8216 ) | ( n8086 & n8216 ) ;
  assign n8227 = n8216 | n8226 ;
  assign n8228 = n8219 | n8220 ;
  assign n8229 = ( ~n6885 & n8034 ) | ( ~n6885 & n8228 ) | ( n8034 & n8228 ) ;
  assign n8230 = n8228 | n8229 ;
  assign n8231 = ( ~n6731 & n8088 ) | ( ~n6731 & n8216 ) | ( n8088 & n8216 ) ;
  assign n8232 = n8230 ^ x5 ^ 1'b0 ;
  assign n8233 = n8227 | n8231 ;
  assign n8234 = ( n7994 & n8192 ) | ( n7994 & n8232 ) | ( n8192 & n8232 ) ;
  assign n8235 = n8224 | n8233 ;
  assign n8236 = n8235 ^ x2 ^ 1'b0 ;
  assign n8237 = n8232 ^ n8192 ^ n7994 ;
  assign n8238 = ( n8225 & n8236 ) | ( n8225 & n8237 ) | ( n8236 & n8237 ) ;
  assign n8239 = n6256 & n8037 ;
  assign n8240 = ( ~n6617 & n8029 ) | ( ~n6617 & n8239 ) | ( n8029 & n8239 ) ;
  assign n8241 = n8239 | n8240 ;
  assign n8242 = ( ~n6718 & n8033 ) | ( ~n6718 & n8239 ) | ( n8033 & n8239 ) ;
  assign n8243 = n8241 | n8242 ;
  assign n8244 = ( n6877 & n8034 ) | ( n6877 & n8243 ) | ( n8034 & n8243 ) ;
  assign n8245 = n8243 | n8244 ;
  assign n8246 = n8245 ^ x5 ^ 1'b0 ;
  assign n8247 = n8246 ^ n8234 ^ n8003 ;
  assign n8248 = ( n8003 & n8234 ) | ( n8003 & n8246 ) | ( n8234 & n8246 ) ;
  assign n8249 = n6603 & n8088 ;
  assign n8250 = ( ~n6731 & n8086 ) | ( ~n6731 & n8249 ) | ( n8086 & n8249 ) ;
  assign n8251 = n8249 | n8250 ;
  assign n8252 = ( ~n6602 & n8090 ) | ( ~n6602 & n8249 ) | ( n8090 & n8249 ) ;
  assign n8253 = n8251 | n8252 ;
  assign n8254 = n7125 & n8089 ;
  assign n8255 = n8253 | n8254 ;
  assign n8256 = n8255 ^ x2 ^ 1'b0 ;
  assign n8257 = n6256 & n7833 ;
  assign n8258 = ( n8238 & n8247 ) | ( n8238 & n8256 ) | ( n8247 & n8256 ) ;
  assign n8259 = ( ~n6617 & n7829 ) | ( ~n6617 & n8257 ) | ( n7829 & n8257 ) ;
  assign n8260 = n8257 | n8259 ;
  assign n8261 = ( ~n6718 & n7834 ) | ( ~n6718 & n8257 ) | ( n7834 & n8257 ) ;
  assign n8262 = ~n6718 & n8029 ;
  assign n8263 = n8260 | n8261 ;
  assign n8264 = ( ~n6617 & n8037 ) | ( ~n6617 & n8262 ) | ( n8037 & n8262 ) ;
  assign n8265 = n8262 | n8264 ;
  assign n8266 = ( ~n6731 & n8033 ) | ( ~n6731 & n8262 ) | ( n8033 & n8262 ) ;
  assign n8267 = n6256 & n7943 ;
  assign n8268 = n8265 | n8266 ;
  assign n8269 = ( ~n6617 & n7932 ) | ( ~n6617 & n8267 ) | ( n7932 & n8267 ) ;
  assign n8270 = n8267 | n8269 ;
  assign n8271 = ( ~n6718 & n7929 ) | ( ~n6718 & n8267 ) | ( n7929 & n8267 ) ;
  assign n8272 = n8270 | n8271 ;
  assign n8273 = ( n6877 & n7930 ) | ( n6877 & n8272 ) | ( n7930 & n8272 ) ;
  assign n8274 = n8272 | n8273 ;
  assign n8275 = n6603 & n8086 ;
  assign n8276 = n8274 ^ x8 ^ 1'b0 ;
  assign n8277 = ( n6877 & n7838 ) | ( n6877 & n8263 ) | ( n7838 & n8263 ) ;
  assign n8278 = n8263 | n8277 ;
  assign n8279 = ~n6917 & n8034 ;
  assign n8280 = n8268 | n8279 ;
  assign n8281 = ( n7904 & n8023 ) | ( n7904 & n8276 ) | ( n8023 & n8276 ) ;
  assign n8282 = n8280 ^ x5 ^ 1'b0 ;
  assign n8283 = n8276 ^ n8023 ^ n7904 ;
  assign n8284 = n8282 ^ n8248 ^ n8013 ;
  assign n8285 = ( n8013 & n8248 ) | ( n8013 & n8282 ) | ( n8248 & n8282 ) ;
  assign n8286 = ( ~n6602 & n8088 ) | ( ~n6602 & n8275 ) | ( n8088 & n8275 ) ;
  assign n8287 = n8275 | n8286 ;
  assign n8288 = n8278 ^ x11 ^ 1'b0 ;
  assign n8289 = ( ~n6533 & n8090 ) | ( ~n6533 & n8275 ) | ( n8090 & n8275 ) ;
  assign n8290 = n8287 | n8289 ;
  assign n8291 = ( ~n7135 & n8089 ) | ( ~n7135 & n8290 ) | ( n8089 & n8290 ) ;
  assign n8292 = n8290 | n8291 ;
  assign n8293 = n8292 ^ x2 ^ 1'b0 ;
  assign n8294 = ( n8258 & n8284 ) | ( n8258 & n8293 ) | ( n8284 & n8293 ) ;
  assign n8295 = ( n7749 & n7924 ) | ( n7749 & n8288 ) | ( n7924 & n8288 ) ;
  assign n8296 = n8288 ^ n7924 ^ n7749 ;
  assign n8297 = ~n6718 & n7829 ;
  assign n8298 = ( ~n6617 & n7833 ) | ( ~n6617 & n8297 ) | ( n7833 & n8297 ) ;
  assign n8299 = n8297 | n8298 ;
  assign n8300 = ( ~n6731 & n7834 ) | ( ~n6731 & n8297 ) | ( n7834 & n8297 ) ;
  assign n8301 = n8299 | n8300 ;
  assign n8302 = ~n6917 & n7838 ;
  assign n8303 = n8301 | n8302 ;
  assign n8304 = n8303 ^ x11 ^ 1'b0 ;
  assign n8305 = n8304 ^ n8295 ^ n7748 ;
  assign n8306 = ( n7748 & n8295 ) | ( n7748 & n8304 ) | ( n8295 & n8304 ) ;
  assign n8307 = ~n6718 & n7932 ;
  assign n8308 = ( ~n6617 & n7943 ) | ( ~n6617 & n8307 ) | ( n7943 & n8307 ) ;
  assign n8309 = n8307 | n8308 ;
  assign n8310 = ( ~n6731 & n7929 ) | ( ~n6731 & n8307 ) | ( n7929 & n8307 ) ;
  assign n8311 = n8309 | n8310 ;
  assign n8312 = ~n6917 & n7930 ;
  assign n8313 = n8311 | n8312 ;
  assign n8314 = n8313 ^ x8 ^ 1'b0 ;
  assign n8315 = ( n7914 & n8281 ) | ( n7914 & n8314 ) | ( n8281 & n8314 ) ;
  assign n8316 = n8314 ^ n8281 ^ n7914 ;
  assign n8317 = ~n6718 & n6791 ;
  assign n8318 = ( ~n6731 & n6788 ) | ( ~n6731 & n8317 ) | ( n6788 & n8317 ) ;
  assign n8319 = ( ~n6617 & n6790 ) | ( ~n6617 & n8317 ) | ( n6790 & n8317 ) ;
  assign n8320 = n8317 | n8318 ;
  assign n8321 = n8319 | n8320 ;
  assign n8322 = n6603 & n8033 ;
  assign n8323 = n6789 & ~n6917 ;
  assign n8324 = ( ~n6731 & n8029 ) | ( ~n6731 & n8322 ) | ( n8029 & n8322 ) ;
  assign n8325 = n8321 | n8323 ;
  assign n8326 = n8322 | n8324 ;
  assign n8327 = ( ~n6718 & n8037 ) | ( ~n6718 & n8322 ) | ( n8037 & n8322 ) ;
  assign n8328 = n8326 | n8327 ;
  assign n8329 = n6724 & n8090 ;
  assign n8330 = ( ~n6602 & n8086 ) | ( ~n6602 & n8329 ) | ( n8086 & n8329 ) ;
  assign n8331 = n8329 | n8330 ;
  assign n8332 = ( ~n6533 & n8088 ) | ( ~n6533 & n8329 ) | ( n8088 & n8329 ) ;
  assign n8333 = n8331 | n8332 ;
  assign n8334 = n7147 & n8034 ;
  assign n8335 = n8328 | n8334 ;
  assign n8336 = n8335 ^ x5 ^ 1'b0 ;
  assign n8337 = n8336 ^ n8285 ^ n8024 ;
  assign n8338 = ( n8024 & n8285 ) | ( n8024 & n8336 ) | ( n8285 & n8336 ) ;
  assign n8339 = ( n7624 & n8089 ) | ( n7624 & n8333 ) | ( n8089 & n8333 ) ;
  assign n8340 = n8333 | n8339 ;
  assign n8341 = n8340 ^ x2 ^ 1'b0 ;
  assign n8342 = ( n8294 & n8337 ) | ( n8294 & n8341 ) | ( n8337 & n8341 ) ;
  assign n8343 = n7147 & n7930 ;
  assign n8344 = n6603 & n7929 ;
  assign n8345 = ( ~n6731 & n7932 ) | ( ~n6731 & n8344 ) | ( n7932 & n8344 ) ;
  assign n8346 = n8344 | n8345 ;
  assign n8347 = ( ~n6718 & n7943 ) | ( ~n6718 & n8344 ) | ( n7943 & n8344 ) ;
  assign n8348 = n8346 | n8347 ;
  assign n8349 = n8343 | n8348 ;
  assign n8350 = n8349 ^ x8 ^ 1'b0 ;
  assign n8351 = ( n7925 & n8315 ) | ( n7925 & n8350 ) | ( n8315 & n8350 ) ;
  assign n8352 = n8350 ^ n8315 ^ n7925 ;
  assign n8353 = n6724 & n6907 ;
  assign n8354 = ( ~n6533 & n6901 ) | ( ~n6533 & n8353 ) | ( n6901 & n8353 ) ;
  assign n8355 = ( ~n6602 & n6906 ) | ( ~n6602 & n8353 ) | ( n6906 & n8353 ) ;
  assign n8356 = n8353 | n8354 ;
  assign n8357 = n6603 & n7834 ;
  assign n8358 = n8355 | n8356 ;
  assign n8359 = ( n6918 & n7624 ) | ( n6918 & n8358 ) | ( n7624 & n8358 ) ;
  assign n8360 = n8358 | n8359 ;
  assign n8361 = ( ~n6731 & n7829 ) | ( ~n6731 & n8357 ) | ( n7829 & n8357 ) ;
  assign n8362 = n8357 | n8361 ;
  assign n8363 = ( ~n6718 & n7833 ) | ( ~n6718 & n8357 ) | ( n7833 & n8357 ) ;
  assign n8364 = n8362 | n8363 ;
  assign n8365 = n7147 & n7838 ;
  assign n8366 = n8364 | n8365 ;
  assign n8367 = n8366 ^ x11 ^ 1'b0 ;
  assign n8368 = n8367 ^ n8306 ^ n7758 ;
  assign n8369 = ( n7758 & n8306 ) | ( n7758 & n8367 ) | ( n8306 & n8367 ) ;
  assign n8370 = ( x2 & x5 ) | ( x2 & ~n6745 ) | ( x5 & ~n6745 ) ;
  assign n8371 = n6745 ^ x5 ^ x2 ;
  assign n8372 = ( n6884 & n8325 ) | ( n6884 & n8371 ) | ( n8325 & n8371 ) ;
  assign n8373 = n8371 ^ n8325 ^ n6884 ;
  assign n8374 = ~n6731 & n6791 ;
  assign n8375 = ( n6603 & n6788 ) | ( n6603 & n8374 ) | ( n6788 & n8374 ) ;
  assign n8376 = n8374 | n8375 ;
  assign n8377 = n8360 ^ x29 ^ 1'b0 ;
  assign n8378 = ( ~n6718 & n6790 ) | ( ~n6718 & n8374 ) | ( n6790 & n8374 ) ;
  assign n8379 = n8376 | n8378 ;
  assign n8380 = n6789 & ~n7147 ;
  assign n8381 = ( n6789 & n8379 ) | ( n6789 & ~n8380 ) | ( n8379 & ~n8380 ) ;
  assign n8382 = n8381 ^ n8370 ^ n6753 ;
  assign n8383 = ( n6753 & ~n8370 ) | ( n6753 & n8381 ) | ( ~n8370 & n8381 ) ;
  assign n8384 = n8382 ^ n8377 ^ n8372 ;
  assign n8385 = ( n8372 & n8377 ) | ( n8372 & ~n8382 ) | ( n8377 & ~n8382 ) ;
  assign n8386 = n6603 & n6907 ;
  assign n8387 = ( ~n6731 & n6901 ) | ( ~n6731 & n8386 ) | ( n6901 & n8386 ) ;
  assign n8388 = n8386 | n8387 ;
  assign n8389 = ( ~n6718 & n6906 ) | ( ~n6718 & n8386 ) | ( n6906 & n8386 ) ;
  assign n8390 = n8388 | n8389 ;
  assign n8391 = ( n6918 & n7147 ) | ( n6918 & n8390 ) | ( n7147 & n8390 ) ;
  assign n8392 = n8390 | n8391 ;
  assign n8393 = ( n6545 & n6753 ) | ( n6545 & n8383 ) | ( n6753 & n8383 ) ;
  assign n8394 = n8383 ^ n6753 ^ n6545 ;
  assign n8395 = n8394 ^ n8385 ^ n7826 ;
  assign n8396 = ( n7826 & n8385 ) | ( n7826 & n8394 ) | ( n8385 & n8394 ) ;
  assign n8397 = n6603 & n8029 ;
  assign n8398 = ( ~n6731 & n8037 ) | ( ~n6731 & n8397 ) | ( n8037 & n8397 ) ;
  assign n8399 = n8397 | n8398 ;
  assign n8400 = ( ~n6602 & n8033 ) | ( ~n6602 & n8397 ) | ( n8033 & n8397 ) ;
  assign n8401 = n8399 | n8400 ;
  assign n8402 = n7125 & n8034 ;
  assign n8403 = n8401 | n8402 ;
  assign n8404 = n8403 ^ x5 ^ 1'b0 ;
  assign n8405 = n8404 ^ n8338 ^ n8283 ;
  assign n8406 = ( n8283 & n8338 ) | ( n8283 & n8404 ) | ( n8338 & n8404 ) ;
  assign n8407 = n6603 & n7932 ;
  assign n8408 = ( ~n6731 & n7943 ) | ( ~n6731 & n8407 ) | ( n7943 & n8407 ) ;
  assign n8409 = n8407 | n8408 ;
  assign n8410 = ( ~n6602 & n7929 ) | ( ~n6602 & n8407 ) | ( n7929 & n8407 ) ;
  assign n8411 = n8409 | n8410 ;
  assign n8412 = n7125 & n7930 ;
  assign n8413 = n8411 | n8412 ;
  assign n8414 = n8413 ^ x8 ^ 1'b0 ;
  assign n8415 = ( n8296 & n8351 ) | ( n8296 & n8414 ) | ( n8351 & n8414 ) ;
  assign n8416 = n8414 ^ n8351 ^ n8296 ;
  assign n8417 = n6603 & n6901 ;
  assign n8418 = ( ~n6731 & n6906 ) | ( ~n6731 & n8417 ) | ( n6906 & n8417 ) ;
  assign n8419 = n8417 | n8418 ;
  assign n8420 = ( ~n6602 & n6907 ) | ( ~n6602 & n8417 ) | ( n6907 & n8417 ) ;
  assign n8421 = n8419 | n8420 ;
  assign n8422 = n6603 & n7829 ;
  assign n8423 = ( ~n6731 & n7833 ) | ( ~n6731 & n8422 ) | ( n7833 & n8422 ) ;
  assign n8424 = n8422 | n8423 ;
  assign n8425 = ( ~n6602 & n7834 ) | ( ~n6602 & n8422 ) | ( n7834 & n8422 ) ;
  assign n8426 = n8424 | n8425 ;
  assign n8427 = n7125 & n7838 ;
  assign n8428 = ( n6918 & n7125 ) | ( n6918 & n8421 ) | ( n7125 & n8421 ) ;
  assign n8429 = n8421 | n8428 ;
  assign n8430 = n8426 | n8427 ;
  assign n8431 = n8430 ^ x11 ^ 1'b0 ;
  assign n8432 = n8431 ^ n8369 ^ n7768 ;
  assign n8433 = ( n7768 & n8369 ) | ( n7768 & n8431 ) | ( n8369 & n8431 ) ;
  assign n8434 = n6603 & n7833 ;
  assign n8435 = ( ~n6602 & n7829 ) | ( ~n6602 & n8434 ) | ( n7829 & n8434 ) ;
  assign n8436 = n8434 | n8435 ;
  assign n8437 = ( ~n6533 & n7834 ) | ( ~n6533 & n8434 ) | ( n7834 & n8434 ) ;
  assign n8438 = n8436 | n8437 ;
  assign n8439 = ( ~n7135 & n7838 ) | ( ~n7135 & n8438 ) | ( n7838 & n8438 ) ;
  assign n8440 = n8438 | n8439 ;
  assign n8441 = n8440 ^ x11 ^ 1'b0 ;
  assign n8442 = ( n7779 & n8433 ) | ( n7779 & n8441 ) | ( n8433 & n8441 ) ;
  assign n8443 = n8441 ^ n8433 ^ n7779 ;
  assign n8444 = n6603 & n6906 ;
  assign n8445 = ( ~n6602 & n6901 ) | ( ~n6602 & n8444 ) | ( n6901 & n8444 ) ;
  assign n8446 = n8444 | n8445 ;
  assign n8447 = ( ~n6533 & n6907 ) | ( ~n6533 & n8444 ) | ( n6907 & n8444 ) ;
  assign n8448 = n8446 | n8447 ;
  assign n8449 = n6918 & ~n7135 ;
  assign n8450 = n8448 | n8449 ;
  assign n8451 = n8450 ^ x29 ^ 1'b0 ;
  assign n8452 = ( n6926 & n8373 ) | ( n6926 & n8451 ) | ( n8373 & n8451 ) ;
  assign n8453 = n8451 ^ n8373 ^ n6926 ;
  assign n8454 = n6603 & n7943 ;
  assign n8455 = ( ~n6602 & n7932 ) | ( ~n6602 & n8454 ) | ( n7932 & n8454 ) ;
  assign n8456 = n8454 | n8455 ;
  assign n8457 = ( ~n6533 & n7929 ) | ( ~n6533 & n8454 ) | ( n7929 & n8454 ) ;
  assign n8458 = n8456 | n8457 ;
  assign n8459 = ( ~n7135 & n7930 ) | ( ~n7135 & n8458 ) | ( n7930 & n8458 ) ;
  assign n8460 = n8458 | n8459 ;
  assign n8461 = n8460 ^ x8 ^ 1'b0 ;
  assign n8462 = ( n8305 & n8415 ) | ( n8305 & n8461 ) | ( n8415 & n8461 ) ;
  assign n8463 = n8461 ^ n8415 ^ n8305 ;
  assign n8464 = ~n6602 & n6791 ;
  assign n8465 = ( n6603 & n6790 ) | ( n6603 & n8464 ) | ( n6790 & n8464 ) ;
  assign n8466 = n8464 | n8465 ;
  assign n8467 = ( ~n6533 & n6788 ) | ( ~n6533 & n8464 ) | ( n6788 & n8464 ) ;
  assign n8468 = n8466 | n8467 ;
  assign n8469 = n6789 & ~n7135 ;
  assign n8470 = n8468 | n8469 ;
  assign n8471 = ( x8 & ~n6623 ) | ( x8 & n6753 ) | ( ~n6623 & n6753 ) ;
  assign n8472 = n6753 ^ n6623 ^ x8 ;
  assign n8473 = ( n8393 & n8470 ) | ( n8393 & n8472 ) | ( n8470 & n8472 ) ;
  assign n8474 = n8472 ^ n8470 ^ n8393 ;
  assign n8475 = n6603 & n8037 ;
  assign n8476 = ( ~n6602 & n8029 ) | ( ~n6602 & n8475 ) | ( n8029 & n8475 ) ;
  assign n8477 = n8475 | n8476 ;
  assign n8478 = ( ~n6533 & n8033 ) | ( ~n6533 & n8475 ) | ( n8033 & n8475 ) ;
  assign n8479 = n8477 | n8478 ;
  assign n8480 = ( ~n7135 & n8034 ) | ( ~n7135 & n8479 ) | ( n8034 & n8479 ) ;
  assign n8481 = n8479 | n8480 ;
  assign n8482 = n8481 ^ x5 ^ 1'b0 ;
  assign n8483 = ( n8316 & n8406 ) | ( n8316 & n8482 ) | ( n8406 & n8482 ) ;
  assign n8484 = n8482 ^ n8406 ^ n8316 ;
  assign n8485 = n6724 & n7037 ;
  assign n8486 = ( ~n6533 & n7036 ) | ( ~n6533 & n8485 ) | ( n7036 & n8485 ) ;
  assign n8487 = n8485 | n8486 ;
  assign n8488 = ( ~n6602 & n7052 ) | ( ~n6602 & n8485 ) | ( n7052 & n8485 ) ;
  assign n8489 = n8487 | n8488 ;
  assign n8490 = n7035 & n7624 ;
  assign n8491 = n8489 | n8490 ;
  assign n8492 = n8491 ^ x26 ^ 1'b0 ;
  assign n8493 = n8392 ^ x29 ^ 1'b0 ;
  assign n8494 = ( n6924 & n8492 ) | ( n6924 & n8493 ) | ( n8492 & n8493 ) ;
  assign n8495 = n8493 ^ n8492 ^ n6924 ;
  assign n8496 = n6724 & n7929 ;
  assign n8497 = ( ~n6533 & n7932 ) | ( ~n6533 & n8496 ) | ( n7932 & n8496 ) ;
  assign n8498 = n8496 | n8497 ;
  assign n8499 = ( ~n6602 & n7943 ) | ( ~n6602 & n8496 ) | ( n7943 & n8496 ) ;
  assign n8500 = n8498 | n8499 ;
  assign n8501 = ( n7624 & n7930 ) | ( n7624 & n8500 ) | ( n7930 & n8500 ) ;
  assign n8502 = n8500 | n8501 ;
  assign n8503 = n8502 ^ x8 ^ 1'b0 ;
  assign n8504 = n8503 ^ n8462 ^ n8368 ;
  assign n8505 = ( n8368 & n8462 ) | ( n8368 & n8503 ) | ( n8462 & n8503 ) ;
  assign n8506 = n6724 & n8033 ;
  assign n8507 = ( ~n6533 & n8029 ) | ( ~n6533 & n8506 ) | ( n8029 & n8506 ) ;
  assign n8508 = n8506 | n8507 ;
  assign n8509 = ( ~n6602 & n8037 ) | ( ~n6602 & n8506 ) | ( n8037 & n8506 ) ;
  assign n8510 = n8508 | n8509 ;
  assign n8511 = ( n7624 & n8034 ) | ( n7624 & n8510 ) | ( n8034 & n8510 ) ;
  assign n8512 = n8510 | n8511 ;
  assign n8513 = n8512 ^ x5 ^ 1'b0 ;
  assign n8514 = ( n8352 & n8483 ) | ( n8352 & n8513 ) | ( n8483 & n8513 ) ;
  assign n8515 = n8513 ^ n8483 ^ n8352 ;
  assign n8516 = n6724 & n7834 ;
  assign n8517 = ( ~n6533 & n7829 ) | ( ~n6533 & n8516 ) | ( n7829 & n8516 ) ;
  assign n8518 = n8516 | n8517 ;
  assign n8519 = ( ~n6602 & n7833 ) | ( ~n6602 & n8516 ) | ( n7833 & n8516 ) ;
  assign n8520 = n8518 | n8519 ;
  assign n8521 = ( n7624 & n7838 ) | ( n7624 & n8520 ) | ( n7838 & n8520 ) ;
  assign n8522 = n6789 & ~n7624 ;
  assign n8523 = n8520 | n8521 ;
  assign n8524 = n8523 ^ x11 ^ 1'b0 ;
  assign n8525 = n8524 ^ n8442 ^ n7789 ;
  assign n8526 = ( n7789 & n8442 ) | ( n7789 & n8524 ) | ( n8442 & n8524 ) ;
  assign n8527 = ~n6533 & n6791 ;
  assign n8528 = ( n6724 & n6788 ) | ( n6724 & n8527 ) | ( n6788 & n8527 ) ;
  assign n8529 = ( ~n6602 & n6790 ) | ( ~n6602 & n8527 ) | ( n6790 & n8527 ) ;
  assign n8530 = n8527 | n8528 ;
  assign n8531 = n8529 | n8530 ;
  assign n8532 = ( n6789 & ~n8522 ) | ( n6789 & n8531 ) | ( ~n8522 & n8531 ) ;
  assign n8533 = ( n6721 & n8471 ) | ( n6721 & ~n8532 ) | ( n8471 & ~n8532 ) ;
  assign n8534 = ( ~n6627 & n6721 ) | ( ~n6627 & n8533 ) | ( n6721 & n8533 ) ;
  assign n8535 = n8532 ^ n8471 ^ n6721 ;
  assign n8536 = n8533 ^ n6721 ^ n6627 ;
  assign n8537 = n6600 & n8090 ;
  assign n8538 = ( n6724 & n8088 ) | ( n6724 & n8537 ) | ( n8088 & n8537 ) ;
  assign n8539 = n8537 | n8538 ;
  assign n8540 = ( n6600 & n6724 ) | ( n6600 & ~n7653 ) | ( n6724 & ~n7653 ) ;
  assign n8541 = ( ~n6533 & n8086 ) | ( ~n6533 & n8537 ) | ( n8086 & n8537 ) ;
  assign n8542 = n7653 ^ n6724 ^ n6600 ;
  assign n8543 = n8539 | n8541 ;
  assign n8544 = ( n8089 & ~n8542 ) | ( n8089 & n8543 ) | ( ~n8542 & n8543 ) ;
  assign n8545 = n8543 | n8544 ;
  assign n8546 = n8540 ^ n6600 ^ n6170 ;
  assign n8547 = n8545 ^ x2 ^ 1'b0 ;
  assign n8548 = ( n8342 & n8405 ) | ( n8342 & n8547 ) | ( n8405 & n8547 ) ;
  assign n8549 = n6600 & n8088 ;
  assign n8550 = ( n6724 & n8086 ) | ( n6724 & n8549 ) | ( n8086 & n8549 ) ;
  assign n8551 = n8549 | n8550 ;
  assign n8552 = ( ~n6170 & n8090 ) | ( ~n6170 & n8549 ) | ( n8090 & n8549 ) ;
  assign n8553 = n8551 | n8552 ;
  assign n8554 = n8089 & ~n8546 ;
  assign n8555 = n8553 | n8554 ;
  assign n8556 = ( ~x11 & n6721 ) | ( ~x11 & n6754 ) | ( n6721 & n6754 ) ;
  assign n8557 = n6754 ^ n6721 ^ x11 ;
  assign n8558 = n6789 & ~n8546 ;
  assign n8559 = n8555 ^ x2 ^ 1'b0 ;
  assign n8560 = ( n8484 & n8548 ) | ( n8484 & n8559 ) | ( n8548 & n8559 ) ;
  assign n8561 = ( n6600 & n6791 ) | ( n6600 & n8558 ) | ( n6791 & n8558 ) ;
  assign n8562 = n8558 | n8561 ;
  assign n8563 = n6170 & n6788 ;
  assign n8564 = ( n6724 & n6790 ) | ( n6724 & n8558 ) | ( n6790 & n8558 ) ;
  assign n8565 = n8562 | n8564 ;
  assign n8566 = ( n6788 & ~n8563 ) | ( n6788 & n8565 ) | ( ~n8563 & n8565 ) ;
  assign n8567 = n8566 ^ n8557 ^ n8534 ;
  assign n8568 = ( n8534 & n8557 ) | ( n8534 & ~n8566 ) | ( n8557 & ~n8566 ) ;
  assign n8569 = n6600 & n8033 ;
  assign n8570 = ( n6724 & n8029 ) | ( n6724 & n8569 ) | ( n8029 & n8569 ) ;
  assign n8571 = n8569 | n8570 ;
  assign n8572 = ( ~n6533 & n8037 ) | ( ~n6533 & n8569 ) | ( n8037 & n8569 ) ;
  assign n8573 = n8571 | n8572 ;
  assign n8574 = ( n8034 & ~n8542 ) | ( n8034 & n8573 ) | ( ~n8542 & n8573 ) ;
  assign n8575 = n8573 | n8574 ;
  assign n8576 = n8575 ^ x5 ^ 1'b0 ;
  assign n8577 = ( n8416 & n8514 ) | ( n8416 & n8576 ) | ( n8514 & n8576 ) ;
  assign n8578 = n8576 ^ n8514 ^ n8416 ;
  assign n8579 = n6600 & n8029 ;
  assign n8580 = ( n6724 & n8037 ) | ( n6724 & n8579 ) | ( n8037 & n8579 ) ;
  assign n8581 = n8579 | n8580 ;
  assign n8582 = ( ~n6170 & n8033 ) | ( ~n6170 & n8579 ) | ( n8033 & n8579 ) ;
  assign n8583 = n8581 | n8582 ;
  assign n8584 = n8034 & ~n8546 ;
  assign n8585 = n8583 | n8584 ;
  assign n8586 = n8585 ^ x5 ^ 1'b0 ;
  assign n8587 = n6529 & n8090 ;
  assign n8588 = ( n8463 & n8577 ) | ( n8463 & n8586 ) | ( n8577 & n8586 ) ;
  assign n8589 = n8586 ^ n8577 ^ n8463 ;
  assign n8590 = ( ~n6170 & n6600 ) | ( ~n6170 & n8540 ) | ( n6600 & n8540 ) ;
  assign n8591 = ( n6600 & n8086 ) | ( n6600 & n8587 ) | ( n8086 & n8587 ) ;
  assign n8592 = n8587 | n8591 ;
  assign n8593 = n8590 ^ n6529 ^ n6170 ;
  assign n8594 = ( ~n6170 & n8088 ) | ( ~n6170 & n8587 ) | ( n8088 & n8587 ) ;
  assign n8595 = n8592 | n8594 ;
  assign n8596 = n8089 & ~n8593 ;
  assign n8597 = n8595 | n8596 ;
  assign n8598 = n8597 ^ x2 ^ 1'b0 ;
  assign n8599 = n8034 & ~n8593 ;
  assign n8600 = ( n8515 & n8560 ) | ( n8515 & n8598 ) | ( n8560 & n8598 ) ;
  assign n8601 = n6529 & n8033 ;
  assign n8602 = ( n6600 & n8037 ) | ( n6600 & n8601 ) | ( n8037 & n8601 ) ;
  assign n8603 = n8601 | n8602 ;
  assign n8604 = ( ~n6170 & n8029 ) | ( ~n6170 & n8601 ) | ( n8029 & n8601 ) ;
  assign n8605 = n8603 | n8604 ;
  assign n8606 = n8599 | n8605 ;
  assign n8607 = n8606 ^ x5 ^ 1'b0 ;
  assign n8608 = ( n8504 & n8588 ) | ( n8504 & n8607 ) | ( n8588 & n8607 ) ;
  assign n8609 = n8607 ^ n8588 ^ n8504 ;
  assign n8610 = n6600 & n7486 ;
  assign n8611 = ( n6724 & n7485 ) | ( n6724 & n8610 ) | ( n7485 & n8610 ) ;
  assign n8612 = n8610 | n8611 ;
  assign n8613 = ( ~n6533 & n7493 ) | ( ~n6533 & n8610 ) | ( n7493 & n8610 ) ;
  assign n8614 = n8612 | n8613 ;
  assign n8615 = n6600 & n7192 ;
  assign n8616 = ( n6724 & n7190 ) | ( n6724 & n8615 ) | ( n7190 & n8615 ) ;
  assign n8617 = n8615 | n8616 ;
  assign n8618 = ( ~n6170 & n7188 ) | ( ~n6170 & n8615 ) | ( n7188 & n8615 ) ;
  assign n8619 = n8617 | n8618 ;
  assign n8620 = n6600 & n7667 ;
  assign n8621 = n6600 & n7929 ;
  assign n8622 = ( n6724 & n7932 ) | ( n6724 & n8621 ) | ( n7932 & n8621 ) ;
  assign n8623 = ( ~n6533 & n7943 ) | ( ~n6533 & n8621 ) | ( n7943 & n8621 ) ;
  assign n8624 = n8621 | n8622 ;
  assign n8625 = n8623 | n8624 ;
  assign n8626 = ( n7930 & ~n8542 ) | ( n7930 & n8625 ) | ( ~n8542 & n8625 ) ;
  assign n8627 = n8625 | n8626 ;
  assign n8628 = n8627 ^ x8 ^ 1'b0 ;
  assign n8629 = ( n8432 & n8505 ) | ( n8432 & n8628 ) | ( n8505 & n8628 ) ;
  assign n8630 = n8628 ^ n8505 ^ n8432 ;
  assign n8631 = n6600 & n7188 ;
  assign n8632 = ( ~n6533 & n7190 ) | ( ~n6533 & n8631 ) | ( n7190 & n8631 ) ;
  assign n8633 = n7487 & ~n8542 ;
  assign n8634 = n8614 | n8633 ;
  assign n8635 = ( n6724 & n7192 ) | ( n6724 & n8631 ) | ( n7192 & n8631 ) ;
  assign n8636 = n8631 | n8635 ;
  assign n8637 = n8632 | n8636 ;
  assign n8638 = n8634 ^ x17 ^ 1'b0 ;
  assign n8639 = ( n7469 & n7660 ) | ( n7469 & n8638 ) | ( n7660 & n8638 ) ;
  assign n8640 = n8638 ^ n7660 ^ n7469 ;
  assign n8641 = n6600 & n7337 ;
  assign n8642 = n7340 & ~n8542 ;
  assign n8643 = ( n6724 & n7339 ) | ( n6724 & n8641 ) | ( n7339 & n8641 ) ;
  assign n8644 = n8641 | n8643 ;
  assign n8645 = ( ~n6533 & n7338 ) | ( ~n6533 & n8641 ) | ( n7338 & n8641 ) ;
  assign n8646 = n8644 | n8645 ;
  assign n8647 = n7196 & ~n8542 ;
  assign n8648 = n8637 | n8647 ;
  assign n8649 = n7196 & ~n8546 ;
  assign n8650 = n8619 | n8649 ;
  assign n8651 = ~n8642 & n8646 ;
  assign n8652 = n8650 ^ x23 ^ 1'b0 ;
  assign n8653 = n8652 ^ n7184 ^ n7142 ;
  assign n8654 = ( n7142 & n7184 ) | ( n7142 & n8652 ) | ( n7184 & n8652 ) ;
  assign n8655 = n6600 & n6901 ;
  assign n8656 = ( n6724 & n6906 ) | ( n6724 & n8655 ) | ( n6906 & n8655 ) ;
  assign n8657 = n8655 | n8656 ;
  assign n8658 = ( ~n6170 & n6907 ) | ( ~n6170 & n8655 ) | ( n6907 & n8655 ) ;
  assign n8659 = n8657 | n8658 ;
  assign n8660 = n6918 & ~n8546 ;
  assign n8661 = n8659 | n8660 ;
  assign n8662 = n8661 ^ x29 ^ 1'b0 ;
  assign n8663 = n8648 ^ x23 ^ 1'b0 ;
  assign n8664 = n8663 ^ n7629 ^ n7183 ;
  assign n8665 = ( n7183 & n7629 ) | ( n7183 & n8663 ) | ( n7629 & n8663 ) ;
  assign n8666 = ( n8396 & n8474 ) | ( n8396 & n8662 ) | ( n8474 & n8662 ) ;
  assign n8667 = n8651 ^ n8642 ^ x20 ;
  assign n8668 = ( n6724 & n7669 ) | ( n6724 & n8620 ) | ( n7669 & n8620 ) ;
  assign n8669 = ( ~n6533 & n7674 ) | ( ~n6533 & n8620 ) | ( n7674 & n8620 ) ;
  assign n8670 = n8620 | n8668 ;
  assign n8671 = n8669 | n8670 ;
  assign n8672 = ( n7666 & ~n8542 ) | ( n7666 & n8671 ) | ( ~n8542 & n8671 ) ;
  assign n8673 = n8671 | n8672 ;
  assign n8674 = n8667 ^ n7649 ^ n7327 ;
  assign n8675 = n8673 ^ x14 ^ 1'b0 ;
  assign n8676 = n8675 ^ n7818 ^ n7618 ;
  assign n8677 = ( n7618 & n7818 ) | ( n7618 & n8675 ) | ( n7818 & n8675 ) ;
  assign n8678 = n7930 & ~n8546 ;
  assign n8679 = ( n7327 & n7649 ) | ( n7327 & n8667 ) | ( n7649 & n8667 ) ;
  assign n8680 = n6600 & n7932 ;
  assign n8681 = ( ~n6170 & n7929 ) | ( ~n6170 & n8680 ) | ( n7929 & n8680 ) ;
  assign n8682 = n8662 ^ n8474 ^ n8396 ;
  assign n8683 = ( n6724 & n7943 ) | ( n6724 & n8680 ) | ( n7943 & n8680 ) ;
  assign n8684 = n8680 | n8683 ;
  assign n8685 = n8681 | n8684 ;
  assign n8686 = n8678 | n8685 ;
  assign n8687 = n8686 ^ x8 ^ 1'b0 ;
  assign n8688 = ( n8443 & n8629 ) | ( n8443 & n8687 ) | ( n8629 & n8687 ) ;
  assign n8689 = n8687 ^ n8629 ^ n8443 ;
  assign n8690 = n6600 & n7834 ;
  assign n8691 = ( n6724 & n7829 ) | ( n6724 & n8690 ) | ( n7829 & n8690 ) ;
  assign n8692 = n8690 | n8691 ;
  assign n8693 = ( ~n6533 & n7833 ) | ( ~n6533 & n8690 ) | ( n7833 & n8690 ) ;
  assign n8694 = n8692 | n8693 ;
  assign n8695 = ( n7838 & ~n8542 ) | ( n7838 & n8694 ) | ( ~n8542 & n8694 ) ;
  assign n8696 = n8694 | n8695 ;
  assign n8697 = n8696 ^ x11 ^ 1'b0 ;
  assign n8698 = ( n7798 & n8526 ) | ( n7798 & n8697 ) | ( n8526 & n8697 ) ;
  assign n8699 = n8697 ^ n8526 ^ n7798 ;
  assign n8700 = n6600 & n7339 ;
  assign n8701 = ( n6724 & n7338 ) | ( n6724 & n8700 ) | ( n7338 & n8700 ) ;
  assign n8702 = n8700 | n8701 ;
  assign n8703 = ( ~n6170 & n7337 ) | ( ~n6170 & n8700 ) | ( n7337 & n8700 ) ;
  assign n8704 = n8702 | n8703 ;
  assign n8705 = n7340 & ~n8546 ;
  assign n8706 = n8704 & ~n8705 ;
  assign n8707 = n8706 ^ n8705 ^ x20 ;
  assign n8708 = ( ~n7331 & n8679 ) | ( ~n7331 & n8707 ) | ( n8679 & n8707 ) ;
  assign n8709 = n8707 ^ n8679 ^ n7331 ;
  assign n8710 = n6600 & n7485 ;
  assign n8711 = ( n6724 & n7493 ) | ( n6724 & n8710 ) | ( n7493 & n8710 ) ;
  assign n8712 = n8710 | n8711 ;
  assign n8713 = ( ~n6170 & n7486 ) | ( ~n6170 & n8710 ) | ( n7486 & n8710 ) ;
  assign n8714 = n8712 | n8713 ;
  assign n8715 = n7487 & ~n8546 ;
  assign n8716 = n8714 | n8715 ;
  assign n8717 = n8716 ^ x17 ^ 1'b0 ;
  assign n8718 = ( ~n7480 & n8639 ) | ( ~n7480 & n8717 ) | ( n8639 & n8717 ) ;
  assign n8719 = n8717 ^ n8639 ^ n7480 ;
  assign n8720 = n6600 & n7669 ;
  assign n8721 = ( n6724 & n7674 ) | ( n6724 & n8720 ) | ( n7674 & n8720 ) ;
  assign n8722 = n8720 | n8721 ;
  assign n8723 = ( ~n6170 & n7667 ) | ( ~n6170 & n8720 ) | ( n7667 & n8720 ) ;
  assign n8724 = n8722 | n8723 ;
  assign n8725 = n7666 & ~n8546 ;
  assign n8726 = n8724 | n8725 ;
  assign n8727 = n8726 ^ x14 ^ 1'b0 ;
  assign n8728 = ( n7639 & n8677 ) | ( n7639 & n8727 ) | ( n8677 & n8727 ) ;
  assign n8729 = n8727 ^ n8677 ^ n7639 ;
  assign n8730 = n6600 & n7829 ;
  assign n8731 = ( n6724 & n7833 ) | ( n6724 & n8730 ) | ( n7833 & n8730 ) ;
  assign n8732 = n8730 | n8731 ;
  assign n8733 = ( ~n6170 & n7834 ) | ( ~n6170 & n8730 ) | ( n7834 & n8730 ) ;
  assign n8734 = n8732 | n8733 ;
  assign n8735 = n7838 & ~n8546 ;
  assign n8736 = n8734 | n8735 ;
  assign n8737 = n8736 ^ x11 ^ 1'b0 ;
  assign n8738 = n8737 ^ n8698 ^ n7808 ;
  assign n8739 = ( n7808 & n8698 ) | ( n7808 & n8737 ) | ( n8698 & n8737 ) ;
  assign n8740 = n6600 & n7037 ;
  assign n8741 = ( n6724 & n7036 ) | ( n6724 & n8740 ) | ( n7036 & n8740 ) ;
  assign n8742 = n8740 | n8741 ;
  assign n8743 = ( ~n6533 & n7052 ) | ( ~n6533 & n8740 ) | ( n7052 & n8740 ) ;
  assign n8744 = n8742 | n8743 ;
  assign n8745 = n7035 & ~n8542 ;
  assign n8746 = n8429 ^ x29 ^ 1'b0 ;
  assign n8747 = n8744 | n8745 ;
  assign n8748 = n8747 ^ x26 ^ 1'b0 ;
  assign n8749 = n8748 ^ n8746 ^ n6925 ;
  assign n8750 = ( ~n6925 & n8746 ) | ( ~n6925 & n8748 ) | ( n8746 & n8748 ) ;
  assign n8751 = n6600 & n6907 ;
  assign n8752 = n7035 & ~n8546 ;
  assign n8753 = ( n6724 & n6901 ) | ( n6724 & n8751 ) | ( n6901 & n8751 ) ;
  assign n8754 = n8751 | n8753 ;
  assign n8755 = ( ~n6533 & n6906 ) | ( ~n6533 & n8751 ) | ( n6906 & n8751 ) ;
  assign n8756 = n8754 | n8755 ;
  assign n8757 = n6789 & ~n8542 ;
  assign n8758 = n6918 & ~n8542 ;
  assign n8759 = n8756 & ~n8758 ;
  assign n8760 = n8759 ^ n8758 ^ x29 ;
  assign n8761 = ( n6724 & n6791 ) | ( n6724 & n8757 ) | ( n6791 & n8757 ) ;
  assign n8762 = n8757 | n8761 ;
  assign n8763 = ( ~n6533 & n6790 ) | ( ~n6533 & n8757 ) | ( n6790 & n8757 ) ;
  assign n8764 = n6600 & n7036 ;
  assign n8765 = ( n6724 & n7052 ) | ( n6724 & n8764 ) | ( n7052 & n8764 ) ;
  assign n8766 = n8764 | n8765 ;
  assign n8767 = ( ~n6170 & n7037 ) | ( ~n6170 & n8764 ) | ( n7037 & n8764 ) ;
  assign n8768 = n8766 | n8767 ;
  assign n8769 = n8762 | n8763 ;
  assign n8770 = ~n8752 & n8768 ;
  assign n8771 = n8770 ^ n8752 ^ x26 ;
  assign n8772 = n8771 ^ n8750 ^ n8453 ;
  assign n8773 = ( n8453 & n8750 ) | ( n8453 & n8771 ) | ( n8750 & n8771 ) ;
  assign n8774 = n6529 & n7188 ;
  assign n8775 = ( n6600 & n7190 ) | ( n6600 & n8774 ) | ( n7190 & n8774 ) ;
  assign n8776 = n8774 | n8775 ;
  assign n8777 = ( ~n6170 & n7192 ) | ( ~n6170 & n8774 ) | ( n7192 & n8774 ) ;
  assign n8778 = n8776 | n8777 ;
  assign n8779 = n7196 & ~n8593 ;
  assign n8780 = ( ~n6170 & n6529 ) | ( ~n6170 & n8590 ) | ( n6529 & n8590 ) ;
  assign n8781 = n8778 | n8779 ;
  assign n8782 = n8781 ^ x23 ^ 1'b0 ;
  assign n8783 = n8782 ^ n8495 ^ n7141 ;
  assign n8784 = ( n7141 & n8495 ) | ( n7141 & n8782 ) | ( n8495 & n8782 ) ;
  assign n8785 = n6529 & n7667 ;
  assign n8786 = ( n6600 & n7674 ) | ( n6600 & n8785 ) | ( n7674 & n8785 ) ;
  assign n8787 = n8785 | n8786 ;
  assign n8788 = ( ~n6170 & n7669 ) | ( ~n6170 & n8785 ) | ( n7669 & n8785 ) ;
  assign n8789 = n8787 | n8788 ;
  assign n8790 = n7666 & ~n8593 ;
  assign n8791 = n8789 | n8790 ;
  assign n8792 = n8791 ^ x14 ^ 1'b0 ;
  assign n8793 = ( n7659 & n8728 ) | ( n7659 & n8792 ) | ( n8728 & n8792 ) ;
  assign n8794 = n8792 ^ n8728 ^ n7659 ;
  assign n8795 = n6529 & n7486 ;
  assign n8796 = ( n6600 & n7493 ) | ( n6600 & n8795 ) | ( n7493 & n8795 ) ;
  assign n8797 = n8795 | n8796 ;
  assign n8798 = ( ~n6170 & n7485 ) | ( ~n6170 & n8795 ) | ( n7485 & n8795 ) ;
  assign n8799 = n8797 | n8798 ;
  assign n8800 = n7487 & ~n8593 ;
  assign n8801 = n8799 | n8800 ;
  assign n8802 = n8801 ^ x17 ^ 1'b0 ;
  assign n8803 = ( ~n7648 & n8718 ) | ( ~n7648 & n8802 ) | ( n8718 & n8802 ) ;
  assign n8804 = n8802 ^ n8718 ^ n7648 ;
  assign n8805 = n6529 & n7037 ;
  assign n8806 = ( n6600 & n7052 ) | ( n6600 & n8805 ) | ( n7052 & n8805 ) ;
  assign n8807 = n8805 | n8806 ;
  assign n8808 = ( ~n6170 & n7036 ) | ( ~n6170 & n8805 ) | ( n7036 & n8805 ) ;
  assign n8809 = n8807 | n8808 ;
  assign n8810 = n7035 & ~n8593 ;
  assign n8811 = n8809 | n8810 ;
  assign n8812 = n8811 ^ x26 ^ 1'b0 ;
  assign n8813 = n8812 ^ n8452 ^ n8384 ;
  assign n8814 = ( ~n8384 & n8452 ) | ( ~n8384 & n8812 ) | ( n8452 & n8812 ) ;
  assign n8815 = n6529 & n7337 ;
  assign n8816 = ( n6600 & n7338 ) | ( n6600 & n8815 ) | ( n7338 & n8815 ) ;
  assign n8817 = n8815 | n8816 ;
  assign n8818 = ( ~n6170 & n7339 ) | ( ~n6170 & n8815 ) | ( n7339 & n8815 ) ;
  assign n8819 = n8817 | n8818 ;
  assign n8820 = n7340 & ~n8593 ;
  assign n8821 = n8819 & ~n8820 ;
  assign n8822 = n8821 ^ n8820 ^ x20 ;
  assign n8823 = n8822 ^ n8708 ^ n7628 ;
  assign n8824 = ( n7628 & n8708 ) | ( n7628 & n8822 ) | ( n8708 & n8822 ) ;
  assign n8825 = n6529 & n6907 ;
  assign n8826 = ( n6600 & n6906 ) | ( n6600 & n8825 ) | ( n6906 & n8825 ) ;
  assign n8827 = n8825 | n8826 ;
  assign n8828 = ( ~n6170 & n6901 ) | ( ~n6170 & n8825 ) | ( n6901 & n8825 ) ;
  assign n8829 = n8827 | n8828 ;
  assign n8830 = n6600 & ~n6788 ;
  assign n8831 = ( n6600 & n8769 ) | ( n6600 & ~n8830 ) | ( n8769 & ~n8830 ) ;
  assign n8832 = n6918 & ~n8593 ;
  assign n8833 = n8829 & ~n8832 ;
  assign n8834 = n8833 ^ n8832 ^ x29 ;
  assign n8835 = ( n8473 & n8535 ) | ( n8473 & n8834 ) | ( n8535 & n8834 ) ;
  assign n8836 = n8834 ^ n8535 ^ n8473 ;
  assign n8837 = n6529 & n7834 ;
  assign n8838 = ( n6600 & n7833 ) | ( n6600 & n8837 ) | ( n7833 & n8837 ) ;
  assign n8839 = n8837 | n8838 ;
  assign n8840 = ( ~n6170 & n7829 ) | ( ~n6170 & n8837 ) | ( n7829 & n8837 ) ;
  assign n8841 = n8839 | n8840 ;
  assign n8842 = n7838 & ~n8593 ;
  assign n8843 = n8841 | n8842 ;
  assign n8844 = n8843 ^ x11 ^ 1'b0 ;
  assign n8845 = n8844 ^ n8739 ^ n7819 ;
  assign n8846 = ( n7819 & n8739 ) | ( n7819 & n8844 ) | ( n8739 & n8844 ) ;
  assign n8847 = n6529 & n7929 ;
  assign n8848 = ( n6600 & n7943 ) | ( n6600 & n8847 ) | ( n7943 & n8847 ) ;
  assign n8849 = n8847 | n8848 ;
  assign n8850 = ( ~n6170 & n7932 ) | ( ~n6170 & n8847 ) | ( n7932 & n8847 ) ;
  assign n8851 = n8849 | n8850 ;
  assign n8852 = n7930 & ~n8593 ;
  assign n8853 = n8851 | n8852 ;
  assign n8854 = n8853 ^ x8 ^ 1'b0 ;
  assign n8855 = n6789 & ~n8593 ;
  assign n8856 = n8854 ^ n8688 ^ n8525 ;
  assign n8857 = ( n8525 & n8688 ) | ( n8525 & n8854 ) | ( n8688 & n8854 ) ;
  assign n8858 = ~n6170 & n6791 ;
  assign n8859 = ( n6529 & n6788 ) | ( n6529 & n8858 ) | ( n6788 & n8858 ) ;
  assign n8860 = n8858 | n8859 ;
  assign n8861 = ( n6600 & n6790 ) | ( n6600 & n8858 ) | ( n6790 & n8858 ) ;
  assign n8862 = n8860 | n8861 ;
  assign n8863 = n8855 | n8862 ;
  assign n8864 = n6529 & n8088 ;
  assign n8865 = n8780 ^ n6729 ^ n6529 ;
  assign n8866 = ( ~n6170 & n8086 ) | ( ~n6170 & n8864 ) | ( n8086 & n8864 ) ;
  assign n8867 = n8864 | n8866 ;
  assign n8868 = ( ~n6729 & n8090 ) | ( ~n6729 & n8864 ) | ( n8090 & n8864 ) ;
  assign n8869 = n8867 | n8868 ;
  assign n8870 = n8089 & ~n8865 ;
  assign n8871 = n8869 | n8870 ;
  assign n8872 = n8871 ^ x2 ^ 1'b0 ;
  assign n8873 = ( n8578 & n8600 ) | ( n8578 & n8872 ) | ( n8600 & n8872 ) ;
  assign n8874 = n6204 & n8090 ;
  assign n8875 = ( n6529 & ~n6729 ) | ( n6529 & n8780 ) | ( ~n6729 & n8780 ) ;
  assign n8876 = ( ~n6729 & n8088 ) | ( ~n6729 & n8874 ) | ( n8088 & n8874 ) ;
  assign n8877 = ( n6529 & n8086 ) | ( n6529 & n8874 ) | ( n8086 & n8874 ) ;
  assign n8878 = n8874 | n8877 ;
  assign n8879 = n8875 ^ n6729 ^ n6204 ;
  assign n8880 = n8876 | n8878 ;
  assign n8881 = ( n8089 & ~n8879 ) | ( n8089 & n8880 ) | ( ~n8879 & n8880 ) ;
  assign n8882 = n8880 | n8881 ;
  assign n8883 = n8882 ^ x2 ^ 1'b0 ;
  assign n8884 = ( n8589 & n8873 ) | ( n8589 & n8883 ) | ( n8873 & n8883 ) ;
  assign n8885 = n6597 & n8090 ;
  assign n8886 = ( n6204 & n8088 ) | ( n6204 & n8885 ) | ( n8088 & n8885 ) ;
  assign n8887 = ( ~n6729 & n8086 ) | ( ~n6729 & n8885 ) | ( n8086 & n8885 ) ;
  assign n8888 = n8885 | n8886 ;
  assign n8889 = ( n6204 & ~n6729 ) | ( n6204 & n8875 ) | ( ~n6729 & n8875 ) ;
  assign n8890 = n8887 | n8888 ;
  assign n8891 = n8889 ^ n6597 ^ n6204 ;
  assign n8892 = ( n8089 & n8890 ) | ( n8089 & n8891 ) | ( n8890 & n8891 ) ;
  assign n8893 = n8890 | n8892 ;
  assign n8894 = n6597 & n6907 ;
  assign n8895 = n8893 ^ x2 ^ 1'b0 ;
  assign n8896 = ( n8609 & n8884 ) | ( n8609 & n8895 ) | ( n8884 & n8895 ) ;
  assign n8897 = ( n6204 & n6901 ) | ( n6204 & n8894 ) | ( n6901 & n8894 ) ;
  assign n8898 = ( ~n6729 & n6906 ) | ( ~n6729 & n8894 ) | ( n6906 & n8894 ) ;
  assign n8899 = n8894 | n8897 ;
  assign n8900 = n8898 | n8899 ;
  assign n8901 = ( ~n6758 & n8556 ) | ( ~n6758 & n8863 ) | ( n8556 & n8863 ) ;
  assign n8902 = ( n6918 & n8891 ) | ( n6918 & n8900 ) | ( n8891 & n8900 ) ;
  assign n8903 = n8556 ^ n6758 ^ 1'b0 ;
  assign n8904 = n8900 | n8902 ;
  assign n8905 = n8903 ^ n8863 ^ 1'b0 ;
  assign n8906 = n6529 & n7339 ;
  assign n8907 = n8904 ^ x29 ^ 1'b0 ;
  assign n8908 = n8907 ^ n8905 ^ n8568 ;
  assign n8909 = ( n8568 & n8905 ) | ( n8568 & ~n8907 ) | ( n8905 & ~n8907 ) ;
  assign n8910 = n6529 & n6791 ;
  assign n8911 = ( ~n6729 & n6788 ) | ( ~n6729 & n8910 ) | ( n6788 & n8910 ) ;
  assign n8912 = n8910 | n8911 ;
  assign n8913 = ( ~n6170 & n6790 ) | ( ~n6170 & n8910 ) | ( n6790 & n8910 ) ;
  assign n8914 = n8912 | n8913 ;
  assign n8915 = n6789 & ~n8865 ;
  assign n8916 = n8914 | n8915 ;
  assign n8917 = ( ~n6729 & n7337 ) | ( ~n6729 & n8906 ) | ( n7337 & n8906 ) ;
  assign n8918 = n8906 | n8917 ;
  assign n8919 = ( ~n6170 & n7338 ) | ( ~n6170 & n8906 ) | ( n7338 & n8906 ) ;
  assign n8920 = n8918 | n8919 ;
  assign n8921 = ( n6716 & ~n6758 ) | ( n6716 & n8916 ) | ( ~n6758 & n8916 ) ;
  assign n8922 = n8916 ^ n6758 ^ n6716 ;
  assign n8923 = n7340 & ~n8865 ;
  assign n8924 = n8920 & ~n8923 ;
  assign n8925 = n8924 ^ n8923 ^ x20 ;
  assign n8926 = ( n8664 & n8824 ) | ( n8664 & n8925 ) | ( n8824 & n8925 ) ;
  assign n8927 = n8925 ^ n8824 ^ n8664 ;
  assign n8928 = ( ~n8901 & n8909 ) | ( ~n8901 & n8922 ) | ( n8909 & n8922 ) ;
  assign n8929 = n8922 ^ n8909 ^ n8901 ;
  assign n8930 = n6529 & n7669 ;
  assign n8931 = ( ~n6170 & n7674 ) | ( ~n6170 & n8930 ) | ( n7674 & n8930 ) ;
  assign n8932 = n8930 | n8931 ;
  assign n8933 = ( ~n6729 & n7667 ) | ( ~n6729 & n8930 ) | ( n7667 & n8930 ) ;
  assign n8934 = n8932 | n8933 ;
  assign n8935 = ( n7666 & ~n8865 ) | ( n7666 & n8934 ) | ( ~n8865 & n8934 ) ;
  assign n8936 = n8934 | n8935 ;
  assign n8937 = n8936 ^ x14 ^ 1'b0 ;
  assign n8938 = ( n8640 & n8793 ) | ( n8640 & n8937 ) | ( n8793 & n8937 ) ;
  assign n8939 = n8937 ^ n8793 ^ n8640 ;
  assign n8940 = n6529 & n6901 ;
  assign n8941 = ( ~n6170 & n6906 ) | ( ~n6170 & n8940 ) | ( n6906 & n8940 ) ;
  assign n8942 = n8940 | n8941 ;
  assign n8943 = ( ~n6729 & n6907 ) | ( ~n6729 & n8940 ) | ( n6907 & n8940 ) ;
  assign n8944 = n8942 | n8943 ;
  assign n8945 = n6918 & ~n8865 ;
  assign n8946 = n8944 | n8945 ;
  assign n8947 = n8946 ^ x29 ^ 1'b0 ;
  assign n8948 = n8947 ^ n8831 ^ n8536 ;
  assign n8949 = ( n8536 & n8831 ) | ( n8536 & n8947 ) | ( n8831 & n8947 ) ;
  assign n8950 = n6204 & n6907 ;
  assign n8951 = ( n6529 & n6906 ) | ( n6529 & n8950 ) | ( n6906 & n8950 ) ;
  assign n8952 = n8950 | n8951 ;
  assign n8953 = ( ~n6729 & n6901 ) | ( ~n6729 & n8950 ) | ( n6901 & n8950 ) ;
  assign n8954 = n8952 | n8953 ;
  assign n8955 = n6918 & ~n8879 ;
  assign n8956 = n8954 | n8955 ;
  assign n8957 = n8956 ^ x29 ^ 1'b0 ;
  assign n8958 = ( n8567 & n8949 ) | ( n8567 & n8957 ) | ( n8949 & n8957 ) ;
  assign n8959 = n8957 ^ n8949 ^ n8567 ;
  assign n8960 = n6529 & n7036 ;
  assign n8961 = ( ~n6729 & n7037 ) | ( ~n6729 & n8960 ) | ( n7037 & n8960 ) ;
  assign n8962 = n8960 | n8961 ;
  assign n8963 = ( ~n6170 & n7052 ) | ( ~n6170 & n8960 ) | ( n7052 & n8960 ) ;
  assign n8964 = n8962 | n8963 ;
  assign n8965 = n7035 & ~n8865 ;
  assign n8966 = n8964 | n8965 ;
  assign n8967 = n8966 ^ x26 ^ 1'b0 ;
  assign n8968 = ( n8395 & n8760 ) | ( n8395 & n8967 ) | ( n8760 & n8967 ) ;
  assign n8969 = n8967 ^ n8760 ^ n8395 ;
  assign n8970 = n6529 & n7485 ;
  assign n8971 = ( ~n6729 & n7486 ) | ( ~n6729 & n8970 ) | ( n7486 & n8970 ) ;
  assign n8972 = n8970 | n8971 ;
  assign n8973 = ( ~n6170 & n7493 ) | ( ~n6170 & n8970 ) | ( n7493 & n8970 ) ;
  assign n8974 = n8972 | n8973 ;
  assign n8975 = n7487 & ~n8865 ;
  assign n8976 = n8974 | n8975 ;
  assign n8977 = n8976 ^ x17 ^ 1'b0 ;
  assign n8978 = ( n8674 & n8803 ) | ( n8674 & n8977 ) | ( n8803 & n8977 ) ;
  assign n8979 = n8977 ^ n8803 ^ n8674 ;
  assign n8980 = n6529 & n7829 ;
  assign n8981 = ( ~n6170 & n7833 ) | ( ~n6170 & n8980 ) | ( n7833 & n8980 ) ;
  assign n8982 = n8980 | n8981 ;
  assign n8983 = ( ~n6729 & n7834 ) | ( ~n6729 & n8980 ) | ( n7834 & n8980 ) ;
  assign n8984 = n8982 | n8983 ;
  assign n8985 = n7838 & ~n8865 ;
  assign n8986 = n8984 | n8985 ;
  assign n8987 = n8986 ^ x11 ^ 1'b0 ;
  assign n8988 = ( n8676 & n8846 ) | ( n8676 & n8987 ) | ( n8846 & n8987 ) ;
  assign n8989 = n8987 ^ n8846 ^ n8676 ;
  assign n8990 = n6529 & n7932 ;
  assign n8991 = ( ~n6170 & n7943 ) | ( ~n6170 & n8990 ) | ( n7943 & n8990 ) ;
  assign n8992 = n8990 | n8991 ;
  assign n8993 = ( ~n6729 & n7929 ) | ( ~n6729 & n8990 ) | ( n7929 & n8990 ) ;
  assign n8994 = n8992 | n8993 ;
  assign n8995 = n7930 & ~n8865 ;
  assign n8996 = n8994 | n8995 ;
  assign n8997 = n8996 ^ x8 ^ 1'b0 ;
  assign n8998 = ( n8699 & n8857 ) | ( n8699 & n8997 ) | ( n8857 & n8997 ) ;
  assign n8999 = n8997 ^ n8857 ^ n8699 ;
  assign n9000 = n6529 & n7192 ;
  assign n9001 = ( ~n6729 & n7188 ) | ( ~n6729 & n9000 ) | ( n7188 & n9000 ) ;
  assign n9002 = n9000 | n9001 ;
  assign n9003 = ( ~n6170 & n7190 ) | ( ~n6170 & n9000 ) | ( n7190 & n9000 ) ;
  assign n9004 = n9002 | n9003 ;
  assign n9005 = n7196 & ~n8865 ;
  assign n9006 = n9004 | n9005 ;
  assign n9007 = n6529 & n8029 ;
  assign n9008 = ( ~n6170 & n8037 ) | ( ~n6170 & n9007 ) | ( n8037 & n9007 ) ;
  assign n9009 = n9007 | n9008 ;
  assign n9010 = n8034 & ~n8865 ;
  assign n9011 = ( ~n6729 & n8033 ) | ( ~n6729 & n9007 ) | ( n8033 & n9007 ) ;
  assign n9012 = n9009 | n9011 ;
  assign n9013 = n6759 ^ n6758 ^ x14 ;
  assign n9014 = n9010 | n9012 ;
  assign n9015 = n6789 & ~n8879 ;
  assign n9016 = n9006 ^ x23 ^ 1'b0 ;
  assign n9017 = ( x14 & ~n6758 ) | ( x14 & n6759 ) | ( ~n6758 & n6759 ) ;
  assign n9018 = n9014 ^ x5 ^ 1'b0 ;
  assign n9019 = n9018 ^ n8630 ^ n8608 ;
  assign n9020 = ( n8608 & n8630 ) | ( n8608 & n9018 ) | ( n8630 & n9018 ) ;
  assign n9021 = ~n6729 & n6791 ;
  assign n9022 = n9016 ^ n8749 ^ n8494 ;
  assign n9023 = ( n8494 & ~n8749 ) | ( n8494 & n9016 ) | ( ~n8749 & n9016 ) ;
  assign n9024 = ( n6204 & n6788 ) | ( n6204 & n9021 ) | ( n6788 & n9021 ) ;
  assign n9025 = n9021 | n9024 ;
  assign n9026 = n7196 & ~n8879 ;
  assign n9027 = ( n6529 & n6790 ) | ( n6529 & n9021 ) | ( n6790 & n9021 ) ;
  assign n9028 = n9025 | n9027 ;
  assign n9029 = n9015 | n9028 ;
  assign n9030 = n9029 ^ n9013 ^ n8921 ;
  assign n9031 = ( n8921 & n9013 ) | ( n8921 & n9029 ) | ( n9013 & n9029 ) ;
  assign n9032 = n6204 & n7337 ;
  assign n9033 = ( ~n6729 & n7339 ) | ( ~n6729 & n9032 ) | ( n7339 & n9032 ) ;
  assign n9034 = ( n6529 & n7338 ) | ( n6529 & n9032 ) | ( n7338 & n9032 ) ;
  assign n9035 = n9032 | n9034 ;
  assign n9036 = n9033 | n9035 ;
  assign n9037 = n7340 & ~n8879 ;
  assign n9038 = n9036 | n9037 ;
  assign n9039 = n6204 & n7188 ;
  assign n9040 = n9038 ^ x20 ^ 1'b0 ;
  assign n9041 = ( n6529 & n7190 ) | ( n6529 & n9039 ) | ( n7190 & n9039 ) ;
  assign n9042 = n9039 | n9041 ;
  assign n9043 = ( ~n6729 & n7192 ) | ( ~n6729 & n9039 ) | ( n7192 & n9039 ) ;
  assign n9044 = n9042 | n9043 ;
  assign n9045 = ( n8653 & n8665 ) | ( n8653 & n9040 ) | ( n8665 & n9040 ) ;
  assign n9046 = n9026 | n9044 ;
  assign n9047 = n9046 ^ x23 ^ 1'b0 ;
  assign n9048 = ( n8772 & n9023 ) | ( n8772 & n9047 ) | ( n9023 & n9047 ) ;
  assign n9049 = n9047 ^ n9023 ^ n8772 ;
  assign n9050 = n9040 ^ n8665 ^ n8653 ;
  assign n9051 = n6204 & n7834 ;
  assign n9052 = ( n6529 & n7833 ) | ( n6529 & n9051 ) | ( n7833 & n9051 ) ;
  assign n9053 = n9051 | n9052 ;
  assign n9054 = ( ~n6729 & n7829 ) | ( ~n6729 & n9051 ) | ( n7829 & n9051 ) ;
  assign n9055 = n9053 | n9054 ;
  assign n9056 = ( n7838 & ~n8879 ) | ( n7838 & n9055 ) | ( ~n8879 & n9055 ) ;
  assign n9057 = n9055 | n9056 ;
  assign n9058 = n9057 ^ x11 ^ 1'b0 ;
  assign n9059 = n9058 ^ n8988 ^ n8729 ;
  assign n9060 = ( n8729 & n8988 ) | ( n8729 & n9058 ) | ( n8988 & n9058 ) ;
  assign n9061 = n6204 & n7929 ;
  assign n9062 = ( n6529 & n7943 ) | ( n6529 & n9061 ) | ( n7943 & n9061 ) ;
  assign n9063 = n9061 | n9062 ;
  assign n9064 = ( ~n6729 & n7932 ) | ( ~n6729 & n9061 ) | ( n7932 & n9061 ) ;
  assign n9065 = n9063 | n9064 ;
  assign n9066 = ( n7930 & ~n8879 ) | ( n7930 & n9065 ) | ( ~n8879 & n9065 ) ;
  assign n9067 = n9065 | n9066 ;
  assign n9068 = n9067 ^ x8 ^ 1'b0 ;
  assign n9069 = n9068 ^ n8998 ^ n8738 ;
  assign n9070 = ( n8738 & n8998 ) | ( n8738 & n9068 ) | ( n8998 & n9068 ) ;
  assign n9071 = n6204 & n7667 ;
  assign n9072 = ( n6529 & n7674 ) | ( n6529 & n9071 ) | ( n7674 & n9071 ) ;
  assign n9073 = n9071 | n9072 ;
  assign n9074 = ( ~n6729 & n7669 ) | ( ~n6729 & n9071 ) | ( n7669 & n9071 ) ;
  assign n9075 = n9073 | n9074 ;
  assign n9076 = ( n7666 & ~n8879 ) | ( n7666 & n9075 ) | ( ~n8879 & n9075 ) ;
  assign n9077 = n9075 | n9076 ;
  assign n9078 = n9077 ^ x14 ^ 1'b0 ;
  assign n9079 = ( ~n8719 & n8938 ) | ( ~n8719 & n9078 ) | ( n8938 & n9078 ) ;
  assign n9080 = n9078 ^ n8938 ^ n8719 ;
  assign n9081 = n6204 & n7037 ;
  assign n9082 = ( n6529 & n7052 ) | ( n6529 & n9081 ) | ( n7052 & n9081 ) ;
  assign n9083 = n9081 | n9082 ;
  assign n9084 = ( ~n6729 & n7036 ) | ( ~n6729 & n9081 ) | ( n7036 & n9081 ) ;
  assign n9085 = n9083 | n9084 ;
  assign n9086 = n7035 & ~n8879 ;
  assign n9087 = n9085 & ~n9086 ;
  assign n9088 = n9087 ^ n9086 ^ x26 ;
  assign n9089 = n9088 ^ n8968 ^ n8682 ;
  assign n9090 = ( n8682 & n8968 ) | ( n8682 & n9088 ) | ( n8968 & n9088 ) ;
  assign n9091 = n6204 & n8033 ;
  assign n9092 = ( n6529 & n8037 ) | ( n6529 & n9091 ) | ( n8037 & n9091 ) ;
  assign n9093 = n9091 | n9092 ;
  assign n9094 = ( ~n6729 & n8029 ) | ( ~n6729 & n9091 ) | ( n8029 & n9091 ) ;
  assign n9095 = n9093 | n9094 ;
  assign n9096 = ( n8034 & ~n8879 ) | ( n8034 & n9095 ) | ( ~n8879 & n9095 ) ;
  assign n9097 = n9095 | n9096 ;
  assign n9098 = n6204 & n7486 ;
  assign n9099 = ( n6529 & n7493 ) | ( n6529 & n9098 ) | ( n7493 & n9098 ) ;
  assign n9100 = n9098 | n9099 ;
  assign n9101 = ( ~n6729 & n7485 ) | ( ~n6729 & n9098 ) | ( n7485 & n9098 ) ;
  assign n9102 = n9100 | n9101 ;
  assign n9103 = n7487 & ~n8879 ;
  assign n9104 = n6597 & n7486 ;
  assign n9105 = n9097 ^ x5 ^ 1'b0 ;
  assign n9106 = n9102 | n9103 ;
  assign n9107 = n9106 ^ x17 ^ 1'b0 ;
  assign n9108 = ( ~n8709 & n8978 ) | ( ~n8709 & n9107 ) | ( n8978 & n9107 ) ;
  assign n9109 = n9107 ^ n8978 ^ n8709 ;
  assign n9110 = ( n8689 & n9020 ) | ( n8689 & n9105 ) | ( n9020 & n9105 ) ;
  assign n9111 = n7487 & n8891 ;
  assign n9112 = n9105 ^ n9020 ^ n8689 ;
  assign n9113 = ( n6204 & n7485 ) | ( n6204 & n9104 ) | ( n7485 & n9104 ) ;
  assign n9114 = n9104 | n9113 ;
  assign n9115 = ( ~n6729 & n7493 ) | ( ~n6729 & n9104 ) | ( n7493 & n9104 ) ;
  assign n9116 = n9114 | n9115 ;
  assign n9117 = n9111 | n9116 ;
  assign n9118 = n9117 ^ x17 ^ 1'b0 ;
  assign n9119 = ( n8823 & n9108 ) | ( n8823 & n9118 ) | ( n9108 & n9118 ) ;
  assign n9120 = n9118 ^ n9108 ^ n8823 ;
  assign n9121 = n6597 & n7188 ;
  assign n9122 = ( ~n6729 & n7190 ) | ( ~n6729 & n9121 ) | ( n7190 & n9121 ) ;
  assign n9123 = n6597 & n7929 ;
  assign n9124 = ( n6204 & n7192 ) | ( n6204 & n9121 ) | ( n7192 & n9121 ) ;
  assign n9125 = n9121 | n9124 ;
  assign n9126 = ( n6204 & n7932 ) | ( n6204 & n9123 ) | ( n7932 & n9123 ) ;
  assign n9127 = n9122 | n9125 ;
  assign n9128 = n7196 & n8891 ;
  assign n9129 = n9127 | n9128 ;
  assign n9130 = n9129 ^ x23 ^ 1'b0 ;
  assign n9131 = ( n8773 & ~n8813 ) | ( n8773 & n9130 ) | ( ~n8813 & n9130 ) ;
  assign n9132 = n9123 | n9126 ;
  assign n9133 = ( ~n6729 & n7943 ) | ( ~n6729 & n9123 ) | ( n7943 & n9123 ) ;
  assign n9134 = n9132 | n9133 ;
  assign n9135 = ( n7930 & n8891 ) | ( n7930 & n9134 ) | ( n8891 & n9134 ) ;
  assign n9136 = n9134 | n9135 ;
  assign n9137 = n9136 ^ x8 ^ 1'b0 ;
  assign n9138 = ( n8845 & n9070 ) | ( n8845 & n9137 ) | ( n9070 & n9137 ) ;
  assign n9139 = n9137 ^ n9070 ^ n8845 ;
  assign n9140 = n6597 & n7667 ;
  assign n9141 = ( n6204 & n7669 ) | ( n6204 & n9140 ) | ( n7669 & n9140 ) ;
  assign n9142 = n9140 | n9141 ;
  assign n9143 = ( ~n6729 & n7674 ) | ( ~n6729 & n9140 ) | ( n7674 & n9140 ) ;
  assign n9144 = n9130 ^ n8813 ^ n8773 ;
  assign n9145 = n6597 & n7834 ;
  assign n9146 = ( ~n6729 & n7833 ) | ( ~n6729 & n9145 ) | ( n7833 & n9145 ) ;
  assign n9147 = n9142 | n9143 ;
  assign n9148 = ( n6204 & n7829 ) | ( n6204 & n9145 ) | ( n7829 & n9145 ) ;
  assign n9149 = n9145 | n9148 ;
  assign n9150 = n9146 | n9149 ;
  assign n9151 = ( n7838 & n8891 ) | ( n7838 & n9150 ) | ( n8891 & n9150 ) ;
  assign n9152 = ( n7666 & n8891 ) | ( n7666 & n9147 ) | ( n8891 & n9147 ) ;
  assign n9153 = n9147 | n9152 ;
  assign n9154 = n9153 ^ x14 ^ 1'b0 ;
  assign n9155 = n9154 ^ n9079 ^ n8804 ;
  assign n9156 = ( ~n8804 & n9079 ) | ( ~n8804 & n9154 ) | ( n9079 & n9154 ) ;
  assign n9157 = n9150 | n9151 ;
  assign n9158 = n9157 ^ x11 ^ 1'b0 ;
  assign n9159 = n9158 ^ n9060 ^ n8794 ;
  assign n9160 = n6597 & n8033 ;
  assign n9161 = ( n6204 & n8029 ) | ( n6204 & n9160 ) | ( n8029 & n9160 ) ;
  assign n9162 = n9160 | n9161 ;
  assign n9163 = ( n8794 & n9060 ) | ( n8794 & n9158 ) | ( n9060 & n9158 ) ;
  assign n9164 = ( ~n6729 & n8037 ) | ( ~n6729 & n9160 ) | ( n8037 & n9160 ) ;
  assign n9165 = n6597 & n7337 ;
  assign n9166 = n6204 & n6791 ;
  assign n9167 = n9162 | n9164 ;
  assign n9168 = ( n6597 & n6788 ) | ( n6597 & n9166 ) | ( n6788 & n9166 ) ;
  assign n9169 = n9166 | n9168 ;
  assign n9170 = ( ~n6729 & n6790 ) | ( ~n6729 & n9166 ) | ( n6790 & n9166 ) ;
  assign n9171 = n9169 | n9170 ;
  assign n9172 = ( n6204 & n7339 ) | ( n6204 & n9165 ) | ( n7339 & n9165 ) ;
  assign n9173 = n9165 | n9172 ;
  assign n9174 = ( ~n6729 & n7338 ) | ( ~n6729 & n9165 ) | ( n7338 & n9165 ) ;
  assign n9175 = n9173 | n9174 ;
  assign n9176 = n6789 & ~n8891 ;
  assign n9177 = ( n6789 & n9171 ) | ( n6789 & ~n9176 ) | ( n9171 & ~n9176 ) ;
  assign n9178 = n7340 & n8891 ;
  assign n9179 = n9175 | n9178 ;
  assign n9180 = n7035 & n8891 ;
  assign n9181 = n9179 ^ x20 ^ 1'b0 ;
  assign n9182 = ( n8034 & n8891 ) | ( n8034 & n9167 ) | ( n8891 & n9167 ) ;
  assign n9183 = n9167 | n9182 ;
  assign n9184 = ( n8654 & n8783 ) | ( n8654 & n9181 ) | ( n8783 & n9181 ) ;
  assign n9185 = n9181 ^ n8783 ^ n8654 ;
  assign n9186 = n6597 & n7037 ;
  assign n9187 = ( n6204 & n7036 ) | ( n6204 & n9186 ) | ( n7036 & n9186 ) ;
  assign n9188 = ( ~n6729 & n7052 ) | ( ~n6729 & n9186 ) | ( n7052 & n9186 ) ;
  assign n9189 = n9183 ^ x5 ^ 1'b0 ;
  assign n9190 = n9186 | n9187 ;
  assign n9191 = n9189 ^ n9110 ^ n8856 ;
  assign n9192 = ( n8856 & n9110 ) | ( n8856 & n9189 ) | ( n9110 & n9189 ) ;
  assign n9193 = n9188 | n9190 ;
  assign n9194 = n9180 | n9193 ;
  assign n9195 = n9194 ^ x26 ^ 1'b0 ;
  assign n9196 = n9195 ^ n8836 ^ n8666 ;
  assign n9197 = ( n8666 & n8836 ) | ( n8666 & n9195 ) | ( n8836 & n9195 ) ;
  assign n9198 = ( n6204 & n6597 ) | ( n6204 & n8889 ) | ( n6597 & n8889 ) ;
  assign n9199 = n6596 & n8090 ;
  assign n9200 = ( n6597 & n8088 ) | ( n6597 & n9199 ) | ( n8088 & n9199 ) ;
  assign n9201 = n9199 | n9200 ;
  assign n9202 = ( n6204 & n8086 ) | ( n6204 & n9199 ) | ( n8086 & n9199 ) ;
  assign n9203 = n9201 | n9202 ;
  assign n9204 = n9198 ^ n6597 ^ n6596 ;
  assign n9205 = ( n8089 & n9203 ) | ( n8089 & n9204 ) | ( n9203 & n9204 ) ;
  assign n9206 = n9203 | n9205 ;
  assign n9207 = n9206 ^ x2 ^ 1'b0 ;
  assign n9208 = ( n8896 & n9019 ) | ( n8896 & n9207 ) | ( n9019 & n9207 ) ;
  assign n9209 = n9177 ^ n9017 ^ n6819 ;
  assign n9210 = n6596 & n7188 ;
  assign n9211 = ( n6819 & n9017 ) | ( n6819 & ~n9177 ) | ( n9017 & ~n9177 ) ;
  assign n9212 = n6596 & n7929 ;
  assign n9213 = ( n6597 & n7192 ) | ( n6597 & n9210 ) | ( n7192 & n9210 ) ;
  assign n9214 = n9210 | n9213 ;
  assign n9215 = ( n6204 & n7190 ) | ( n6204 & n9210 ) | ( n7190 & n9210 ) ;
  assign n9216 = n9214 | n9215 ;
  assign n9217 = n7196 & n9204 ;
  assign n9218 = n9216 | n9217 ;
  assign n9219 = ( n6597 & n7932 ) | ( n6597 & n9212 ) | ( n7932 & n9212 ) ;
  assign n9220 = n9212 | n9219 ;
  assign n9221 = ( n6204 & n7943 ) | ( n6204 & n9212 ) | ( n7943 & n9212 ) ;
  assign n9222 = n9220 | n9221 ;
  assign n9223 = n9211 ^ n6819 ^ n6629 ;
  assign n9224 = ( n6629 & n6819 ) | ( n6629 & ~n9211 ) | ( n6819 & ~n9211 ) ;
  assign n9225 = ( n6596 & n6597 ) | ( n6596 & n9198 ) | ( n6597 & n9198 ) ;
  assign n9226 = n9218 ^ x23 ^ 1'b0 ;
  assign n9227 = ( n8814 & n8969 ) | ( n8814 & n9226 ) | ( n8969 & n9226 ) ;
  assign n9228 = n9226 ^ n8969 ^ n8814 ;
  assign n9229 = ( n7930 & n9204 ) | ( n7930 & n9222 ) | ( n9204 & n9222 ) ;
  assign n9230 = n6596 & n7037 ;
  assign n9231 = n9222 | n9229 ;
  assign n9232 = ( x17 & n6629 ) | ( x17 & ~n6691 ) | ( n6629 & ~n6691 ) ;
  assign n9233 = n6691 ^ n6629 ^ x17 ;
  assign n9234 = n9231 ^ x8 ^ 1'b0 ;
  assign n9235 = ( n8989 & n9138 ) | ( n8989 & n9234 ) | ( n9138 & n9234 ) ;
  assign n9236 = n9234 ^ n9138 ^ n8989 ;
  assign n9237 = ( n6597 & n7036 ) | ( n6597 & n9230 ) | ( n7036 & n9230 ) ;
  assign n9238 = n7035 & n9204 ;
  assign n9239 = n9230 | n9237 ;
  assign n9240 = ( n6204 & n7052 ) | ( n6204 & n9230 ) | ( n7052 & n9230 ) ;
  assign n9241 = n9239 | n9240 ;
  assign n9242 = n9238 | n9241 ;
  assign n9243 = n9242 ^ x26 ^ 1'b0 ;
  assign n9244 = n9243 ^ n8948 ^ n8835 ;
  assign n9245 = ( n8835 & n8948 ) | ( n8835 & n9243 ) | ( n8948 & n9243 ) ;
  assign n9246 = n6596 & n8033 ;
  assign n9247 = ( n6597 & n8029 ) | ( n6597 & n9246 ) | ( n8029 & n9246 ) ;
  assign n9248 = n9246 | n9247 ;
  assign n9249 = ( n6204 & n8037 ) | ( n6204 & n9246 ) | ( n8037 & n9246 ) ;
  assign n9250 = n9248 | n9249 ;
  assign n9251 = n6596 & n7036 ;
  assign n9252 = ( n8034 & n9204 ) | ( n8034 & n9250 ) | ( n9204 & n9250 ) ;
  assign n9253 = n9250 | n9252 ;
  assign n9254 = ( n6597 & n7052 ) | ( n6597 & n9251 ) | ( n7052 & n9251 ) ;
  assign n9255 = n9251 | n9254 ;
  assign n9256 = n9253 ^ x5 ^ 1'b0 ;
  assign n9257 = ( ~n6728 & n7037 ) | ( ~n6728 & n9251 ) | ( n7037 & n9251 ) ;
  assign n9258 = n9255 | n9257 ;
  assign n9259 = n9256 ^ n9192 ^ n8999 ;
  assign n9260 = ( n8999 & n9192 ) | ( n8999 & n9256 ) | ( n9192 & n9256 ) ;
  assign n9261 = n9225 ^ n6728 ^ n6596 ;
  assign n9262 = n7035 & ~n9261 ;
  assign n9263 = n9258 & ~n9262 ;
  assign n9264 = n9263 ^ n9262 ^ x26 ;
  assign n9265 = ( n8959 & n9245 ) | ( n8959 & n9264 ) | ( n9245 & n9264 ) ;
  assign n9266 = n9264 ^ n9245 ^ n8959 ;
  assign n9267 = n6596 & n8088 ;
  assign n9268 = ( n6597 & n8086 ) | ( n6597 & n9267 ) | ( n8086 & n9267 ) ;
  assign n9269 = n9267 | n9268 ;
  assign n9270 = ( ~n6728 & n8090 ) | ( ~n6728 & n9267 ) | ( n8090 & n9267 ) ;
  assign n9271 = n9269 | n9270 ;
  assign n9272 = n8089 & ~n9261 ;
  assign n9273 = n9271 | n9272 ;
  assign n9274 = n6596 & n7932 ;
  assign n9275 = n9273 ^ x2 ^ 1'b0 ;
  assign n9276 = ( n9112 & n9208 ) | ( n9112 & n9275 ) | ( n9208 & n9275 ) ;
  assign n9277 = ( n6597 & n7943 ) | ( n6597 & n9274 ) | ( n7943 & n9274 ) ;
  assign n9278 = ( ~n6728 & n7929 ) | ( ~n6728 & n9274 ) | ( n7929 & n9274 ) ;
  assign n9279 = n9274 | n9277 ;
  assign n9280 = n7930 & ~n9261 ;
  assign n9281 = n9278 | n9279 ;
  assign n9282 = n9280 | n9281 ;
  assign n9283 = n7340 & n9204 ;
  assign n9284 = n9282 ^ x8 ^ 1'b0 ;
  assign n9285 = ( n9059 & n9235 ) | ( n9059 & n9284 ) | ( n9235 & n9284 ) ;
  assign n9286 = n9284 ^ n9235 ^ n9059 ;
  assign n9287 = n6596 & n7337 ;
  assign n9288 = ( n6597 & n7339 ) | ( n6597 & n9287 ) | ( n7339 & n9287 ) ;
  assign n9289 = n9287 | n9288 ;
  assign n9290 = ( n6204 & n7338 ) | ( n6204 & n9287 ) | ( n7338 & n9287 ) ;
  assign n9291 = n9289 | n9290 ;
  assign n9292 = n9283 | n9291 ;
  assign n9293 = n9292 ^ x20 ^ 1'b0 ;
  assign n9294 = n9293 ^ n9022 ^ n8784 ;
  assign n9295 = ( n8784 & ~n9022 ) | ( n8784 & n9293 ) | ( ~n9022 & n9293 ) ;
  assign n9296 = n6596 & n7834 ;
  assign n9297 = ( n6597 & n7829 ) | ( n6597 & n9296 ) | ( n7829 & n9296 ) ;
  assign n9298 = n9296 | n9297 ;
  assign n9299 = ( n6204 & n7833 ) | ( n6204 & n9296 ) | ( n7833 & n9296 ) ;
  assign n9300 = n9298 | n9299 ;
  assign n9301 = n7838 & n9204 ;
  assign n9302 = n9300 | n9301 ;
  assign n9303 = n9302 ^ x11 ^ 1'b0 ;
  assign n9304 = n9303 ^ n9163 ^ n8939 ;
  assign n9305 = ( n8939 & n9163 ) | ( n8939 & n9303 ) | ( n9163 & n9303 ) ;
  assign n9306 = n6596 & n7829 ;
  assign n9307 = ( n6597 & n7833 ) | ( n6597 & n9306 ) | ( n7833 & n9306 ) ;
  assign n9308 = n9306 | n9307 ;
  assign n9309 = ( ~n6728 & n7834 ) | ( ~n6728 & n9306 ) | ( n7834 & n9306 ) ;
  assign n9310 = n9308 | n9309 ;
  assign n9311 = n7838 & ~n9261 ;
  assign n9312 = n9310 | n9311 ;
  assign n9313 = n9312 ^ x11 ^ 1'b0 ;
  assign n9314 = ( ~n9080 & n9305 ) | ( ~n9080 & n9313 ) | ( n9305 & n9313 ) ;
  assign n9315 = n9313 ^ n9305 ^ n9080 ;
  assign n9316 = n6596 & n7339 ;
  assign n9317 = ( n6597 & n7338 ) | ( n6597 & n9316 ) | ( n7338 & n9316 ) ;
  assign n9318 = n9316 | n9317 ;
  assign n9319 = ( ~n6728 & n7337 ) | ( ~n6728 & n9316 ) | ( n7337 & n9316 ) ;
  assign n9320 = n9318 | n9319 ;
  assign n9321 = ( n7340 & ~n9261 ) | ( n7340 & n9320 ) | ( ~n9261 & n9320 ) ;
  assign n9322 = n9320 | n9321 ;
  assign n9323 = n9322 ^ x20 ^ 1'b0 ;
  assign n9324 = ( n9049 & n9295 ) | ( n9049 & n9323 ) | ( n9295 & n9323 ) ;
  assign n9325 = n9323 ^ n9295 ^ n9049 ;
  assign n9326 = n6596 & n7486 ;
  assign n9327 = ( n6597 & n7485 ) | ( n6597 & n9326 ) | ( n7485 & n9326 ) ;
  assign n9328 = n9326 | n9327 ;
  assign n9329 = ( n6204 & n7493 ) | ( n6204 & n9326 ) | ( n7493 & n9326 ) ;
  assign n9330 = n9328 | n9329 ;
  assign n9331 = n7487 & n9204 ;
  assign n9332 = n9330 | n9331 ;
  assign n9333 = n9332 ^ x17 ^ 1'b0 ;
  assign n9334 = ( n8927 & n9119 ) | ( n8927 & n9333 ) | ( n9119 & n9333 ) ;
  assign n9335 = n9333 ^ n9119 ^ n8927 ;
  assign n9336 = n6596 & n7667 ;
  assign n9337 = ( n6597 & n7669 ) | ( n6597 & n9336 ) | ( n7669 & n9336 ) ;
  assign n9338 = n9336 | n9337 ;
  assign n9339 = ( n6204 & n7674 ) | ( n6204 & n9336 ) | ( n7674 & n9336 ) ;
  assign n9340 = n9338 | n9339 ;
  assign n9341 = ( n7666 & n9204 ) | ( n7666 & n9340 ) | ( n9204 & n9340 ) ;
  assign n9342 = n9340 | n9341 ;
  assign n9343 = n9342 ^ x14 ^ 1'b0 ;
  assign n9344 = n9343 ^ n9156 ^ n8979 ;
  assign n9345 = ( n8979 & n9156 ) | ( n8979 & n9343 ) | ( n9156 & n9343 ) ;
  assign n9346 = n6596 & n7669 ;
  assign n9347 = ( n6597 & n7674 ) | ( n6597 & n9346 ) | ( n7674 & n9346 ) ;
  assign n9348 = n9346 | n9347 ;
  assign n9349 = ( ~n6728 & n7667 ) | ( ~n6728 & n9346 ) | ( n7667 & n9346 ) ;
  assign n9350 = n9348 | n9349 ;
  assign n9351 = ( n7666 & ~n9261 ) | ( n7666 & n9350 ) | ( ~n9261 & n9350 ) ;
  assign n9352 = n9350 | n9351 ;
  assign n9353 = n9352 ^ x14 ^ 1'b0 ;
  assign n9354 = n9353 ^ n9345 ^ n9109 ;
  assign n9355 = ( ~n9109 & n9345 ) | ( ~n9109 & n9353 ) | ( n9345 & n9353 ) ;
  assign n9356 = n6789 & ~n9261 ;
  assign n9357 = ( n6596 & n6791 ) | ( n6596 & n9356 ) | ( n6791 & n9356 ) ;
  assign n9358 = n9356 | n9357 ;
  assign n9359 = ( n6597 & n6790 ) | ( n6597 & n9356 ) | ( n6790 & n9356 ) ;
  assign n9360 = n9358 | n9359 ;
  assign n9361 = n6728 & n6788 ;
  assign n9362 = ( n6788 & n9360 ) | ( n6788 & ~n9361 ) | ( n9360 & ~n9361 ) ;
  assign n9363 = ( n9224 & n9233 ) | ( n9224 & n9362 ) | ( n9233 & n9362 ) ;
  assign n9364 = n9362 ^ n9233 ^ n9224 ;
  assign n9365 = n6596 & n6907 ;
  assign n9366 = ( n6597 & n6901 ) | ( n6597 & n9365 ) | ( n6901 & n9365 ) ;
  assign n9367 = n9365 | n9366 ;
  assign n9368 = ( n6204 & n6906 ) | ( n6204 & n9365 ) | ( n6906 & n9365 ) ;
  assign n9369 = n9367 | n9368 ;
  assign n9370 = n6789 & n9204 ;
  assign n9371 = ( n6204 & n6790 ) | ( n6204 & n9370 ) | ( n6790 & n9370 ) ;
  assign n9372 = ( n6918 & n9204 ) | ( n6918 & n9369 ) | ( n9204 & n9369 ) ;
  assign n9373 = n9369 | n9372 ;
  assign n9374 = ( n6597 & n6791 ) | ( n6597 & n9370 ) | ( n6791 & n9370 ) ;
  assign n9375 = n9370 | n9374 ;
  assign n9376 = n9371 | n9375 ;
  assign n9377 = n6596 & n8029 ;
  assign n9378 = n6596 & n7192 ;
  assign n9379 = ( n6597 & n8037 ) | ( n6597 & n9377 ) | ( n8037 & n9377 ) ;
  assign n9380 = n9377 | n9379 ;
  assign n9381 = ( ~n6728 & n8033 ) | ( ~n6728 & n9377 ) | ( n8033 & n9377 ) ;
  assign n9382 = n9380 | n9381 ;
  assign n9383 = n8034 & ~n9261 ;
  assign n9384 = n9382 | n9383 ;
  assign n9385 = ( n6597 & n7190 ) | ( n6597 & n9378 ) | ( n7190 & n9378 ) ;
  assign n9386 = n9378 | n9385 ;
  assign n9387 = ( n6596 & ~n6728 ) | ( n6596 & n9225 ) | ( ~n6728 & n9225 ) ;
  assign n9388 = n9384 ^ x5 ^ 1'b0 ;
  assign n9389 = ( ~n6728 & n7188 ) | ( ~n6728 & n9378 ) | ( n7188 & n9378 ) ;
  assign n9390 = n9386 | n9389 ;
  assign n9391 = n7196 & ~n9261 ;
  assign n9392 = n9390 | n9391 ;
  assign n9393 = n9392 ^ x23 ^ 1'b0 ;
  assign n9394 = n9393 ^ n9227 ^ n9089 ;
  assign n9395 = ( n9089 & n9227 ) | ( n9089 & n9393 ) | ( n9227 & n9393 ) ;
  assign n9396 = ( n9069 & n9260 ) | ( n9069 & n9388 ) | ( n9260 & n9388 ) ;
  assign n9397 = n6596 & n7485 ;
  assign n9398 = n9388 ^ n9260 ^ n9069 ;
  assign n9399 = ( n6597 & n7493 ) | ( n6597 & n9397 ) | ( n7493 & n9397 ) ;
  assign n9400 = n9397 | n9399 ;
  assign n9401 = ( ~n6728 & n7486 ) | ( ~n6728 & n9397 ) | ( n7486 & n9397 ) ;
  assign n9402 = n9400 | n9401 ;
  assign n9403 = n6371 & n7337 ;
  assign n9404 = n7487 & ~n9261 ;
  assign n9405 = n9402 | n9404 ;
  assign n9406 = n9405 ^ x17 ^ 1'b0 ;
  assign n9407 = ( n6596 & n7338 ) | ( n6596 & n9403 ) | ( n7338 & n9403 ) ;
  assign n9408 = n9403 | n9407 ;
  assign n9409 = ( ~n6728 & n7339 ) | ( ~n6728 & n9403 ) | ( n7339 & n9403 ) ;
  assign n9410 = n9408 | n9409 ;
  assign n9411 = n9406 ^ n9050 ^ n8926 ;
  assign n9412 = ( n8926 & n9050 ) | ( n8926 & n9406 ) | ( n9050 & n9406 ) ;
  assign n9413 = n9387 ^ n6728 ^ n6371 ;
  assign n9414 = n6596 & n6901 ;
  assign n9415 = ( n6597 & n6906 ) | ( n6597 & n9414 ) | ( n6906 & n9414 ) ;
  assign n9416 = n6918 & ~n9261 ;
  assign n9417 = n9414 | n9415 ;
  assign n9418 = ( ~n6728 & n6907 ) | ( ~n6728 & n9414 ) | ( n6907 & n9414 ) ;
  assign n9419 = n9417 | n9418 ;
  assign n9420 = n9416 | n9419 ;
  assign n9421 = n6371 & n8090 ;
  assign n9422 = ( n6596 & n8086 ) | ( n6596 & n9421 ) | ( n8086 & n9421 ) ;
  assign n9423 = n9421 | n9422 ;
  assign n9424 = ( ~n6728 & n8088 ) | ( ~n6728 & n9421 ) | ( n8088 & n9421 ) ;
  assign n9425 = n9420 ^ x29 ^ 1'b0 ;
  assign n9426 = n9423 | n9424 ;
  assign n9427 = n7340 & ~n9413 ;
  assign n9428 = n9410 | n9427 ;
  assign n9429 = ( ~n8928 & n9030 ) | ( ~n8928 & n9425 ) | ( n9030 & n9425 ) ;
  assign n9430 = n9425 ^ n9030 ^ n8928 ;
  assign n9431 = n9428 ^ x20 ^ 1'b0 ;
  assign n9432 = n8089 & ~n9413 ;
  assign n9433 = ( n9048 & ~n9144 ) | ( n9048 & n9431 ) | ( ~n9144 & n9431 ) ;
  assign n9434 = n9431 ^ n9144 ^ n9048 ;
  assign n9435 = n6371 & n7486 ;
  assign n9436 = n9426 | n9432 ;
  assign n9437 = n9436 ^ x2 ^ 1'b0 ;
  assign n9438 = ( n6596 & n7493 ) | ( n6596 & n9435 ) | ( n7493 & n9435 ) ;
  assign n9439 = ( ~n6728 & n7485 ) | ( ~n6728 & n9435 ) | ( n7485 & n9435 ) ;
  assign n9440 = ( n9191 & n9276 ) | ( n9191 & n9437 ) | ( n9276 & n9437 ) ;
  assign n9441 = n9435 | n9438 ;
  assign n9442 = n9439 | n9441 ;
  assign n9443 = n7487 & ~n9413 ;
  assign n9444 = n9442 | n9443 ;
  assign n9445 = n9444 ^ x17 ^ 1'b0 ;
  assign n9446 = ( n9045 & n9185 ) | ( n9045 & n9445 ) | ( n9185 & n9445 ) ;
  assign n9447 = n9445 ^ n9185 ^ n9045 ;
  assign n9448 = n6371 & n8033 ;
  assign n9449 = ( n6596 & n8037 ) | ( n6596 & n9448 ) | ( n8037 & n9448 ) ;
  assign n9450 = n9448 | n9449 ;
  assign n9451 = ( ~n6728 & n8029 ) | ( ~n6728 & n9448 ) | ( n8029 & n9448 ) ;
  assign n9452 = n9450 | n9451 ;
  assign n9453 = n8034 & ~n9413 ;
  assign n9454 = n9452 | n9453 ;
  assign n9455 = n9454 ^ x5 ^ 1'b0 ;
  assign n9456 = ( n9139 & n9396 ) | ( n9139 & n9455 ) | ( n9396 & n9455 ) ;
  assign n9457 = n9455 ^ n9396 ^ n9139 ;
  assign n9458 = n6371 & n6907 ;
  assign n9459 = ( n6596 & n6906 ) | ( n6596 & n9458 ) | ( n6906 & n9458 ) ;
  assign n9460 = n9458 | n9459 ;
  assign n9461 = ( ~n6728 & n6901 ) | ( ~n6728 & n9458 ) | ( n6901 & n9458 ) ;
  assign n9462 = n9460 | n9461 ;
  assign n9463 = n6918 & ~n9413 ;
  assign n9464 = n9462 & ~n9463 ;
  assign n9465 = n9464 ^ n9463 ^ x29 ;
  assign n9466 = n6371 & n7929 ;
  assign n9467 = ( n6596 & n7943 ) | ( n6596 & n9466 ) | ( n7943 & n9466 ) ;
  assign n9468 = n9466 | n9467 ;
  assign n9469 = ( ~n6728 & n7932 ) | ( ~n6728 & n9466 ) | ( n7932 & n9466 ) ;
  assign n9470 = n9468 | n9469 ;
  assign n9471 = n7930 & ~n9413 ;
  assign n9472 = n9470 | n9471 ;
  assign n9473 = n9472 ^ x8 ^ 1'b0 ;
  assign n9474 = ( n9159 & n9285 ) | ( n9159 & n9473 ) | ( n9285 & n9473 ) ;
  assign n9475 = n9473 ^ n9285 ^ n9159 ;
  assign n9476 = n6371 & n7667 ;
  assign n9477 = ( n6596 & n7674 ) | ( n6596 & n9476 ) | ( n7674 & n9476 ) ;
  assign n9478 = n9476 | n9477 ;
  assign n9479 = ( ~n6728 & n7669 ) | ( ~n6728 & n9476 ) | ( n7669 & n9476 ) ;
  assign n9480 = n9478 | n9479 ;
  assign n9481 = ( n7666 & ~n9413 ) | ( n7666 & n9480 ) | ( ~n9413 & n9480 ) ;
  assign n9482 = n9480 | n9481 ;
  assign n9483 = ( n9031 & n9209 ) | ( n9031 & n9465 ) | ( n9209 & n9465 ) ;
  assign n9484 = n9465 ^ n9209 ^ n9031 ;
  assign n9485 = n6371 & n7037 ;
  assign n9486 = ( n6596 & n7052 ) | ( n6596 & n9485 ) | ( n7052 & n9485 ) ;
  assign n9487 = n9485 | n9486 ;
  assign n9488 = ( ~n6728 & n7036 ) | ( ~n6728 & n9485 ) | ( n7036 & n9485 ) ;
  assign n9489 = n9487 | n9488 ;
  assign n9490 = n7035 & ~n9413 ;
  assign n9491 = n9489 | n9490 ;
  assign n9492 = n9491 ^ x26 ^ 1'b0 ;
  assign n9493 = n9492 ^ n8958 ^ n8908 ;
  assign n9494 = ( n8908 & n8958 ) | ( n8908 & n9492 ) | ( n8958 & n9492 ) ;
  assign n9495 = n6371 & n7834 ;
  assign n9496 = ( n6596 & n7833 ) | ( n6596 & n9495 ) | ( n7833 & n9495 ) ;
  assign n9497 = n9495 | n9496 ;
  assign n9498 = ( ~n6728 & n7829 ) | ( ~n6728 & n9495 ) | ( n7829 & n9495 ) ;
  assign n9499 = n9497 | n9498 ;
  assign n9500 = n9482 ^ x14 ^ 1'b0 ;
  assign n9501 = n9500 ^ n9355 ^ n9120 ;
  assign n9502 = ( n9120 & n9355 ) | ( n9120 & n9500 ) | ( n9355 & n9500 ) ;
  assign n9503 = ~n6728 & n6791 ;
  assign n9504 = ( n6371 & n6788 ) | ( n6371 & n9503 ) | ( n6788 & n9503 ) ;
  assign n9505 = n9503 | n9504 ;
  assign n9506 = ( n6596 & n6790 ) | ( n6596 & n9503 ) | ( n6790 & n9503 ) ;
  assign n9507 = n9505 | n9506 ;
  assign n9508 = n7838 & ~n9413 ;
  assign n9509 = n9499 | n9508 ;
  assign n9510 = n6596 & ~n6788 ;
  assign n9511 = ( n6596 & n9376 ) | ( n6596 & ~n9510 ) | ( n9376 & ~n9510 ) ;
  assign n9512 = n6789 & ~n9413 ;
  assign n9513 = n9509 ^ x11 ^ 1'b0 ;
  assign n9514 = n7196 & ~n9413 ;
  assign n9515 = n9507 | n9512 ;
  assign n9516 = n6371 & n7188 ;
  assign n9517 = ( n6596 & n7190 ) | ( n6596 & n9516 ) | ( n7190 & n9516 ) ;
  assign n9518 = n9516 | n9517 ;
  assign n9519 = ( ~n6728 & n7192 ) | ( ~n6728 & n9516 ) | ( n7192 & n9516 ) ;
  assign n9520 = n9518 | n9519 ;
  assign n9521 = ( ~n9155 & n9314 ) | ( ~n9155 & n9513 ) | ( n9314 & n9513 ) ;
  assign n9522 = n9513 ^ n9314 ^ n9155 ;
  assign n9523 = n9514 | n9520 ;
  assign n9524 = n9523 ^ x23 ^ 1'b0 ;
  assign n9525 = n9524 ^ n9196 ^ n9090 ;
  assign n9526 = ( n9090 & n9196 ) | ( n9090 & n9524 ) | ( n9196 & n9524 ) ;
  assign n9527 = n6524 & n8033 ;
  assign n9528 = ( n6371 & n8029 ) | ( n6371 & n9527 ) | ( n8029 & n9527 ) ;
  assign n9529 = n9527 | n9528 ;
  assign n9530 = ( n6371 & ~n6728 ) | ( n6371 & n9387 ) | ( ~n6728 & n9387 ) ;
  assign n9531 = ( ~n6728 & n8037 ) | ( ~n6728 & n9527 ) | ( n8037 & n9527 ) ;
  assign n9532 = n9373 ^ x29 ^ 1'b0 ;
  assign n9533 = n9529 | n9531 ;
  assign n9534 = n9530 ^ n6524 ^ n6371 ;
  assign n9535 = n8034 & n9534 ;
  assign n9536 = n9533 | n9535 ;
  assign n9537 = n9536 ^ x5 ^ 1'b0 ;
  assign n9538 = ( n9236 & n9456 ) | ( n9236 & n9537 ) | ( n9456 & n9537 ) ;
  assign n9539 = n9537 ^ n9456 ^ n9236 ;
  assign n9540 = n6524 & n7337 ;
  assign n9541 = ( n6371 & n7339 ) | ( n6371 & n9540 ) | ( n7339 & n9540 ) ;
  assign n9542 = n9540 | n9541 ;
  assign n9543 = ( ~n6728 & n7338 ) | ( ~n6728 & n9540 ) | ( n7338 & n9540 ) ;
  assign n9544 = n9542 | n9543 ;
  assign n9545 = n7340 & n9534 ;
  assign n9546 = n9544 | n9545 ;
  assign n9547 = n9546 ^ x20 ^ 1'b0 ;
  assign n9548 = ( n9131 & n9228 ) | ( n9131 & n9547 ) | ( n9228 & n9547 ) ;
  assign n9549 = n9547 ^ n9228 ^ n9131 ;
  assign n9550 = n6524 & n8090 ;
  assign n9551 = ( n6371 & n8088 ) | ( n6371 & n9550 ) | ( n8088 & n9550 ) ;
  assign n9552 = n9550 | n9551 ;
  assign n9553 = ( ~n6728 & n8086 ) | ( ~n6728 & n9550 ) | ( n8086 & n9550 ) ;
  assign n9554 = n9552 | n9553 ;
  assign n9555 = n8089 & n9534 ;
  assign n9556 = n9554 | n9555 ;
  assign n9557 = n9556 ^ x2 ^ 1'b0 ;
  assign n9558 = ( n9259 & n9440 ) | ( n9259 & n9557 ) | ( n9440 & n9557 ) ;
  assign n9559 = n6524 & n7667 ;
  assign n9560 = ( n6371 & n7669 ) | ( n6371 & n9559 ) | ( n7669 & n9559 ) ;
  assign n9561 = n9559 | n9560 ;
  assign n9562 = ( ~n6728 & n7674 ) | ( ~n6728 & n9559 ) | ( n7674 & n9559 ) ;
  assign n9563 = n9561 | n9562 ;
  assign n9564 = ( n7666 & n9534 ) | ( n7666 & n9563 ) | ( n9534 & n9563 ) ;
  assign n9565 = n9563 | n9564 ;
  assign n9566 = n9565 ^ x14 ^ 1'b0 ;
  assign n9567 = n9566 ^ n9502 ^ n9335 ;
  assign n9568 = ( n9335 & n9502 ) | ( n9335 & n9566 ) | ( n9502 & n9566 ) ;
  assign n9569 = n6524 & n7486 ;
  assign n9570 = ( n6371 & n7485 ) | ( n6371 & n9569 ) | ( n7485 & n9569 ) ;
  assign n9571 = n9569 | n9570 ;
  assign n9572 = ( ~n6728 & n7493 ) | ( ~n6728 & n9569 ) | ( n7493 & n9569 ) ;
  assign n9573 = n9571 | n9572 ;
  assign n9574 = n7487 & n9534 ;
  assign n9575 = n9573 | n9574 ;
  assign n9576 = n9575 ^ x17 ^ 1'b0 ;
  assign n9577 = n9576 ^ n9294 ^ n9184 ;
  assign n9578 = ( n9184 & ~n9294 ) | ( n9184 & n9576 ) | ( ~n9294 & n9576 ) ;
  assign n9579 = n6524 & n7037 ;
  assign n9580 = ( n6371 & n7036 ) | ( n6371 & n9579 ) | ( n7036 & n9579 ) ;
  assign n9581 = n9579 | n9580 ;
  assign n9582 = ( ~n6728 & n7052 ) | ( ~n6728 & n9579 ) | ( n7052 & n9579 ) ;
  assign n9583 = n9581 | n9582 ;
  assign n9584 = n7035 & n9534 ;
  assign n9585 = n9583 | n9584 ;
  assign n9586 = n9585 ^ x26 ^ 1'b0 ;
  assign n9587 = ( n8929 & n9532 ) | ( n8929 & n9586 ) | ( n9532 & n9586 ) ;
  assign n9588 = n9586 ^ n9532 ^ n8929 ;
  assign n9589 = n6524 & n7929 ;
  assign n9590 = ( n6371 & n7932 ) | ( n6371 & n9589 ) | ( n7932 & n9589 ) ;
  assign n9591 = n9589 | n9590 ;
  assign n9592 = ( ~n6728 & n7943 ) | ( ~n6728 & n9589 ) | ( n7943 & n9589 ) ;
  assign n9593 = n9591 | n9592 ;
  assign n9594 = ( n7930 & n9534 ) | ( n7930 & n9593 ) | ( n9534 & n9593 ) ;
  assign n9595 = n9593 | n9594 ;
  assign n9596 = n9595 ^ x8 ^ 1'b0 ;
  assign n9597 = ( n9304 & n9474 ) | ( n9304 & n9596 ) | ( n9474 & n9596 ) ;
  assign n9598 = n9596 ^ n9474 ^ n9304 ;
  assign n9599 = n6524 & n7188 ;
  assign n9600 = ( n6371 & n7192 ) | ( n6371 & n9599 ) | ( n7192 & n9599 ) ;
  assign n9601 = n9599 | n9600 ;
  assign n9602 = ( ~n6728 & n7190 ) | ( ~n6728 & n9599 ) | ( n7190 & n9599 ) ;
  assign n9603 = n9601 | n9602 ;
  assign n9604 = n7196 & n9534 ;
  assign n9605 = n9603 | n9604 ;
  assign n9606 = n9605 ^ x23 ^ 1'b0 ;
  assign n9607 = ( n9197 & n9244 ) | ( n9197 & n9606 ) | ( n9244 & n9606 ) ;
  assign n9608 = n9606 ^ n9244 ^ n9197 ;
  assign n9609 = n6524 & n8088 ;
  assign n9610 = n6524 & n6906 ;
  assign n9611 = ( n6371 & n6524 ) | ( n6371 & n9530 ) | ( n6524 & n9530 ) ;
  assign n9612 = ( ~n6741 & n8090 ) | ( ~n6741 & n9609 ) | ( n8090 & n9609 ) ;
  assign n9613 = ( n6371 & n8086 ) | ( n6371 & n9609 ) | ( n8086 & n9609 ) ;
  assign n9614 = n9609 | n9613 ;
  assign n9615 = n9611 ^ n6741 ^ n6524 ;
  assign n9616 = n9612 | n9614 ;
  assign n9617 = ( n6524 & ~n6741 ) | ( n6524 & n9611 ) | ( ~n6741 & n9611 ) ;
  assign n9618 = ( n8089 & ~n9615 ) | ( n8089 & n9616 ) | ( ~n9615 & n9616 ) ;
  assign n9619 = n9616 | n9618 ;
  assign n9620 = n9619 ^ x2 ^ 1'b0 ;
  assign n9621 = ( ~n6741 & n6901 ) | ( ~n6741 & n9610 ) | ( n6901 & n9610 ) ;
  assign n9622 = ( n9398 & n9558 ) | ( n9398 & n9620 ) | ( n9558 & n9620 ) ;
  assign n9623 = ( ~n6746 & n6907 ) | ( ~n6746 & n9610 ) | ( n6907 & n9610 ) ;
  assign n9624 = n9610 | n9621 ;
  assign n9625 = n9623 | n9624 ;
  assign n9626 = n6524 & n7834 ;
  assign n9627 = ( ~n6728 & n7833 ) | ( ~n6728 & n9626 ) | ( n7833 & n9626 ) ;
  assign n9628 = ( n6371 & n7829 ) | ( n6371 & n9626 ) | ( n7829 & n9626 ) ;
  assign n9629 = n9626 | n9628 ;
  assign n9630 = n9627 | n9629 ;
  assign n9631 = n6524 & n8029 ;
  assign n9632 = ( n6371 & n8037 ) | ( n6371 & n9631 ) | ( n8037 & n9631 ) ;
  assign n9633 = n9631 | n9632 ;
  assign n9634 = ( ~n6741 & n8033 ) | ( ~n6741 & n9631 ) | ( n8033 & n9631 ) ;
  assign n9635 = n9633 | n9634 ;
  assign n9636 = ( n8034 & ~n9615 ) | ( n8034 & n9635 ) | ( ~n9615 & n9635 ) ;
  assign n9637 = n9635 | n9636 ;
  assign n9638 = n9637 ^ x5 ^ 1'b0 ;
  assign n9639 = ( n9286 & n9538 ) | ( n9286 & n9638 ) | ( n9538 & n9638 ) ;
  assign n9640 = n9638 ^ n9538 ^ n9286 ;
  assign n9641 = n9617 ^ n6746 ^ n6741 ;
  assign n9642 = ( n6918 & n9625 ) | ( n6918 & n9641 ) | ( n9625 & n9641 ) ;
  assign n9643 = n9625 | n9642 ;
  assign n9644 = n9643 ^ x29 ^ 1'b0 ;
  assign n9645 = ( n6701 & n9232 ) | ( n6701 & ~n9515 ) | ( n9232 & ~n9515 ) ;
  assign n9646 = ( ~n6701 & n9515 ) | ( ~n6701 & n9645 ) | ( n9515 & n9645 ) ;
  assign n9647 = ( ~n9232 & n9645 ) | ( ~n9232 & n9646 ) | ( n9645 & n9646 ) ;
  assign n9648 = n9647 ^ n9644 ^ n9363 ;
  assign n9649 = ( n9363 & n9644 ) | ( n9363 & n9647 ) | ( n9644 & n9647 ) ;
  assign n9650 = n7838 & n9534 ;
  assign n9651 = n6524 & n8086 ;
  assign n9652 = n9630 | n9650 ;
  assign n9653 = ( ~n6741 & n8088 ) | ( ~n6741 & n9651 ) | ( n8088 & n9651 ) ;
  assign n9654 = n9651 | n9653 ;
  assign n9655 = ( ~n6746 & n8090 ) | ( ~n6746 & n9651 ) | ( n8090 & n9651 ) ;
  assign n9656 = n9654 | n9655 ;
  assign n9657 = ( n8089 & n9641 ) | ( n8089 & n9656 ) | ( n9641 & n9656 ) ;
  assign n9658 = n9656 | n9657 ;
  assign n9659 = n9652 ^ x11 ^ 1'b0 ;
  assign n9660 = n9658 ^ x2 ^ 1'b0 ;
  assign n9661 = n6524 & n6907 ;
  assign n9662 = ( n9457 & n9622 ) | ( n9457 & n9660 ) | ( n9622 & n9660 ) ;
  assign n9663 = n6789 & ~n9534 ;
  assign n9664 = ( n6371 & n6901 ) | ( n6371 & n9661 ) | ( n6901 & n9661 ) ;
  assign n9665 = n9661 | n9664 ;
  assign n9666 = n6918 & n9534 ;
  assign n9667 = ( ~n6728 & n6906 ) | ( ~n6728 & n9661 ) | ( n6906 & n9661 ) ;
  assign n9668 = n9665 | n9667 ;
  assign n9669 = n9666 | n9668 ;
  assign n9670 = ( n9344 & n9521 ) | ( n9344 & n9659 ) | ( n9521 & n9659 ) ;
  assign n9671 = n6371 & n6791 ;
  assign n9672 = n9669 ^ x29 ^ 1'b0 ;
  assign n9673 = n9659 ^ n9521 ^ n9344 ;
  assign n9674 = n9672 ^ n9511 ^ n9223 ;
  assign n9675 = ( ~n9223 & n9511 ) | ( ~n9223 & n9672 ) | ( n9511 & n9672 ) ;
  assign n9676 = ( n6524 & n6788 ) | ( n6524 & n9671 ) | ( n6788 & n9671 ) ;
  assign n9677 = ( ~n6728 & n6790 ) | ( ~n6728 & n9671 ) | ( n6790 & n9671 ) ;
  assign n9678 = n9671 | n9676 ;
  assign n9679 = n9677 | n9678 ;
  assign n9680 = ( n6789 & ~n9663 ) | ( n6789 & n9679 ) | ( ~n9663 & n9679 ) ;
  assign n9681 = n9680 ^ n6701 ^ n6490 ;
  assign n9682 = ( n6490 & n6701 ) | ( n6490 & ~n9680 ) | ( n6701 & ~n9680 ) ;
  assign n9683 = n9681 ^ n9649 ^ n9645 ;
  assign n9684 = ( ~n9645 & n9649 ) | ( ~n9645 & n9681 ) | ( n9649 & n9681 ) ;
  assign n9685 = n6524 & n7669 ;
  assign n9686 = ( n6371 & n7674 ) | ( n6371 & n9685 ) | ( n7674 & n9685 ) ;
  assign n9687 = n9685 | n9686 ;
  assign n9688 = ( ~n6741 & n7667 ) | ( ~n6741 & n9685 ) | ( n7667 & n9685 ) ;
  assign n9689 = n9687 | n9688 ;
  assign n9690 = n7666 & ~n9615 ;
  assign n9691 = n9689 | n9690 ;
  assign n9692 = n9691 ^ x14 ^ 1'b0 ;
  assign n9693 = n9692 ^ n9411 ^ n9334 ;
  assign n9694 = ( n9334 & n9411 ) | ( n9334 & n9692 ) | ( n9411 & n9692 ) ;
  assign n9695 = n6524 & n7192 ;
  assign n9696 = ( n6371 & n7190 ) | ( n6371 & n9695 ) | ( n7190 & n9695 ) ;
  assign n9697 = n9695 | n9696 ;
  assign n9698 = ( ~n6741 & n7188 ) | ( ~n6741 & n9695 ) | ( n7188 & n9695 ) ;
  assign n9699 = n9697 | n9698 ;
  assign n9700 = n7196 & ~n9615 ;
  assign n9701 = n9699 | n9700 ;
  assign n9702 = n9701 ^ x23 ^ 1'b0 ;
  assign n9703 = ( n9266 & n9607 ) | ( n9266 & n9702 ) | ( n9607 & n9702 ) ;
  assign n9704 = n9702 ^ n9607 ^ n9266 ;
  assign n9705 = n6701 ^ n6554 ^ x20 ;
  assign n9706 = ( ~x20 & n6554 ) | ( ~x20 & n6701 ) | ( n6554 & n6701 ) ;
  assign n9707 = n6524 & n7829 ;
  assign n9708 = ( n6371 & n7833 ) | ( n6371 & n9707 ) | ( n7833 & n9707 ) ;
  assign n9709 = n9707 | n9708 ;
  assign n9710 = ( ~n6741 & n7834 ) | ( ~n6741 & n9707 ) | ( n7834 & n9707 ) ;
  assign n9711 = n9709 | n9710 ;
  assign n9712 = n7838 & ~n9615 ;
  assign n9713 = n9711 | n9712 ;
  assign n9714 = n9713 ^ x11 ^ 1'b0 ;
  assign n9715 = ( ~n9354 & n9670 ) | ( ~n9354 & n9714 ) | ( n9670 & n9714 ) ;
  assign n9716 = n9714 ^ n9670 ^ n9354 ;
  assign n9717 = n6524 & n7339 ;
  assign n9718 = ( n6371 & n7338 ) | ( n6371 & n9717 ) | ( n7338 & n9717 ) ;
  assign n9719 = n9717 | n9718 ;
  assign n9720 = ( ~n6741 & n7337 ) | ( ~n6741 & n9717 ) | ( n7337 & n9717 ) ;
  assign n9721 = n9719 | n9720 ;
  assign n9722 = ( n7340 & ~n9615 ) | ( n7340 & n9721 ) | ( ~n9615 & n9721 ) ;
  assign n9723 = n9721 | n9722 ;
  assign n9724 = n9723 ^ x20 ^ 1'b0 ;
  assign n9725 = n9724 ^ n9548 ^ n9394 ;
  assign n9726 = ( n9394 & n9548 ) | ( n9394 & n9724 ) | ( n9548 & n9724 ) ;
  assign n9727 = n6524 & n7932 ;
  assign n9728 = ( n6371 & n7943 ) | ( n6371 & n9727 ) | ( n7943 & n9727 ) ;
  assign n9729 = n9727 | n9728 ;
  assign n9730 = ( ~n6741 & n7929 ) | ( ~n6741 & n9727 ) | ( n7929 & n9727 ) ;
  assign n9731 = n9729 | n9730 ;
  assign n9732 = ( n7930 & ~n9615 ) | ( n7930 & n9731 ) | ( ~n9615 & n9731 ) ;
  assign n9733 = n9731 | n9732 ;
  assign n9734 = n9733 ^ x8 ^ 1'b0 ;
  assign n9735 = n9734 ^ n9597 ^ n9315 ;
  assign n9736 = ( ~n9315 & n9597 ) | ( ~n9315 & n9734 ) | ( n9597 & n9734 ) ;
  assign n9737 = n6524 & n7036 ;
  assign n9738 = ( n6371 & n7052 ) | ( n6371 & n9737 ) | ( n7052 & n9737 ) ;
  assign n9739 = n9737 | n9738 ;
  assign n9740 = ( ~n6741 & n7037 ) | ( ~n6741 & n9737 ) | ( n7037 & n9737 ) ;
  assign n9741 = n9739 | n9740 ;
  assign n9742 = n7035 & ~n9615 ;
  assign n9743 = n9741 & ~n9742 ;
  assign n9744 = n9743 ^ n9742 ^ x26 ;
  assign n9745 = ( ~n9430 & n9587 ) | ( ~n9430 & n9744 ) | ( n9587 & n9744 ) ;
  assign n9746 = n9744 ^ n9587 ^ n9430 ;
  assign n9747 = n6524 & n6901 ;
  assign n9748 = ( n6371 & n6906 ) | ( n6371 & n9747 ) | ( n6906 & n9747 ) ;
  assign n9749 = n9747 | n9748 ;
  assign n9750 = ( ~n6741 & n6907 ) | ( ~n6741 & n9747 ) | ( n6907 & n9747 ) ;
  assign n9751 = n9749 | n9750 ;
  assign n9752 = n6918 & ~n9615 ;
  assign n9753 = n9751 | n9752 ;
  assign n9754 = n9753 ^ x29 ^ 1'b0 ;
  assign n9755 = ( n9364 & n9675 ) | ( n9364 & n9754 ) | ( n9675 & n9754 ) ;
  assign n9756 = n9754 ^ n9675 ^ n9364 ;
  assign n9757 = n6524 & n7485 ;
  assign n9758 = ( n6371 & n7493 ) | ( n6371 & n9757 ) | ( n7493 & n9757 ) ;
  assign n9759 = n9757 | n9758 ;
  assign n9760 = ( ~n6741 & n7486 ) | ( ~n6741 & n9757 ) | ( n7486 & n9757 ) ;
  assign n9761 = n9759 | n9760 ;
  assign n9762 = n7487 & ~n9615 ;
  assign n9763 = n9761 | n9762 ;
  assign n9764 = n9763 ^ x17 ^ 1'b0 ;
  assign n9765 = ( n9325 & n9578 ) | ( n9325 & n9764 ) | ( n9578 & n9764 ) ;
  assign n9766 = n6789 & ~n9615 ;
  assign n9767 = n9764 ^ n9578 ^ n9325 ;
  assign n9768 = n6524 & n6791 ;
  assign n9769 = ( n6371 & n6790 ) | ( n6371 & n9768 ) | ( n6790 & n9768 ) ;
  assign n9770 = n9768 | n9769 ;
  assign n9771 = ( ~n6741 & n6788 ) | ( ~n6741 & n9768 ) | ( n6788 & n9768 ) ;
  assign n9772 = n9770 | n9771 ;
  assign n9773 = n9766 | n9772 ;
  assign n9774 = ( n9682 & n9705 ) | ( n9682 & ~n9773 ) | ( n9705 & ~n9773 ) ;
  assign n9775 = n9773 ^ n9705 ^ n9682 ;
  assign n9776 = n6524 & n7943 ;
  assign n9777 = ( ~n6741 & n7932 ) | ( ~n6741 & n9776 ) | ( n7932 & n9776 ) ;
  assign n9778 = n9776 | n9777 ;
  assign n9779 = ( ~n6746 & n7929 ) | ( ~n6746 & n9776 ) | ( n7929 & n9776 ) ;
  assign n9780 = n9778 | n9779 ;
  assign n9781 = ( n7930 & n9641 ) | ( n7930 & n9780 ) | ( n9641 & n9780 ) ;
  assign n9782 = n9780 | n9781 ;
  assign n9783 = n9782 ^ x8 ^ 1'b0 ;
  assign n9784 = n9783 ^ n9736 ^ n9522 ;
  assign n9785 = ( ~n9522 & n9736 ) | ( ~n9522 & n9783 ) | ( n9736 & n9783 ) ;
  assign n9786 = n6524 & n7493 ;
  assign n9787 = ( ~n6741 & n7485 ) | ( ~n6741 & n9786 ) | ( n7485 & n9786 ) ;
  assign n9788 = n9786 | n9787 ;
  assign n9789 = ( ~n6746 & n7486 ) | ( ~n6746 & n9786 ) | ( n7486 & n9786 ) ;
  assign n9790 = n9788 | n9789 ;
  assign n9791 = n7487 & n9641 ;
  assign n9792 = n9790 | n9791 ;
  assign n9793 = n9792 ^ x17 ^ 1'b0 ;
  assign n9794 = n9793 ^ n9434 ^ n9324 ;
  assign n9795 = ( n9324 & ~n9434 ) | ( n9324 & n9793 ) | ( ~n9434 & n9793 ) ;
  assign n9796 = n6524 & n7833 ;
  assign n9797 = ( ~n6741 & n7829 ) | ( ~n6741 & n9796 ) | ( n7829 & n9796 ) ;
  assign n9798 = n9796 | n9797 ;
  assign n9799 = ( ~n6746 & n7834 ) | ( ~n6746 & n9796 ) | ( n7834 & n9796 ) ;
  assign n9800 = n9798 | n9799 ;
  assign n9801 = n7838 & n9641 ;
  assign n9802 = n9800 | n9801 ;
  assign n9803 = n9802 ^ x11 ^ 1'b0 ;
  assign n9804 = ( n9501 & n9715 ) | ( n9501 & n9803 ) | ( n9715 & n9803 ) ;
  assign n9805 = n9803 ^ n9715 ^ n9501 ;
  assign n9806 = n6524 & n7674 ;
  assign n9807 = ( ~n6741 & n7669 ) | ( ~n6741 & n9806 ) | ( n7669 & n9806 ) ;
  assign n9808 = n9806 | n9807 ;
  assign n9809 = ( ~n6746 & n7667 ) | ( ~n6746 & n9806 ) | ( n7667 & n9806 ) ;
  assign n9810 = n9808 | n9809 ;
  assign n9811 = n7666 & n9641 ;
  assign n9812 = n9810 | n9811 ;
  assign n9813 = n9812 ^ x14 ^ 1'b0 ;
  assign n9814 = ( n9412 & n9447 ) | ( n9412 & n9813 ) | ( n9447 & n9813 ) ;
  assign n9815 = n9813 ^ n9447 ^ n9412 ;
  assign n9816 = n6524 & n7190 ;
  assign n9817 = ( ~n6746 & n7188 ) | ( ~n6746 & n9816 ) | ( n7188 & n9816 ) ;
  assign n9818 = n9816 | n9817 ;
  assign n9819 = ( ~n6741 & n7192 ) | ( ~n6741 & n9816 ) | ( n7192 & n9816 ) ;
  assign n9820 = n9818 | n9819 ;
  assign n9821 = n7196 & n9641 ;
  assign n9822 = n9820 | n9821 ;
  assign n9823 = n9822 ^ x23 ^ 1'b0 ;
  assign n9824 = ( n9265 & n9493 ) | ( n9265 & n9823 ) | ( n9493 & n9823 ) ;
  assign n9825 = n9823 ^ n9493 ^ n9265 ;
  assign n9826 = n6524 & n8037 ;
  assign n9827 = ( ~n6741 & n8029 ) | ( ~n6741 & n9826 ) | ( n8029 & n9826 ) ;
  assign n9828 = n9826 | n9827 ;
  assign n9829 = ( ~n6746 & n8033 ) | ( ~n6746 & n9826 ) | ( n8033 & n9826 ) ;
  assign n9830 = n9828 | n9829 ;
  assign n9831 = ( n8034 & n9641 ) | ( n8034 & n9830 ) | ( n9641 & n9830 ) ;
  assign n9832 = n9830 | n9831 ;
  assign n9833 = n9832 ^ x5 ^ 1'b0 ;
  assign n9834 = ( n9475 & n9639 ) | ( n9475 & n9833 ) | ( n9639 & n9833 ) ;
  assign n9835 = n9833 ^ n9639 ^ n9475 ;
  assign n9836 = n6524 & n7338 ;
  assign n9837 = ( ~n6741 & n7339 ) | ( ~n6741 & n9836 ) | ( n7339 & n9836 ) ;
  assign n9838 = n9836 | n9837 ;
  assign n9839 = ( ~n6746 & n7337 ) | ( ~n6746 & n9836 ) | ( n7337 & n9836 ) ;
  assign n9840 = n9838 | n9839 ;
  assign n9841 = n7340 & n9641 ;
  assign n9842 = n9840 | n9841 ;
  assign n9843 = n9842 ^ x20 ^ 1'b0 ;
  assign n9844 = ( n9395 & n9525 ) | ( n9395 & n9843 ) | ( n9525 & n9843 ) ;
  assign n9845 = n9843 ^ n9525 ^ n9395 ;
  assign n9846 = ~n6741 & n6791 ;
  assign n9847 = ( n6524 & n6790 ) | ( n6524 & n9846 ) | ( n6790 & n9846 ) ;
  assign n9848 = n6524 & n7052 ;
  assign n9849 = n9846 | n9847 ;
  assign n9850 = ( ~n6746 & n6788 ) | ( ~n6746 & n9846 ) | ( n6788 & n9846 ) ;
  assign n9851 = n9849 | n9850 ;
  assign n9852 = ( ~n6746 & n7037 ) | ( ~n6746 & n9848 ) | ( n7037 & n9848 ) ;
  assign n9853 = n9848 | n9852 ;
  assign n9854 = ( ~n6741 & n7036 ) | ( ~n6741 & n9848 ) | ( n7036 & n9848 ) ;
  assign n9855 = n9853 | n9854 ;
  assign n9856 = n7035 & n9641 ;
  assign n9857 = n9855 | n9856 ;
  assign n9858 = n6789 & ~n9641 ;
  assign n9859 = ( n6789 & n9851 ) | ( n6789 & ~n9858 ) | ( n9851 & ~n9858 ) ;
  assign n9860 = n9857 ^ x26 ^ 1'b0 ;
  assign n9861 = n9860 ^ n9484 ^ n9429 ;
  assign n9862 = ( n9429 & n9484 ) | ( n9429 & n9860 ) | ( n9484 & n9860 ) ;
  assign n9863 = n6747 & n8090 ;
  assign n9864 = ( n6741 & n6746 ) | ( n6741 & ~n9617 ) | ( n6746 & ~n9617 ) ;
  assign n9865 = n9864 ^ n6747 ^ n6746 ;
  assign n9866 = ( ~n6741 & n8086 ) | ( ~n6741 & n9863 ) | ( n8086 & n9863 ) ;
  assign n9867 = ( n6746 & ~n6747 ) | ( n6746 & n9864 ) | ( ~n6747 & n9864 ) ;
  assign n9868 = n9863 | n9866 ;
  assign n9869 = ( ~n6746 & n8088 ) | ( ~n6746 & n9863 ) | ( n8088 & n9863 ) ;
  assign n9870 = n9868 | n9869 ;
  assign n9871 = ( n8089 & n9865 ) | ( n8089 & n9870 ) | ( n9865 & n9870 ) ;
  assign n9872 = n9870 | n9871 ;
  assign n9873 = n6823 & n7834 ;
  assign n9874 = n9872 ^ x2 ^ 1'b0 ;
  assign n9875 = ( n9539 & n9662 ) | ( n9539 & n9874 ) | ( n9662 & n9874 ) ;
  assign n9876 = ( n6747 & n7829 ) | ( n6747 & n9873 ) | ( n7829 & n9873 ) ;
  assign n9877 = n9867 ^ n6823 ^ n6747 ;
  assign n9878 = n9873 | n9876 ;
  assign n9879 = ( ~n6746 & n7833 ) | ( ~n6746 & n9873 ) | ( n7833 & n9873 ) ;
  assign n9880 = n9878 | n9879 ;
  assign n9881 = n7838 & ~n9877 ;
  assign n9882 = n9880 | n9881 ;
  assign n9883 = n9882 ^ x11 ^ 1'b0 ;
  assign n9884 = n9883 ^ n9693 ^ n9568 ;
  assign n9885 = ( n9568 & n9693 ) | ( n9568 & n9883 ) | ( n9693 & n9883 ) ;
  assign n9886 = n6747 & n7834 ;
  assign n9887 = ( ~n6746 & n7829 ) | ( ~n6746 & n9886 ) | ( n7829 & n9886 ) ;
  assign n9888 = n9886 | n9887 ;
  assign n9889 = ( ~n6741 & n7833 ) | ( ~n6741 & n9886 ) | ( n7833 & n9886 ) ;
  assign n9890 = n9888 | n9889 ;
  assign n9891 = n7838 & n9865 ;
  assign n9892 = n9890 | n9891 ;
  assign n9893 = n9892 ^ x11 ^ 1'b0 ;
  assign n9894 = ( n9567 & n9804 ) | ( n9567 & n9893 ) | ( n9804 & n9893 ) ;
  assign n9895 = n9893 ^ n9804 ^ n9567 ;
  assign n9896 = n6747 & n7337 ;
  assign n9897 = ( ~n6746 & n7339 ) | ( ~n6746 & n9896 ) | ( n7339 & n9896 ) ;
  assign n9898 = n9896 | n9897 ;
  assign n9899 = ( ~n6741 & n7338 ) | ( ~n6741 & n9896 ) | ( n7338 & n9896 ) ;
  assign n9900 = n9898 | n9899 ;
  assign n9901 = n7340 & n9865 ;
  assign n9902 = n9900 | n9901 ;
  assign n9903 = n9902 ^ x20 ^ 1'b0 ;
  assign n9904 = n5913 | n6687 ;
  assign n9905 = n9903 ^ n9608 ^ n9526 ;
  assign n9906 = ( n9526 & n9608 ) | ( n9526 & n9903 ) | ( n9608 & n9903 ) ;
  assign n9907 = n6747 & n7667 ;
  assign n9908 = ( ~n6746 & n7669 ) | ( ~n6746 & n9907 ) | ( n7669 & n9907 ) ;
  assign n9909 = n9907 | n9908 ;
  assign n9910 = ( ~n6741 & n7674 ) | ( ~n6741 & n9907 ) | ( n7674 & n9907 ) ;
  assign n9911 = n9909 | n9910 ;
  assign n9912 = n6035 & ~n6687 ;
  assign n9913 = n7666 & n9865 ;
  assign n9914 = n9911 | n9913 ;
  assign n9915 = n9914 ^ x14 ^ 1'b0 ;
  assign n9916 = n9915 ^ n9577 ^ n9446 ;
  assign n9917 = ( n9446 & ~n9577 ) | ( n9446 & n9915 ) | ( ~n9577 & n9915 ) ;
  assign n9918 = n6747 & n8033 ;
  assign n9919 = ( ~n6746 & n8029 ) | ( ~n6746 & n9918 ) | ( n8029 & n9918 ) ;
  assign n9920 = n9918 | n9919 ;
  assign n9921 = ( ~n6741 & n8037 ) | ( ~n6741 & n9918 ) | ( n8037 & n9918 ) ;
  assign n9922 = n9920 | n9921 ;
  assign n9923 = n8034 & n9865 ;
  assign n9924 = n9922 | n9923 ;
  assign n9925 = n9924 ^ x5 ^ 1'b0 ;
  assign n9926 = ( n9598 & n9834 ) | ( n9598 & n9925 ) | ( n9834 & n9925 ) ;
  assign n9927 = n9925 ^ n9834 ^ n9598 ;
  assign n9928 = n6823 & n8090 ;
  assign n9929 = ( n6747 & n8088 ) | ( n6747 & n9928 ) | ( n8088 & n9928 ) ;
  assign n9930 = n9928 | n9929 ;
  assign n9931 = ( ~n6746 & n8086 ) | ( ~n6746 & n9928 ) | ( n8086 & n9928 ) ;
  assign n9932 = n9930 | n9931 ;
  assign n9933 = n8089 & ~n9877 ;
  assign n9934 = n9932 | n9933 ;
  assign n9935 = n9934 ^ x2 ^ 1'b0 ;
  assign n9936 = ( n9640 & n9875 ) | ( n9640 & n9935 ) | ( n9875 & n9935 ) ;
  assign n9937 = n6823 & n8088 ;
  assign n9938 = ( n6747 & n8086 ) | ( n6747 & n9937 ) | ( n8086 & n9937 ) ;
  assign n9939 = n9937 | n9938 ;
  assign n9940 = ( ~n6752 & n8090 ) | ( ~n6752 & n9937 ) | ( n8090 & n9937 ) ;
  assign n9941 = n9939 | n9940 ;
  assign n9942 = ( n6747 & n6823 ) | ( n6747 & ~n9867 ) | ( n6823 & ~n9867 ) ;
  assign n9943 = n9942 ^ n6823 ^ n6752 ;
  assign n9944 = n8089 & ~n9943 ;
  assign n9945 = n9941 | n9944 ;
  assign n9946 = n9945 ^ x2 ^ 1'b0 ;
  assign n9947 = ( n9835 & n9936 ) | ( n9835 & n9946 ) | ( n9936 & n9946 ) ;
  assign n9948 = n6823 & n8033 ;
  assign n9949 = ( n6747 & n8029 ) | ( n6747 & n9948 ) | ( n8029 & n9948 ) ;
  assign n9950 = n9948 | n9949 ;
  assign n9951 = ( ~n6746 & n8037 ) | ( ~n6746 & n9948 ) | ( n8037 & n9948 ) ;
  assign n9952 = n9950 | n9951 ;
  assign n9953 = n8034 & ~n9877 ;
  assign n9954 = n9952 | n9953 ;
  assign n9955 = n6823 & n8029 ;
  assign n9956 = n9954 ^ x5 ^ 1'b0 ;
  assign n9957 = ( ~n9735 & n9926 ) | ( ~n9735 & n9956 ) | ( n9926 & n9956 ) ;
  assign n9958 = n9956 ^ n9926 ^ n9735 ;
  assign n9959 = ( n6747 & n8037 ) | ( n6747 & n9955 ) | ( n8037 & n9955 ) ;
  assign n9960 = n9955 | n9959 ;
  assign n9961 = ( ~n6752 & n8033 ) | ( ~n6752 & n9955 ) | ( n8033 & n9955 ) ;
  assign n9962 = n9960 | n9961 ;
  assign n9963 = n8034 & ~n9943 ;
  assign n9964 = n9962 | n9963 ;
  assign n9965 = n9964 ^ x5 ^ 1'b0 ;
  assign n9966 = n9965 ^ n9957 ^ n9784 ;
  assign n9967 = ( ~n9784 & n9957 ) | ( ~n9784 & n9965 ) | ( n9957 & n9965 ) ;
  assign n9968 = n6823 & n7669 ;
  assign n9969 = ( n6747 & n7674 ) | ( n6747 & n9968 ) | ( n7674 & n9968 ) ;
  assign n9970 = ( ~n6752 & n7667 ) | ( ~n6752 & n9968 ) | ( n7667 & n9968 ) ;
  assign n9971 = n9968 | n9969 ;
  assign n9972 = n9970 | n9971 ;
  assign n9973 = n7666 & ~n9943 ;
  assign n9974 = n9972 | n9973 ;
  assign n9975 = n6823 & n7486 ;
  assign n9976 = ( n6747 & n7485 ) | ( n6747 & n9975 ) | ( n7485 & n9975 ) ;
  assign n9977 = n9975 | n9976 ;
  assign n9978 = ( ~n6746 & n7493 ) | ( ~n6746 & n9975 ) | ( n7493 & n9975 ) ;
  assign n9979 = n9977 | n9978 ;
  assign n9980 = n7487 & ~n9877 ;
  assign n9981 = n9979 | n9980 ;
  assign n9982 = n9981 ^ x17 ^ 1'b0 ;
  assign n9983 = n9974 ^ x14 ^ 1'b0 ;
  assign n9984 = ( n9765 & ~n9794 ) | ( n9765 & n9983 ) | ( ~n9794 & n9983 ) ;
  assign n9985 = n9983 ^ n9794 ^ n9765 ;
  assign n9986 = n6747 & n7486 ;
  assign n9987 = ( ~n6746 & n7485 ) | ( ~n6746 & n9986 ) | ( n7485 & n9986 ) ;
  assign n9988 = n9986 | n9987 ;
  assign n9989 = ( ~n6741 & n7493 ) | ( ~n6741 & n9986 ) | ( n7493 & n9986 ) ;
  assign n9990 = n9988 | n9989 ;
  assign n9991 = n7487 & n9865 ;
  assign n9992 = n9990 | n9991 ;
  assign n9993 = n9992 ^ x17 ^ 1'b0 ;
  assign n9994 = ( n9433 & n9549 ) | ( n9433 & n9993 ) | ( n9549 & n9993 ) ;
  assign n9995 = n9993 ^ n9549 ^ n9433 ;
  assign n9996 = n9994 ^ n9982 ^ n9725 ;
  assign n9997 = ( n9725 & n9982 ) | ( n9725 & n9994 ) | ( n9982 & n9994 ) ;
  assign n9998 = n6823 & n7667 ;
  assign n9999 = ( ~n6746 & n7674 ) | ( ~n6746 & n9998 ) | ( n7674 & n9998 ) ;
  assign n10000 = ( n6747 & n7669 ) | ( n6747 & n9998 ) | ( n7669 & n9998 ) ;
  assign n10001 = n9998 | n10000 ;
  assign n10002 = n9999 | n10001 ;
  assign n10003 = ( n7666 & ~n9877 ) | ( n7666 & n10002 ) | ( ~n9877 & n10002 ) ;
  assign n10004 = n10002 | n10003 ;
  assign n10005 = n10004 ^ x14 ^ 1'b0 ;
  assign n10006 = ( n9767 & n9917 ) | ( n9767 & n10005 ) | ( n9917 & n10005 ) ;
  assign n10007 = n10005 ^ n9917 ^ n9767 ;
  assign n10008 = n6823 & n8086 ;
  assign n10009 = ( ~n6752 & n8088 ) | ( ~n6752 & n10008 ) | ( n8088 & n10008 ) ;
  assign n10010 = ( n6751 & n8090 ) | ( n6751 & n10008 ) | ( n8090 & n10008 ) ;
  assign n10011 = n10008 | n10010 ;
  assign n10012 = ( ~n6752 & n6823 ) | ( ~n6752 & n9942 ) | ( n6823 & n9942 ) ;
  assign n10013 = n10012 ^ n6752 ^ n6751 ;
  assign n10014 = n10009 | n10011 ;
  assign n10015 = ( n8089 & ~n10013 ) | ( n8089 & n10014 ) | ( ~n10013 & n10014 ) ;
  assign n10016 = n10014 | n10015 ;
  assign n10017 = n10016 ^ x2 ^ 1'b0 ;
  assign n10018 = ( n9927 & n9947 ) | ( n9927 & n10017 ) | ( n9947 & n10017 ) ;
  assign n10019 = n6823 & n7829 ;
  assign n10020 = ( n6747 & n7833 ) | ( n6747 & n10019 ) | ( n7833 & n10019 ) ;
  assign n10021 = n10019 | n10020 ;
  assign n10022 = ( ~n6752 & n7834 ) | ( ~n6752 & n10019 ) | ( n7834 & n10019 ) ;
  assign n10023 = n10021 | n10022 ;
  assign n10024 = n6747 & n7929 ;
  assign n10025 = ( ~n6746 & n7932 ) | ( ~n6746 & n10024 ) | ( n7932 & n10024 ) ;
  assign n10026 = n10024 | n10025 ;
  assign n10027 = ( ~n6741 & n7943 ) | ( ~n6741 & n10024 ) | ( n7943 & n10024 ) ;
  assign n10028 = n10026 | n10027 ;
  assign n10029 = n7838 & ~n9943 ;
  assign n10030 = n10023 | n10029 ;
  assign n10031 = ( n7930 & n9865 ) | ( n7930 & n10028 ) | ( n9865 & n10028 ) ;
  assign n10032 = n10030 ^ x11 ^ 1'b0 ;
  assign n10033 = n10028 | n10031 ;
  assign n10034 = ( n9694 & n9815 ) | ( n9694 & n10032 ) | ( n9815 & n10032 ) ;
  assign n10035 = n10032 ^ n9815 ^ n9694 ;
  assign n10036 = n6823 & n7493 ;
  assign n10037 = ( n6751 & n7486 ) | ( n6751 & n10036 ) | ( n7486 & n10036 ) ;
  assign n10038 = n10036 | n10037 ;
  assign n10039 = n10033 ^ x8 ^ 1'b0 ;
  assign n10040 = ( ~n6752 & n7485 ) | ( ~n6752 & n10036 ) | ( n7485 & n10036 ) ;
  assign n10041 = n10038 | n10040 ;
  assign n10042 = n7487 & ~n10013 ;
  assign n10043 = n10041 | n10042 ;
  assign n10044 = ( n9673 & n9785 ) | ( n9673 & n10039 ) | ( n9785 & n10039 ) ;
  assign n10045 = n10039 ^ n9785 ^ n9673 ;
  assign n10046 = n10043 ^ x17 ^ 1'b0 ;
  assign n10047 = ( n9844 & n9905 ) | ( n9844 & n10046 ) | ( n9905 & n10046 ) ;
  assign n10048 = n10046 ^ n9905 ^ n9844 ;
  assign n10049 = n6823 & n7929 ;
  assign n10050 = ( n6747 & n7932 ) | ( n6747 & n10049 ) | ( n7932 & n10049 ) ;
  assign n10051 = n10049 | n10050 ;
  assign n10052 = ( ~n6746 & n7943 ) | ( ~n6746 & n10049 ) | ( n7943 & n10049 ) ;
  assign n10053 = n10051 | n10052 ;
  assign n10054 = ( n7930 & ~n9877 ) | ( n7930 & n10053 ) | ( ~n9877 & n10053 ) ;
  assign n10055 = n10053 | n10054 ;
  assign n10056 = n10055 ^ x8 ^ 1'b0 ;
  assign n10057 = n6823 & n7932 ;
  assign n10058 = n10056 ^ n10044 ^ n9716 ;
  assign n10059 = ( ~n9716 & n10044 ) | ( ~n9716 & n10056 ) | ( n10044 & n10056 ) ;
  assign n10060 = ( ~n6752 & n7929 ) | ( ~n6752 & n10057 ) | ( n7929 & n10057 ) ;
  assign n10061 = ( n6747 & n7943 ) | ( n6747 & n10057 ) | ( n7943 & n10057 ) ;
  assign n10062 = n10057 | n10061 ;
  assign n10063 = n10060 | n10062 ;
  assign n10064 = ( n7930 & ~n9943 ) | ( n7930 & n10063 ) | ( ~n9943 & n10063 ) ;
  assign n10065 = n10063 | n10064 ;
  assign n10066 = n10065 ^ x8 ^ 1'b0 ;
  assign n10067 = n10066 ^ n10059 ^ n9805 ;
  assign n10068 = ( n9805 & n10059 ) | ( n9805 & n10066 ) | ( n10059 & n10066 ) ;
  assign n10069 = n6823 & n7674 ;
  assign n10070 = ( n6751 & n7667 ) | ( n6751 & n10069 ) | ( n7667 & n10069 ) ;
  assign n10071 = n10069 | n10070 ;
  assign n10072 = ( ~n6752 & n7669 ) | ( ~n6752 & n10069 ) | ( n7669 & n10069 ) ;
  assign n10073 = n10071 | n10072 ;
  assign n10074 = n7666 & ~n10013 ;
  assign n10075 = n10073 | n10074 ;
  assign n10076 = n10075 ^ x14 ^ 1'b0 ;
  assign n10077 = ( n9795 & n9995 ) | ( n9795 & n10076 ) | ( n9995 & n10076 ) ;
  assign n10078 = n10076 ^ n9995 ^ n9795 ;
  assign n10079 = n6823 & n8037 ;
  assign n10080 = ( n6751 & n8033 ) | ( n6751 & n10079 ) | ( n8033 & n10079 ) ;
  assign n10081 = n10079 | n10080 ;
  assign n10082 = ( ~n6752 & n8029 ) | ( ~n6752 & n10079 ) | ( n8029 & n10079 ) ;
  assign n10083 = n10081 | n10082 ;
  assign n10084 = n8034 & ~n10013 ;
  assign n10085 = n10083 | n10084 ;
  assign n10086 = n10085 ^ x5 ^ 1'b0 ;
  assign n10087 = n10086 ^ n10045 ^ n9967 ;
  assign n10088 = ( n9967 & n10045 ) | ( n9967 & n10086 ) | ( n10045 & n10086 ) ;
  assign n10089 = n6823 & n7943 ;
  assign n10090 = ( n6751 & n7929 ) | ( n6751 & n10089 ) | ( n7929 & n10089 ) ;
  assign n10091 = n10089 | n10090 ;
  assign n10092 = ( ~n6752 & n7932 ) | ( ~n6752 & n10089 ) | ( n7932 & n10089 ) ;
  assign n10093 = n10091 | n10092 ;
  assign n10094 = ( n7930 & ~n10013 ) | ( n7930 & n10093 ) | ( ~n10013 & n10093 ) ;
  assign n10095 = n10093 | n10094 ;
  assign n10096 = n10095 ^ x8 ^ 1'b0 ;
  assign n10097 = ( n9895 & n10068 ) | ( n9895 & n10096 ) | ( n10068 & n10096 ) ;
  assign n10098 = n10096 ^ n10068 ^ n9895 ;
  assign n10099 = n6823 & n7337 ;
  assign n10100 = ( n6747 & n7339 ) | ( n6747 & n10099 ) | ( n7339 & n10099 ) ;
  assign n10101 = n10099 | n10100 ;
  assign n10102 = ( ~n6746 & n7338 ) | ( ~n6746 & n10099 ) | ( n7338 & n10099 ) ;
  assign n10103 = n10101 | n10102 ;
  assign n10104 = ( n7340 & ~n9877 ) | ( n7340 & n10103 ) | ( ~n9877 & n10103 ) ;
  assign n10105 = n10103 | n10104 ;
  assign n10106 = n10105 ^ x20 ^ 1'b0 ;
  assign n10107 = ( n6751 & ~n6752 ) | ( n6751 & n10012 ) | ( ~n6752 & n10012 ) ;
  assign n10108 = ( n9704 & n9906 ) | ( n9704 & n10106 ) | ( n9906 & n10106 ) ;
  assign n10109 = n10106 ^ n9906 ^ n9704 ;
  assign n10110 = n6823 & n7485 ;
  assign n10111 = ( n6747 & n7493 ) | ( n6747 & n10110 ) | ( n7493 & n10110 ) ;
  assign n10112 = n10110 | n10111 ;
  assign n10113 = ( ~n6752 & n7486 ) | ( ~n6752 & n10110 ) | ( n7486 & n10110 ) ;
  assign n10114 = n10112 | n10113 ;
  assign n10115 = n7487 & ~n9943 ;
  assign n10116 = n10114 | n10115 ;
  assign n10117 = n10116 ^ x17 ^ 1'b0 ;
  assign n10118 = ( n9726 & n9845 ) | ( n9726 & n10117 ) | ( n9845 & n10117 ) ;
  assign n10119 = n10117 ^ n9845 ^ n9726 ;
  assign n10120 = n6823 & n7833 ;
  assign n10121 = ( n6751 & n7834 ) | ( n6751 & n10120 ) | ( n7834 & n10120 ) ;
  assign n10122 = n10120 | n10121 ;
  assign n10123 = ( ~n6752 & n7829 ) | ( ~n6752 & n10120 ) | ( n7829 & n10120 ) ;
  assign n10124 = n10122 | n10123 ;
  assign n10125 = n7838 & ~n10013 ;
  assign n10126 = n10124 | n10125 ;
  assign n10127 = n10126 ^ x11 ^ 1'b0 ;
  assign n10128 = ( n9814 & ~n9916 ) | ( n9814 & n10127 ) | ( ~n9916 & n10127 ) ;
  assign n10129 = n10127 ^ n9916 ^ n9814 ;
  assign n10130 = n6751 & n8088 ;
  assign n10131 = ( ~n6477 & n8090 ) | ( ~n6477 & n10130 ) | ( n8090 & n10130 ) ;
  assign n10132 = ( ~n6752 & n8086 ) | ( ~n6752 & n10130 ) | ( n8086 & n10130 ) ;
  assign n10133 = n6751 & n8029 ;
  assign n10134 = n10130 | n10132 ;
  assign n10135 = n10107 ^ n6751 ^ n6477 ;
  assign n10136 = n10131 | n10134 ;
  assign n10137 = ( n8089 & ~n10135 ) | ( n8089 & n10136 ) | ( ~n10135 & n10136 ) ;
  assign n10138 = n10136 | n10137 ;
  assign n10139 = ( ~n6752 & n8037 ) | ( ~n6752 & n10133 ) | ( n8037 & n10133 ) ;
  assign n10140 = n10133 | n10139 ;
  assign n10141 = ( ~n6477 & n8033 ) | ( ~n6477 & n10133 ) | ( n8033 & n10133 ) ;
  assign n10142 = n10140 | n10141 ;
  assign n10143 = n6751 & n7932 ;
  assign n10144 = n10138 ^ x2 ^ 1'b0 ;
  assign n10145 = ( ~n9958 & n10018 ) | ( ~n9958 & n10144 ) | ( n10018 & n10144 ) ;
  assign n10146 = n10144 ^ n10018 ^ n9958 ;
  assign n10147 = n8034 & ~n10135 ;
  assign n10148 = ( ~n6752 & n7943 ) | ( ~n6752 & n10143 ) | ( n7943 & n10143 ) ;
  assign n10149 = n10143 | n10148 ;
  assign n10150 = ( ~n6477 & n7929 ) | ( ~n6477 & n10143 ) | ( n7929 & n10143 ) ;
  assign n10151 = n10149 | n10150 ;
  assign n10152 = n7930 & ~n10135 ;
  assign n10153 = n10151 | n10152 ;
  assign n10154 = n6751 & n7943 ;
  assign n10155 = n10142 | n10147 ;
  assign n10156 = n10155 ^ x5 ^ 1'b0 ;
  assign n10157 = n10153 ^ x8 ^ 1'b0 ;
  assign n10158 = n10157 ^ n9894 ^ n9884 ;
  assign n10159 = ( n9884 & n9894 ) | ( n9884 & n10157 ) | ( n9894 & n10157 ) ;
  assign n10160 = n6751 & n8037 ;
  assign n10161 = ( ~n6477 & n8029 ) | ( ~n6477 & n10160 ) | ( n8029 & n10160 ) ;
  assign n10162 = n10160 | n10161 ;
  assign n10163 = ( ~n6477 & n6751 ) | ( ~n6477 & n10107 ) | ( n6751 & n10107 ) ;
  assign n10164 = ( ~n6004 & n8033 ) | ( ~n6004 & n10160 ) | ( n8033 & n10160 ) ;
  assign n10165 = n10162 | n10164 ;
  assign n10166 = n10156 ^ n10088 ^ n10058 ;
  assign n10167 = ( ~n10058 & n10088 ) | ( ~n10058 & n10156 ) | ( n10088 & n10156 ) ;
  assign n10168 = n10163 ^ n6477 ^ n6004 ;
  assign n10169 = n8034 & n10168 ;
  assign n10170 = n10165 | n10169 ;
  assign n10171 = ( ~n6477 & n7932 ) | ( ~n6477 & n10154 ) | ( n7932 & n10154 ) ;
  assign n10172 = n10154 | n10171 ;
  assign n10173 = ( ~n6004 & n7929 ) | ( ~n6004 & n10154 ) | ( n7929 & n10154 ) ;
  assign n10174 = n10170 ^ x5 ^ 1'b0 ;
  assign n10175 = n10172 | n10173 ;
  assign n10176 = ( n10067 & n10167 ) | ( n10067 & n10174 ) | ( n10167 & n10174 ) ;
  assign n10177 = n10174 ^ n10167 ^ n10067 ;
  assign n10178 = n6751 & n8086 ;
  assign n10179 = ( ~n6477 & n8088 ) | ( ~n6477 & n10178 ) | ( n8088 & n10178 ) ;
  assign n10180 = n10178 | n10179 ;
  assign n10181 = ( ~n6004 & n8090 ) | ( ~n6004 & n10178 ) | ( n8090 & n10178 ) ;
  assign n10182 = n10180 | n10181 ;
  assign n10183 = ( n8089 & n10168 ) | ( n8089 & n10182 ) | ( n10168 & n10182 ) ;
  assign n10184 = n10182 | n10183 ;
  assign n10185 = n7930 & n10168 ;
  assign n10186 = n10175 | n10185 ;
  assign n10187 = n10184 ^ x2 ^ 1'b0 ;
  assign n10188 = n10186 ^ x8 ^ 1'b0 ;
  assign n10189 = n10188 ^ n10035 ^ n9885 ;
  assign n10190 = ( n9885 & n10035 ) | ( n9885 & n10188 ) | ( n10035 & n10188 ) ;
  assign n10191 = ~n6477 & n8086 ;
  assign n10192 = ( ~n6004 & n8088 ) | ( ~n6004 & n10191 ) | ( n8088 & n10191 ) ;
  assign n10193 = n10191 | n10192 ;
  assign n10194 = ( ~n6707 & n8090 ) | ( ~n6707 & n10191 ) | ( n8090 & n10191 ) ;
  assign n10195 = n10193 | n10194 ;
  assign n10196 = n10187 ^ n10145 ^ n9966 ;
  assign n10197 = ( n6004 & n6477 ) | ( n6004 & ~n10163 ) | ( n6477 & ~n10163 ) ;
  assign n10198 = ( ~n9966 & n10145 ) | ( ~n9966 & n10187 ) | ( n10145 & n10187 ) ;
  assign n10199 = ( n6004 & n6707 ) | ( n6004 & n10197 ) | ( n6707 & n10197 ) ;
  assign n10200 = n10197 ^ n6707 ^ n6004 ;
  assign n10201 = ( n8089 & n10195 ) | ( n8089 & ~n10200 ) | ( n10195 & ~n10200 ) ;
  assign n10202 = n10195 | n10201 ;
  assign n10203 = n10202 ^ x2 ^ 1'b0 ;
  assign n10204 = ( n10087 & n10198 ) | ( n10087 & n10203 ) | ( n10198 & n10203 ) ;
  assign n10205 = n10203 ^ n10198 ^ n10087 ;
  assign n10206 = ~n6004 & n8029 ;
  assign n10207 = ~n6004 & n8086 ;
  assign n10208 = ( ~n6707 & n8088 ) | ( ~n6707 & n10207 ) | ( n8088 & n10207 ) ;
  assign n10209 = ~n6707 & n8029 ;
  assign n10210 = ( ~n6004 & n8037 ) | ( ~n6004 & n10209 ) | ( n8037 & n10209 ) ;
  assign n10211 = n10209 | n10210 ;
  assign n10212 = ( n8033 & ~n9912 ) | ( n8033 & n10209 ) | ( ~n9912 & n10209 ) ;
  assign n10213 = n10199 ^ n9912 ^ n6707 ;
  assign n10214 = ( ~n6477 & n8037 ) | ( ~n6477 & n10206 ) | ( n8037 & n10206 ) ;
  assign n10215 = n10207 | n10208 ;
  assign n10216 = n10206 | n10214 ;
  assign n10217 = ( n8090 & ~n9912 ) | ( n8090 & n10207 ) | ( ~n9912 & n10207 ) ;
  assign n10218 = n10215 | n10217 ;
  assign n10219 = ( n8089 & ~n10213 ) | ( n8089 & n10218 ) | ( ~n10213 & n10218 ) ;
  assign n10220 = ( ~n6707 & n8033 ) | ( ~n6707 & n10206 ) | ( n8033 & n10206 ) ;
  assign n10221 = n10218 | n10219 ;
  assign n10222 = n10211 | n10212 ;
  assign n10223 = ~n6004 & n7932 ;
  assign n10224 = n10216 | n10220 ;
  assign n10225 = n8034 & ~n10200 ;
  assign n10226 = n10224 | n10225 ;
  assign n10227 = ( ~n6477 & n7943 ) | ( ~n6477 & n10223 ) | ( n7943 & n10223 ) ;
  assign n10228 = n8034 & ~n10213 ;
  assign n10229 = n10223 | n10227 ;
  assign n10230 = ( ~n6707 & n7929 ) | ( ~n6707 & n10223 ) | ( n7929 & n10223 ) ;
  assign n10231 = n10229 | n10230 ;
  assign n10232 = n10221 ^ x2 ^ 1'b0 ;
  assign n10233 = n10232 ^ n10204 ^ n10166 ;
  assign n10234 = ( ~n10166 & n10204 ) | ( ~n10166 & n10232 ) | ( n10204 & n10232 ) ;
  assign n10235 = ( n6707 & n9912 ) | ( n6707 & n10199 ) | ( n9912 & n10199 ) ;
  assign n10236 = n7930 & ~n10200 ;
  assign n10237 = n10222 | n10228 ;
  assign n10238 = n10231 | n10236 ;
  assign n10239 = n10238 ^ x8 ^ 1'b0 ;
  assign n10240 = n10237 ^ x5 ^ 1'b0 ;
  assign n10241 = n9912 | n10235 ;
  assign n10242 = n8089 & ~n10241 ;
  assign n10243 = ( n8086 & ~n9912 ) | ( n8086 & n10242 ) | ( ~n9912 & n10242 ) ;
  assign n10244 = n10242 | n10243 ;
  assign n10245 = ( n10034 & ~n10129 ) | ( n10034 & n10239 ) | ( ~n10129 & n10239 ) ;
  assign n10246 = n10244 ^ x2 ^ 1'b0 ;
  assign n10247 = n10239 ^ n10129 ^ n10034 ;
  assign n10248 = n8034 & ~n10241 ;
  assign n10249 = n8037 & ~n9912 ;
  assign n10250 = ~n10248 & n10249 ;
  assign n10251 = n10235 ^ n9912 ^ 1'b0 ;
  assign n10252 = n10250 ^ n10248 ^ x5 ;
  assign n10253 = n10252 ^ n10247 ^ n10190 ;
  assign n10254 = ( n10190 & ~n10247 ) | ( n10190 & n10252 ) | ( ~n10247 & n10252 ) ;
  assign n10255 = n8089 & n10251 ;
  assign n10256 = ( ~n6707 & n8086 ) | ( ~n6707 & n10255 ) | ( n8086 & n10255 ) ;
  assign n10257 = n10255 | n10256 ;
  assign n10258 = ( n8088 & ~n9912 ) | ( n8088 & n10255 ) | ( ~n9912 & n10255 ) ;
  assign n10259 = n10257 | n10258 ;
  assign n10260 = n10259 ^ x2 ^ 1'b0 ;
  assign n10261 = n10260 ^ n10234 ^ n10177 ;
  assign n10262 = ( n10177 & n10234 ) | ( n10177 & n10260 ) | ( n10234 & n10260 ) ;
  assign n10263 = n10240 ^ n10158 ^ n10097 ;
  assign n10264 = n8034 & n10251 ;
  assign n10265 = n10226 ^ x5 ^ 1'b0 ;
  assign n10266 = ( n10097 & n10158 ) | ( n10097 & n10240 ) | ( n10158 & n10240 ) ;
  assign n10267 = ( n8029 & ~n9912 ) | ( n8029 & n10264 ) | ( ~n9912 & n10264 ) ;
  assign n10268 = n10265 ^ n10246 ^ n10098 ;
  assign n10269 = n10264 | n10267 ;
  assign n10270 = ( ~n6707 & n8037 ) | ( ~n6707 & n10264 ) | ( n8037 & n10264 ) ;
  assign n10271 = n10269 | n10270 ;
  assign n10272 = ( n10098 & n10246 ) | ( n10098 & n10265 ) | ( n10246 & n10265 ) ;
  assign n10273 = ( n10176 & n10262 ) | ( n10176 & n10268 ) | ( n10262 & n10268 ) ;
  assign n10274 = n10271 ^ x5 ^ 1'b0 ;
  assign n10275 = ( n10159 & n10189 ) | ( n10159 & n10274 ) | ( n10189 & n10274 ) ;
  assign n10276 = ( n10263 & n10272 ) | ( n10263 & n10273 ) | ( n10272 & n10273 ) ;
  assign n10277 = n10274 ^ n10189 ^ n10159 ;
  assign n10278 = n10277 ^ n10276 ^ n10266 ;
  assign n10279 = ( n10266 & n10276 ) | ( n10266 & n10277 ) | ( n10276 & n10277 ) ;
  assign n10280 = n10279 ^ n10275 ^ n10253 ;
  assign n10281 = ( ~n10253 & n10275 ) | ( ~n10253 & n10279 ) | ( n10275 & n10279 ) ;
  assign n10282 = n10273 ^ n10272 ^ n10263 ;
  assign n10283 = n10268 ^ n10262 ^ n10176 ;
  assign n10284 = n6751 & n7829 ;
  assign n10285 = ( ~n6752 & n7833 ) | ( ~n6752 & n10284 ) | ( n7833 & n10284 ) ;
  assign n10286 = n10284 | n10285 ;
  assign n10287 = ( ~n6477 & n7834 ) | ( ~n6477 & n10284 ) | ( n7834 & n10284 ) ;
  assign n10288 = n10286 | n10287 ;
  assign n10289 = ( n7838 & ~n10135 ) | ( n7838 & n10288 ) | ( ~n10135 & n10288 ) ;
  assign n10290 = n10288 | n10289 ;
  assign n10291 = n10290 ^ x11 ^ 1'b0 ;
  assign n10292 = ( n10007 & n10128 ) | ( n10007 & n10291 ) | ( n10128 & n10291 ) ;
  assign n10293 = n10291 ^ n10128 ^ n10007 ;
  assign n10294 = ~n6707 & n7932 ;
  assign n10295 = ( ~n6004 & n7943 ) | ( ~n6004 & n10294 ) | ( n7943 & n10294 ) ;
  assign n10296 = n10294 | n10295 ;
  assign n10297 = ( n7929 & ~n9912 ) | ( n7929 & n10294 ) | ( ~n9912 & n10294 ) ;
  assign n10298 = n10296 | n10297 ;
  assign n10299 = ( n7930 & ~n10213 ) | ( n7930 & n10298 ) | ( ~n10213 & n10298 ) ;
  assign n10300 = n10298 | n10299 ;
  assign n10301 = n10300 ^ x8 ^ 1'b0 ;
  assign n10302 = ( n10245 & n10293 ) | ( n10245 & n10301 ) | ( n10293 & n10301 ) ;
  assign n10303 = n10301 ^ n10293 ^ n10245 ;
  assign n10304 = n6751 & n7669 ;
  assign n10305 = ( n10254 & n10281 ) | ( n10254 & n10303 ) | ( n10281 & n10303 ) ;
  assign n10306 = n10303 ^ n10281 ^ n10254 ;
  assign n10307 = n6751 & n7833 ;
  assign n10308 = ( ~n6752 & n7674 ) | ( ~n6752 & n10304 ) | ( n7674 & n10304 ) ;
  assign n10309 = n10304 | n10308 ;
  assign n10310 = ( ~n6477 & n7667 ) | ( ~n6477 & n10304 ) | ( n7667 & n10304 ) ;
  assign n10311 = n10309 | n10310 ;
  assign n10312 = ( n7666 & ~n10135 ) | ( n7666 & n10311 ) | ( ~n10135 & n10311 ) ;
  assign n10313 = n10311 | n10312 ;
  assign n10314 = ( ~n6477 & n7829 ) | ( ~n6477 & n10307 ) | ( n7829 & n10307 ) ;
  assign n10315 = n10307 | n10314 ;
  assign n10316 = ( ~n6004 & n7834 ) | ( ~n6004 & n10307 ) | ( n7834 & n10307 ) ;
  assign n10317 = n10313 ^ x14 ^ 1'b0 ;
  assign n10318 = n10315 | n10316 ;
  assign n10319 = n7838 & n10168 ;
  assign n10320 = n10318 | n10319 ;
  assign n10321 = n10317 ^ n10077 ^ n9996 ;
  assign n10322 = ( n9996 & n10077 ) | ( n9996 & n10317 ) | ( n10077 & n10317 ) ;
  assign n10323 = n10320 ^ x11 ^ 1'b0 ;
  assign n10324 = n7930 & n10251 ;
  assign n10325 = ( n7932 & ~n9912 ) | ( n7932 & n10324 ) | ( ~n9912 & n10324 ) ;
  assign n10326 = n10324 | n10325 ;
  assign n10327 = ( ~n6707 & n7943 ) | ( ~n6707 & n10324 ) | ( n7943 & n10324 ) ;
  assign n10328 = n10326 | n10327 ;
  assign n10329 = n10323 ^ n10006 ^ n9985 ;
  assign n10330 = ( ~n9985 & n10006 ) | ( ~n9985 & n10323 ) | ( n10006 & n10323 ) ;
  assign n10331 = n7943 & ~n9912 ;
  assign n10332 = n7930 & ~n10241 ;
  assign n10333 = n10331 & ~n10332 ;
  assign n10334 = n10328 ^ x8 ^ 1'b0 ;
  assign n10335 = n10333 ^ n10332 ^ x8 ;
  assign n10336 = n10334 ^ n10329 ^ n10292 ;
  assign n10337 = ( n10292 & ~n10329 ) | ( n10292 & n10334 ) | ( ~n10329 & n10334 ) ;
  assign n10338 = ( n10302 & n10305 ) | ( n10302 & ~n10336 ) | ( n10305 & ~n10336 ) ;
  assign n10339 = n7838 & ~n10200 ;
  assign n10340 = n10336 ^ n10305 ^ n10302 ;
  assign n10341 = ~n6004 & n7829 ;
  assign n10342 = ( ~n6477 & n7833 ) | ( ~n6477 & n10341 ) | ( n7833 & n10341 ) ;
  assign n10343 = n10341 | n10342 ;
  assign n10344 = ( ~n6707 & n7834 ) | ( ~n6707 & n10341 ) | ( n7834 & n10341 ) ;
  assign n10345 = n10343 | n10344 ;
  assign n10346 = n10339 | n10345 ;
  assign n10347 = n10346 ^ x11 ^ 1'b0 ;
  assign n10348 = n10347 ^ n10078 ^ n9984 ;
  assign n10349 = ( n10330 & n10335 ) | ( n10330 & n10348 ) | ( n10335 & n10348 ) ;
  assign n10350 = n10348 ^ n10335 ^ n10330 ;
  assign n10351 = ( n9984 & n10078 ) | ( n9984 & n10347 ) | ( n10078 & n10347 ) ;
  assign n10352 = ( n10337 & n10338 ) | ( n10337 & n10350 ) | ( n10338 & n10350 ) ;
  assign n10353 = n10350 ^ n10338 ^ n10337 ;
  assign n10354 = ~n6707 & n7829 ;
  assign n10355 = ( ~n6004 & n7833 ) | ( ~n6004 & n10354 ) | ( n7833 & n10354 ) ;
  assign n10356 = n10354 | n10355 ;
  assign n10357 = ( n7834 & ~n9912 ) | ( n7834 & n10354 ) | ( ~n9912 & n10354 ) ;
  assign n10358 = n10356 | n10357 ;
  assign n10359 = ( n7838 & ~n10213 ) | ( n7838 & n10358 ) | ( ~n10213 & n10358 ) ;
  assign n10360 = n10358 | n10359 ;
  assign n10361 = n10360 ^ x11 ^ 1'b0 ;
  assign n10362 = n10361 ^ n10351 ^ n10321 ;
  assign n10363 = ( n10321 & n10351 ) | ( n10321 & n10361 ) | ( n10351 & n10361 ) ;
  assign n10364 = ~n6004 & n7669 ;
  assign n10365 = ( ~n6477 & n7674 ) | ( ~n6477 & n10364 ) | ( n7674 & n10364 ) ;
  assign n10366 = n10364 | n10365 ;
  assign n10367 = ( ~n6707 & n7667 ) | ( ~n6707 & n10364 ) | ( n7667 & n10364 ) ;
  assign n10368 = n10366 | n10367 ;
  assign n10369 = n7666 & ~n10200 ;
  assign n10370 = n10368 | n10369 ;
  assign n10371 = ( n10349 & n10352 ) | ( n10349 & n10362 ) | ( n10352 & n10362 ) ;
  assign n10372 = n10362 ^ n10352 ^ n10349 ;
  assign n10373 = n6751 & n7674 ;
  assign n10374 = n10370 ^ x14 ^ 1'b0 ;
  assign n10375 = ( ~n6477 & n7669 ) | ( ~n6477 & n10373 ) | ( n7669 & n10373 ) ;
  assign n10376 = n10373 | n10375 ;
  assign n10377 = ( ~n6004 & n7667 ) | ( ~n6004 & n10373 ) | ( n7667 & n10373 ) ;
  assign n10378 = n10376 | n10377 ;
  assign n10379 = ( n10048 & n10118 ) | ( n10048 & n10374 ) | ( n10118 & n10374 ) ;
  assign n10380 = n10374 ^ n10118 ^ n10048 ;
  assign n10381 = n7838 & ~n10241 ;
  assign n10382 = n7666 & n10168 ;
  assign n10383 = n10378 | n10382 ;
  assign n10384 = n10383 ^ x14 ^ 1'b0 ;
  assign n10385 = n10384 ^ n10119 ^ n9997 ;
  assign n10386 = ( n9997 & n10119 ) | ( n9997 & n10384 ) | ( n10119 & n10384 ) ;
  assign n10387 = n6751 & n7485 ;
  assign n10388 = ( ~n6477 & n7486 ) | ( ~n6477 & n10387 ) | ( n7486 & n10387 ) ;
  assign n10389 = n10387 | n10388 ;
  assign n10390 = ( ~n6752 & n7493 ) | ( ~n6752 & n10387 ) | ( n7493 & n10387 ) ;
  assign n10391 = n10389 | n10390 ;
  assign n10392 = n7487 & ~n10135 ;
  assign n10393 = n10391 | n10392 ;
  assign n10394 = n10393 ^ x17 ^ 1'b0 ;
  assign n10395 = ( n10047 & n10109 ) | ( n10047 & n10394 ) | ( n10109 & n10394 ) ;
  assign n10396 = n10394 ^ n10109 ^ n10047 ;
  assign n10397 = n7838 & n10251 ;
  assign n10398 = n7833 & ~n9912 ;
  assign n10399 = ~n10381 & n10398 ;
  assign n10400 = n10399 ^ n10381 ^ x11 ;
  assign n10401 = ( n7829 & ~n9912 ) | ( n7829 & n10397 ) | ( ~n9912 & n10397 ) ;
  assign n10402 = n10397 | n10401 ;
  assign n10403 = ( ~n6707 & n7833 ) | ( ~n6707 & n10397 ) | ( n7833 & n10397 ) ;
  assign n10404 = n10402 | n10403 ;
  assign n10405 = n10404 ^ x11 ^ 1'b0 ;
  assign n10406 = n10405 ^ n10385 ^ n10322 ;
  assign n10407 = ( n10322 & n10385 ) | ( n10322 & n10405 ) | ( n10385 & n10405 ) ;
  assign n10408 = n10406 ^ n10371 ^ n10363 ;
  assign n10409 = ( n10363 & n10371 ) | ( n10363 & n10406 ) | ( n10371 & n10406 ) ;
  assign n10410 = ~n6707 & n7669 ;
  assign n10411 = ( ~n6004 & n7674 ) | ( ~n6004 & n10410 ) | ( n7674 & n10410 ) ;
  assign n10412 = n10410 | n10411 ;
  assign n10413 = ( n10380 & n10386 ) | ( n10380 & n10400 ) | ( n10386 & n10400 ) ;
  assign n10414 = n10400 ^ n10386 ^ n10380 ;
  assign n10415 = ( n7667 & ~n9912 ) | ( n7667 & n10410 ) | ( ~n9912 & n10410 ) ;
  assign n10416 = ( n10407 & n10409 ) | ( n10407 & n10414 ) | ( n10409 & n10414 ) ;
  assign n10417 = n10412 | n10415 ;
  assign n10418 = ( n7666 & ~n10213 ) | ( n7666 & n10417 ) | ( ~n10213 & n10417 ) ;
  assign n10419 = n10414 ^ n10409 ^ n10407 ;
  assign n10420 = n10417 | n10418 ;
  assign n10421 = n10420 ^ x14 ^ 1'b0 ;
  assign n10422 = ( n10379 & n10396 ) | ( n10379 & n10421 ) | ( n10396 & n10421 ) ;
  assign n10423 = n10421 ^ n10396 ^ n10379 ;
  assign n10424 = ( n10413 & n10416 ) | ( n10413 & n10423 ) | ( n10416 & n10423 ) ;
  assign n10425 = n10423 ^ n10416 ^ n10413 ;
  assign n10426 = n6747 & n7188 ;
  assign n10427 = ( ~n6741 & n7190 ) | ( ~n6741 & n10426 ) | ( n7190 & n10426 ) ;
  assign n10428 = n10426 | n10427 ;
  assign n10429 = ( ~n6746 & n7192 ) | ( ~n6746 & n10426 ) | ( n7192 & n10426 ) ;
  assign n10430 = n10428 | n10429 ;
  assign n10431 = n7196 & n9865 ;
  assign n10432 = n10430 | n10431 ;
  assign n10433 = n10432 ^ x23 ^ 1'b0 ;
  assign n10434 = ( n9494 & n9588 ) | ( n9494 & n10433 ) | ( n9588 & n10433 ) ;
  assign n10435 = n10433 ^ n9588 ^ n9494 ;
  assign n10436 = n6823 & n7338 ;
  assign n10437 = ( n6751 & n7337 ) | ( n6751 & n10436 ) | ( n7337 & n10436 ) ;
  assign n10438 = n10436 | n10437 ;
  assign n10439 = ( ~n6752 & n7339 ) | ( ~n6752 & n10436 ) | ( n7339 & n10436 ) ;
  assign n10440 = n10438 | n10439 ;
  assign n10441 = n7340 & ~n10013 ;
  assign n10442 = n10440 | n10441 ;
  assign n10443 = n10442 ^ x20 ^ 1'b0 ;
  assign n10444 = ( n9824 & n10435 ) | ( n9824 & n10443 ) | ( n10435 & n10443 ) ;
  assign n10445 = n10443 ^ n10435 ^ n9824 ;
  assign n10446 = n6823 & n7339 ;
  assign n10447 = ( n6747 & n7338 ) | ( n6747 & n10446 ) | ( n7338 & n10446 ) ;
  assign n10448 = n10446 | n10447 ;
  assign n10449 = ( ~n6752 & n7337 ) | ( ~n6752 & n10446 ) | ( n7337 & n10446 ) ;
  assign n10450 = n10448 | n10449 ;
  assign n10451 = n7340 & ~n9943 ;
  assign n10452 = n10450 | n10451 ;
  assign n10453 = n10452 ^ x20 ^ 1'b0 ;
  assign n10454 = ( n9703 & n9825 ) | ( n9703 & n10453 ) | ( n9825 & n10453 ) ;
  assign n10455 = n10453 ^ n9825 ^ n9703 ;
  assign n10456 = n6751 & n7493 ;
  assign n10457 = ( ~n6477 & n7485 ) | ( ~n6477 & n10456 ) | ( n7485 & n10456 ) ;
  assign n10458 = n10456 | n10457 ;
  assign n10459 = ( ~n6004 & n7486 ) | ( ~n6004 & n10456 ) | ( n7486 & n10456 ) ;
  assign n10460 = n10458 | n10459 ;
  assign n10461 = n7487 & n10168 ;
  assign n10462 = n10460 | n10461 ;
  assign n10463 = n10462 ^ x17 ^ 1'b0 ;
  assign n10464 = ( n10108 & n10455 ) | ( n10108 & n10463 ) | ( n10455 & n10463 ) ;
  assign n10465 = n10463 ^ n10455 ^ n10108 ;
  assign n10466 = ~n6004 & n7485 ;
  assign n10467 = ( ~n6707 & n7486 ) | ( ~n6707 & n10466 ) | ( n7486 & n10466 ) ;
  assign n10468 = n10466 | n10467 ;
  assign n10469 = ( ~n6477 & n7493 ) | ( ~n6477 & n10466 ) | ( n7493 & n10466 ) ;
  assign n10470 = n10468 | n10469 ;
  assign n10471 = n7487 & ~n10200 ;
  assign n10472 = n10470 | n10471 ;
  assign n10473 = n10472 ^ x17 ^ 1'b0 ;
  assign n10474 = ( n10445 & n10454 ) | ( n10445 & n10473 ) | ( n10454 & n10473 ) ;
  assign n10475 = n10473 ^ n10454 ^ n10445 ;
  assign n10476 = n7674 & ~n9912 ;
  assign n10477 = n7666 & ~n10241 ;
  assign n10478 = n10476 & ~n10477 ;
  assign n10479 = n10478 ^ n10477 ^ x14 ;
  assign n10480 = n10479 ^ n10475 ^ n10464 ;
  assign n10481 = ( n10464 & n10475 ) | ( n10464 & n10479 ) | ( n10475 & n10479 ) ;
  assign n10482 = n7666 & n10251 ;
  assign n10483 = ( n7669 & ~n9912 ) | ( n7669 & n10482 ) | ( ~n9912 & n10482 ) ;
  assign n10484 = n10482 | n10483 ;
  assign n10485 = ( ~n6707 & n7674 ) | ( ~n6707 & n10482 ) | ( n7674 & n10482 ) ;
  assign n10486 = n10484 | n10485 ;
  assign n10487 = n10486 ^ x14 ^ 1'b0 ;
  assign n10488 = ( n10395 & n10465 ) | ( n10395 & n10487 ) | ( n10465 & n10487 ) ;
  assign n10489 = n10487 ^ n10465 ^ n10395 ;
  assign n10490 = ( n10422 & n10424 ) | ( n10422 & n10489 ) | ( n10424 & n10489 ) ;
  assign n10491 = n10489 ^ n10424 ^ n10422 ;
  assign n10492 = n10490 ^ n10488 ^ n10480 ;
  assign n10493 = ( n10480 & n10488 ) | ( n10480 & n10490 ) | ( n10488 & n10490 ) ;
  assign n10494 = n6823 & n7188 ;
  assign n10495 = ( n6747 & n7192 ) | ( n6747 & n10494 ) | ( n7192 & n10494 ) ;
  assign n10496 = n10494 | n10495 ;
  assign n10497 = ( ~n6746 & n7190 ) | ( ~n6746 & n10494 ) | ( n7190 & n10494 ) ;
  assign n10498 = n10496 | n10497 ;
  assign n10499 = n7196 & ~n9877 ;
  assign n10500 = n10498 | n10499 ;
  assign n10501 = n10500 ^ x23 ^ 1'b0 ;
  assign n10502 = ( ~n9746 & n10434 ) | ( ~n9746 & n10501 ) | ( n10434 & n10501 ) ;
  assign n10503 = n10501 ^ n10434 ^ n9746 ;
  assign n10504 = n6751 & n7339 ;
  assign n10505 = ( ~n6477 & n7337 ) | ( ~n6477 & n10504 ) | ( n7337 & n10504 ) ;
  assign n10506 = n10504 | n10505 ;
  assign n10507 = ( ~n6752 & n7338 ) | ( ~n6752 & n10504 ) | ( n7338 & n10504 ) ;
  assign n10508 = n10506 | n10507 ;
  assign n10509 = ( n7340 & ~n10135 ) | ( n7340 & n10508 ) | ( ~n10135 & n10508 ) ;
  assign n10510 = n10508 | n10509 ;
  assign n10511 = n10510 ^ x20 ^ 1'b0 ;
  assign n10512 = ( n10444 & ~n10503 ) | ( n10444 & n10511 ) | ( ~n10503 & n10511 ) ;
  assign n10513 = n10511 ^ n10503 ^ n10444 ;
  assign n10514 = n6823 & n7192 ;
  assign n10515 = ( n6747 & n7190 ) | ( n6747 & n10514 ) | ( n7190 & n10514 ) ;
  assign n10516 = n10514 | n10515 ;
  assign n10517 = ( ~n6752 & n7188 ) | ( ~n6752 & n10514 ) | ( n7188 & n10514 ) ;
  assign n10518 = n10516 | n10517 ;
  assign n10519 = n7196 & ~n9943 ;
  assign n10520 = n10518 | n10519 ;
  assign n10521 = n10520 ^ x23 ^ 1'b0 ;
  assign n10522 = ( n9745 & n9861 ) | ( n9745 & n10521 ) | ( n9861 & n10521 ) ;
  assign n10523 = n10521 ^ n9861 ^ n9745 ;
  assign n10524 = ~n6707 & n7485 ;
  assign n10525 = ( n7486 & ~n9912 ) | ( n7486 & n10524 ) | ( ~n9912 & n10524 ) ;
  assign n10526 = n10524 | n10525 ;
  assign n10527 = ( ~n6004 & n7493 ) | ( ~n6004 & n10524 ) | ( n7493 & n10524 ) ;
  assign n10528 = n10526 | n10527 ;
  assign n10529 = ( n7487 & ~n10213 ) | ( n7487 & n10528 ) | ( ~n10213 & n10528 ) ;
  assign n10530 = n10528 | n10529 ;
  assign n10531 = n10530 ^ x17 ^ 1'b0 ;
  assign n10532 = n10531 ^ n10513 ^ n10474 ;
  assign n10533 = ( n10474 & ~n10513 ) | ( n10474 & n10531 ) | ( ~n10513 & n10531 ) ;
  assign n10534 = n6751 & n7338 ;
  assign n10535 = ( ~n6477 & n7339 ) | ( ~n6477 & n10534 ) | ( n7339 & n10534 ) ;
  assign n10536 = n10534 | n10535 ;
  assign n10537 = ( ~n6004 & n7337 ) | ( ~n6004 & n10534 ) | ( n7337 & n10534 ) ;
  assign n10538 = n10536 | n10537 ;
  assign n10539 = n10532 ^ n10493 ^ n10481 ;
  assign n10540 = ( n10481 & n10493 ) | ( n10481 & ~n10532 ) | ( n10493 & ~n10532 ) ;
  assign n10541 = n7487 & n10251 ;
  assign n10542 = n7340 & n10168 ;
  assign n10543 = n10538 | n10542 ;
  assign n10544 = ( n7485 & ~n9912 ) | ( n7485 & n10541 ) | ( ~n9912 & n10541 ) ;
  assign n10545 = n10541 | n10544 ;
  assign n10546 = ( ~n6707 & n7493 ) | ( ~n6707 & n10541 ) | ( n7493 & n10541 ) ;
  assign n10547 = n10543 ^ x20 ^ 1'b0 ;
  assign n10548 = n10545 | n10546 ;
  assign n10549 = n10548 ^ x17 ^ 1'b0 ;
  assign n10550 = n10547 ^ n10523 ^ n10502 ;
  assign n10551 = ( n10502 & n10523 ) | ( n10502 & n10547 ) | ( n10523 & n10547 ) ;
  assign n10552 = ( n10512 & n10549 ) | ( n10512 & n10550 ) | ( n10549 & n10550 ) ;
  assign n10553 = n10550 ^ n10549 ^ n10512 ;
  assign n10554 = ( n10533 & n10540 ) | ( n10533 & n10553 ) | ( n10540 & n10553 ) ;
  assign n10555 = n10553 ^ n10540 ^ n10533 ;
  assign n10556 = ( n6308 & n9706 ) | ( n6308 & n9859 ) | ( n9706 & n9859 ) ;
  assign n10557 = n6747 & n7037 ;
  assign n10558 = ( ~n6746 & n7036 ) | ( ~n6746 & n10557 ) | ( n7036 & n10557 ) ;
  assign n10559 = n10557 | n10558 ;
  assign n10560 = ( ~n6741 & n7052 ) | ( ~n6741 & n10557 ) | ( n7052 & n10557 ) ;
  assign n10561 = n10559 | n10560 ;
  assign n10562 = n7035 & n9865 ;
  assign n10563 = n10561 | n10562 ;
  assign n10564 = n10563 ^ x26 ^ 1'b0 ;
  assign n10565 = ( n9483 & ~n9674 ) | ( n9483 & n10564 ) | ( ~n9674 & n10564 ) ;
  assign n10566 = n10564 ^ n9674 ^ n9483 ;
  assign n10567 = n6823 & n7037 ;
  assign n10568 = ( n6747 & n7036 ) | ( n6747 & n10567 ) | ( n7036 & n10567 ) ;
  assign n10569 = n10567 | n10568 ;
  assign n10570 = n9859 ^ n9706 ^ n6308 ;
  assign n10571 = ( ~n6746 & n7052 ) | ( ~n6746 & n10567 ) | ( n7052 & n10567 ) ;
  assign n10572 = n10569 | n10571 ;
  assign n10573 = ( n7035 & ~n9877 ) | ( n7035 & n10572 ) | ( ~n9877 & n10572 ) ;
  assign n10574 = ( n6308 & n6700 ) | ( n6308 & ~n10556 ) | ( n6700 & ~n10556 ) ;
  assign n10575 = n10572 | n10573 ;
  assign n10576 = n10575 ^ x26 ^ 1'b0 ;
  assign n10577 = n10556 ^ n6700 ^ n6308 ;
  assign n10578 = n10576 ^ n10565 ^ n9756 ;
  assign n10579 = ( n9756 & n10565 ) | ( n9756 & n10576 ) | ( n10565 & n10576 ) ;
  assign n10580 = n6789 & n9865 ;
  assign n10581 = ( ~x23 & n6700 ) | ( ~x23 & n6761 ) | ( n6700 & n6761 ) ;
  assign n10582 = ( ~n6746 & n6791 ) | ( ~n6746 & n10580 ) | ( n6791 & n10580 ) ;
  assign n10583 = n10580 | n10582 ;
  assign n10584 = ( ~n6741 & n6790 ) | ( ~n6741 & n10580 ) | ( n6790 & n10580 ) ;
  assign n10585 = n6761 ^ n6700 ^ x23 ;
  assign n10586 = n6747 & n6907 ;
  assign n10587 = n10583 | n10584 ;
  assign n10588 = n6747 & ~n6788 ;
  assign n10589 = ( n6747 & n10587 ) | ( n6747 & ~n10588 ) | ( n10587 & ~n10588 ) ;
  assign n10590 = ( ~n6746 & n6901 ) | ( ~n6746 & n10586 ) | ( n6901 & n10586 ) ;
  assign n10591 = n10586 | n10590 ;
  assign n10592 = ( ~n6741 & n6906 ) | ( ~n6741 & n10586 ) | ( n6906 & n10586 ) ;
  assign n10593 = n10591 | n10592 ;
  assign n10594 = n6918 & ~n9877 ;
  assign n10595 = ( n6918 & n9865 ) | ( n6918 & n10593 ) | ( n9865 & n10593 ) ;
  assign n10596 = n10593 | n10595 ;
  assign n10597 = n6789 & ~n9877 ;
  assign n10598 = ( n6747 & n6791 ) | ( n6747 & n10597 ) | ( n6791 & n10597 ) ;
  assign n10599 = n10597 | n10598 ;
  assign n10600 = n6823 & n6907 ;
  assign n10601 = ( ~n6746 & n6790 ) | ( ~n6746 & n10597 ) | ( n6790 & n10597 ) ;
  assign n10602 = ( ~n6746 & n6906 ) | ( ~n6746 & n10600 ) | ( n6906 & n10600 ) ;
  assign n10603 = n10599 | n10601 ;
  assign n10604 = ~n6788 & n6823 ;
  assign n10605 = ( n6823 & n10603 ) | ( n6823 & ~n10604 ) | ( n10603 & ~n10604 ) ;
  assign n10606 = ( n10574 & n10585 ) | ( n10574 & ~n10605 ) | ( n10585 & ~n10605 ) ;
  assign n10607 = n10605 ^ n10585 ^ n10574 ;
  assign n10608 = ( n6747 & n6901 ) | ( n6747 & n10600 ) | ( n6901 & n10600 ) ;
  assign n10609 = n10600 | n10608 ;
  assign n10610 = n10602 | n10609 ;
  assign n10611 = n10594 | n10610 ;
  assign n10612 = n10611 ^ x29 ^ 1'b0 ;
  assign n10613 = n10612 ^ n9775 ^ n9684 ;
  assign n10614 = ( n9684 & n9775 ) | ( n9684 & n10612 ) | ( n9775 & n10612 ) ;
  assign n10615 = n6823 & n7036 ;
  assign n10616 = ( n6747 & n7052 ) | ( n6747 & n10615 ) | ( n7052 & n10615 ) ;
  assign n10617 = n10615 | n10616 ;
  assign n10618 = ( ~n6752 & n7037 ) | ( ~n6752 & n10615 ) | ( n7037 & n10615 ) ;
  assign n10619 = n10617 | n10618 ;
  assign n10620 = n7035 & ~n9943 ;
  assign n10621 = n10619 | n10620 ;
  assign n10622 = n10621 ^ x26 ^ 1'b0 ;
  assign n10623 = ( n9648 & n9755 ) | ( n9648 & n10622 ) | ( n9755 & n10622 ) ;
  assign n10624 = n10622 ^ n9755 ^ n9648 ;
  assign n10625 = n6823 & n7190 ;
  assign n10626 = ( n6751 & n7188 ) | ( n6751 & n10625 ) | ( n7188 & n10625 ) ;
  assign n10627 = n10625 | n10626 ;
  assign n10628 = ( ~n6752 & n7192 ) | ( ~n6752 & n10625 ) | ( n7192 & n10625 ) ;
  assign n10629 = n10627 | n10628 ;
  assign n10630 = n7196 & ~n10013 ;
  assign n10631 = n10629 | n10630 ;
  assign n10632 = n10631 ^ x23 ^ 1'b0 ;
  assign n10633 = ( n9862 & ~n10566 ) | ( n9862 & n10632 ) | ( ~n10566 & n10632 ) ;
  assign n10634 = n10632 ^ n10566 ^ n9862 ;
  assign n10635 = n6791 & n6823 ;
  assign n10636 = ( ~n6752 & n6788 ) | ( ~n6752 & n10635 ) | ( n6788 & n10635 ) ;
  assign n10637 = n10635 | n10636 ;
  assign n10638 = ( n6747 & n6790 ) | ( n6747 & n10635 ) | ( n6790 & n10635 ) ;
  assign n10639 = n10637 | n10638 ;
  assign n10640 = n6823 & n6901 ;
  assign n10641 = ( n6747 & n6906 ) | ( n6747 & n10640 ) | ( n6906 & n10640 ) ;
  assign n10642 = n10640 | n10641 ;
  assign n10643 = ( ~n6752 & n6907 ) | ( ~n6752 & n10640 ) | ( n6907 & n10640 ) ;
  assign n10644 = n10642 | n10643 ;
  assign n10645 = n6918 & ~n9943 ;
  assign n10646 = n10644 & ~n10645 ;
  assign n10647 = n10646 ^ n10645 ^ x29 ;
  assign n10648 = ~n6004 & n7339 ;
  assign n10649 = n6789 & ~n9943 ;
  assign n10650 = n10639 | n10649 ;
  assign n10651 = ( ~n6707 & n7337 ) | ( ~n6707 & n10648 ) | ( n7337 & n10648 ) ;
  assign n10652 = n10648 | n10651 ;
  assign n10653 = ( ~n6477 & n7338 ) | ( ~n6477 & n10648 ) | ( n7338 & n10648 ) ;
  assign n10654 = n10652 | n10653 ;
  assign n10655 = n7340 & ~n10200 ;
  assign n10656 = n10654 | n10655 ;
  assign n10657 = ( ~n9774 & n10570 ) | ( ~n9774 & n10647 ) | ( n10570 & n10647 ) ;
  assign n10658 = n10647 ^ n10570 ^ n9774 ;
  assign n10659 = n7487 & ~n10241 ;
  assign n10660 = n10656 ^ x20 ^ 1'b0 ;
  assign n10661 = ( n10522 & ~n10634 ) | ( n10522 & n10660 ) | ( ~n10634 & n10660 ) ;
  assign n10662 = n10660 ^ n10634 ^ n10522 ;
  assign n10663 = ( n10577 & n10589 ) | ( n10577 & n10657 ) | ( n10589 & n10657 ) ;
  assign n10664 = n7493 & ~n9912 ;
  assign n10665 = n10657 ^ n10589 ^ n10577 ;
  assign n10666 = ~n10659 & n10664 ;
  assign n10667 = n10666 ^ n10659 ^ x17 ;
  assign n10668 = n10667 ^ n10662 ^ n10551 ;
  assign n10669 = n10668 ^ n10554 ^ n10552 ;
  assign n10670 = ( n10552 & n10554 ) | ( n10552 & ~n10668 ) | ( n10554 & ~n10668 ) ;
  assign n10671 = ( n10551 & ~n10662 ) | ( n10551 & n10667 ) | ( ~n10662 & n10667 ) ;
  assign n10672 = n6751 & n7192 ;
  assign n10673 = ( ~n6763 & n10581 ) | ( ~n6763 & n10650 ) | ( n10581 & n10650 ) ;
  assign n10674 = ( ~n6477 & n7188 ) | ( ~n6477 & n10672 ) | ( n7188 & n10672 ) ;
  assign n10675 = n10672 | n10674 ;
  assign n10676 = ( ~n6752 & n7190 ) | ( ~n6752 & n10672 ) | ( n7190 & n10672 ) ;
  assign n10677 = n10675 | n10676 ;
  assign n10678 = n7196 & ~n10135 ;
  assign n10679 = n10677 | n10678 ;
  assign n10680 = n10679 ^ x23 ^ 1'b0 ;
  assign n10681 = ( n10578 & n10633 ) | ( n10578 & n10680 ) | ( n10633 & n10680 ) ;
  assign n10682 = n10680 ^ n10633 ^ n10578 ;
  assign n10683 = n6751 & n6906 ;
  assign n10684 = ( ~n6477 & n6901 ) | ( ~n6477 & n10683 ) | ( n6901 & n10683 ) ;
  assign n10685 = n10683 | n10684 ;
  assign n10686 = ( ~n6004 & n6907 ) | ( ~n6004 & n10683 ) | ( n6907 & n10683 ) ;
  assign n10687 = n10596 ^ x29 ^ 1'b0 ;
  assign n10688 = n10685 | n10686 ;
  assign n10689 = n6918 & ~n10168 ;
  assign n10690 = ( n6918 & n10688 ) | ( n6918 & ~n10689 ) | ( n10688 & ~n10689 ) ;
  assign n10691 = n10581 ^ n6763 ^ 1'b0 ;
  assign n10692 = n10691 ^ n10650 ^ 1'b0 ;
  assign n10693 = ~n6707 & n7339 ;
  assign n10694 = ( n7337 & ~n9912 ) | ( n7337 & n10693 ) | ( ~n9912 & n10693 ) ;
  assign n10695 = n10693 | n10694 ;
  assign n10696 = ( ~n6004 & n7338 ) | ( ~n6004 & n10693 ) | ( n7338 & n10693 ) ;
  assign n10697 = n10695 | n10696 ;
  assign n10698 = ( n7340 & ~n10213 ) | ( n7340 & n10697 ) | ( ~n10213 & n10697 ) ;
  assign n10699 = n10697 | n10698 ;
  assign n10700 = n10699 ^ x20 ^ 1'b0 ;
  assign n10701 = ( n10661 & n10682 ) | ( n10661 & n10700 ) | ( n10682 & n10700 ) ;
  assign n10702 = n10700 ^ n10682 ^ n10661 ;
  assign n10703 = n6823 & n7052 ;
  assign n10704 = ( n6751 & n7037 ) | ( n6751 & n10703 ) | ( n7037 & n10703 ) ;
  assign n10705 = n10703 | n10704 ;
  assign n10706 = ( ~n6752 & n7036 ) | ( ~n6752 & n10703 ) | ( n7036 & n10703 ) ;
  assign n10707 = n10705 | n10706 ;
  assign n10708 = n7035 & ~n10013 ;
  assign n10709 = n10707 | n10708 ;
  assign n10710 = ( n10670 & n10671 ) | ( n10670 & n10702 ) | ( n10671 & n10702 ) ;
  assign n10711 = n10702 ^ n10671 ^ n10670 ;
  assign n10712 = n10709 ^ x26 ^ 1'b0 ;
  assign n10713 = n6823 & n6906 ;
  assign n10714 = ( n6751 & n6907 ) | ( n6751 & n10713 ) | ( n6907 & n10713 ) ;
  assign n10715 = n10713 | n10714 ;
  assign n10716 = ( ~n6752 & n6901 ) | ( ~n6752 & n10713 ) | ( n6901 & n10713 ) ;
  assign n10717 = n10715 | n10716 ;
  assign n10718 = ( n6918 & ~n10013 ) | ( n6918 & n10717 ) | ( ~n10013 & n10717 ) ;
  assign n10719 = n10717 | n10718 ;
  assign n10720 = ( ~n9683 & n10687 ) | ( ~n9683 & n10712 ) | ( n10687 & n10712 ) ;
  assign n10721 = n10712 ^ n10687 ^ n9683 ;
  assign n10722 = n10690 ^ x29 ^ 1'b0 ;
  assign n10723 = ( n10606 & n10692 ) | ( n10606 & ~n10722 ) | ( n10692 & ~n10722 ) ;
  assign n10724 = n10722 ^ n10692 ^ n10606 ;
  assign n10725 = n6789 & ~n10013 ;
  assign n10726 = ~n6752 & n6791 ;
  assign n10727 = ( n6790 & n6823 ) | ( n6790 & n10726 ) | ( n6823 & n10726 ) ;
  assign n10728 = ( n6751 & n6788 ) | ( n6751 & n10726 ) | ( n6788 & n10726 ) ;
  assign n10729 = n10726 | n10728 ;
  assign n10730 = n10727 | n10729 ;
  assign n10731 = n10725 | n10730 ;
  assign n10732 = ( n6364 & ~n6763 ) | ( n6364 & n10731 ) | ( ~n6763 & n10731 ) ;
  assign n10733 = n10731 ^ n6763 ^ n6364 ;
  assign n10734 = n10733 ^ n10723 ^ n10673 ;
  assign n10735 = ( ~n10673 & n10723 ) | ( ~n10673 & n10733 ) | ( n10723 & n10733 ) ;
  assign n10736 = n6751 & n7036 ;
  assign n10737 = ( ~n6477 & n7037 ) | ( ~n6477 & n10736 ) | ( n7037 & n10736 ) ;
  assign n10738 = n10736 | n10737 ;
  assign n10739 = ( ~n6752 & n7052 ) | ( ~n6752 & n10736 ) | ( n7052 & n10736 ) ;
  assign n10740 = n10738 | n10739 ;
  assign n10741 = ( n7035 & ~n10135 ) | ( n7035 & n10740 ) | ( ~n10135 & n10740 ) ;
  assign n10742 = n10740 | n10741 ;
  assign n10743 = n10742 ^ x26 ^ 1'b0 ;
  assign n10744 = n10743 ^ n10720 ^ n10613 ;
  assign n10745 = ( n10613 & n10720 ) | ( n10613 & n10743 ) | ( n10720 & n10743 ) ;
  assign n10746 = n6751 & n7052 ;
  assign n10747 = ( ~n6004 & n7037 ) | ( ~n6004 & n10746 ) | ( n7037 & n10746 ) ;
  assign n10748 = n10746 | n10747 ;
  assign n10749 = ( ~n6477 & n7036 ) | ( ~n6477 & n10746 ) | ( n7036 & n10746 ) ;
  assign n10750 = n10748 | n10749 ;
  assign n10751 = n7035 & n10168 ;
  assign n10752 = n10750 | n10751 ;
  assign n10753 = n10752 ^ x26 ^ 1'b0 ;
  assign n10754 = ( n10614 & ~n10658 ) | ( n10614 & n10753 ) | ( ~n10658 & n10753 ) ;
  assign n10755 = n10753 ^ n10658 ^ n10614 ;
  assign n10756 = n6751 & n6791 ;
  assign n10757 = ( ~n6477 & n6788 ) | ( ~n6477 & n10756 ) | ( n6788 & n10756 ) ;
  assign n10758 = n10756 | n10757 ;
  assign n10759 = ( ~n6752 & n6790 ) | ( ~n6752 & n10756 ) | ( n6790 & n10756 ) ;
  assign n10760 = n10758 | n10759 ;
  assign n10761 = n6763 ^ n6042 ^ x26 ;
  assign n10762 = ( ~x26 & n6042 ) | ( ~x26 & n6763 ) | ( n6042 & n6763 ) ;
  assign n10763 = n6751 & n6901 ;
  assign n10764 = ( ~n6752 & n6906 ) | ( ~n6752 & n10763 ) | ( n6906 & n10763 ) ;
  assign n10765 = n10763 | n10764 ;
  assign n10766 = ( ~n6477 & n6907 ) | ( ~n6477 & n10763 ) | ( n6907 & n10763 ) ;
  assign n10767 = n10765 | n10766 ;
  assign n10768 = n6918 & ~n10135 ;
  assign n10769 = n10767 | n10768 ;
  assign n10770 = n6789 & ~n10168 ;
  assign n10771 = n6789 & ~n10135 ;
  assign n10772 = n10760 | n10771 ;
  assign n10773 = n10772 ^ n10761 ^ n10732 ;
  assign n10774 = ( n10732 & ~n10761 ) | ( n10732 & n10772 ) | ( ~n10761 & n10772 ) ;
  assign n10775 = n6751 & n7190 ;
  assign n10776 = ( ~n6004 & n7188 ) | ( ~n6004 & n10775 ) | ( n7188 & n10775 ) ;
  assign n10777 = n10769 ^ x29 ^ 1'b0 ;
  assign n10778 = n10775 | n10776 ;
  assign n10779 = ( ~n6477 & n7192 ) | ( ~n6477 & n10775 ) | ( n7192 & n10775 ) ;
  assign n10780 = n10778 | n10779 ;
  assign n10781 = n7196 & n10168 ;
  assign n10782 = n10780 | n10781 ;
  assign n10783 = n10782 ^ x23 ^ 1'b0 ;
  assign n10784 = ( n10579 & n10624 ) | ( n10579 & n10783 ) | ( n10624 & n10783 ) ;
  assign n10785 = n10777 ^ n10663 ^ n10607 ;
  assign n10786 = ( n10607 & n10663 ) | ( n10607 & n10777 ) | ( n10663 & n10777 ) ;
  assign n10787 = ~n6477 & n6791 ;
  assign n10788 = ( ~n6004 & n6788 ) | ( ~n6004 & n10787 ) | ( n6788 & n10787 ) ;
  assign n10789 = n10787 | n10788 ;
  assign n10790 = ( n6751 & n6790 ) | ( n6751 & n10787 ) | ( n6790 & n10787 ) ;
  assign n10791 = n10789 | n10790 ;
  assign n10792 = ( n6789 & ~n10770 ) | ( n6789 & n10791 ) | ( ~n10770 & n10791 ) ;
  assign n10793 = n10783 ^ n10624 ^ n10579 ;
  assign n10794 = ~n6707 & n7037 ;
  assign n10795 = ( ~n6004 & n7036 ) | ( ~n6004 & n10794 ) | ( n7036 & n10794 ) ;
  assign n10796 = n10794 | n10795 ;
  assign n10797 = ( ~n6477 & n7052 ) | ( ~n6477 & n10794 ) | ( n7052 & n10794 ) ;
  assign n10798 = n10796 | n10797 ;
  assign n10799 = n7035 & ~n10200 ;
  assign n10800 = n10798 | n10799 ;
  assign n10801 = n10800 ^ x26 ^ 1'b0 ;
  assign n10802 = n10719 ^ x29 ^ 1'b0 ;
  assign n10803 = n10802 ^ n10801 ^ n10665 ;
  assign n10804 = ( n10665 & n10801 ) | ( n10665 & n10802 ) | ( n10801 & n10802 ) ;
  assign n10805 = ~n6707 & n7188 ;
  assign n10806 = ( ~n6477 & n7190 ) | ( ~n6477 & n10805 ) | ( n7190 & n10805 ) ;
  assign n10807 = n10805 | n10806 ;
  assign n10808 = ( ~n6004 & n7192 ) | ( ~n6004 & n10805 ) | ( n7192 & n10805 ) ;
  assign n10809 = n10807 | n10808 ;
  assign n10810 = n7196 & ~n10200 ;
  assign n10811 = n10809 | n10810 ;
  assign n10812 = n10811 ^ x23 ^ 1'b0 ;
  assign n10813 = ( n10623 & ~n10721 ) | ( n10623 & n10812 ) | ( ~n10721 & n10812 ) ;
  assign n10814 = n10812 ^ n10721 ^ n10623 ;
  assign n10815 = n7338 & ~n9912 ;
  assign n10816 = n7340 & ~n10241 ;
  assign n10817 = n10815 & ~n10816 ;
  assign n10818 = n10817 ^ n10816 ^ x20 ;
  assign n10819 = ( n10784 & ~n10814 ) | ( n10784 & n10818 ) | ( ~n10814 & n10818 ) ;
  assign n10820 = n10818 ^ n10814 ^ n10784 ;
  assign n10821 = n7190 & ~n9912 ;
  assign n10822 = n7196 & ~n10241 ;
  assign n10823 = n10821 & ~n10822 ;
  assign n10824 = n10823 ^ n10822 ^ x23 ;
  assign n10825 = n10824 ^ n10803 ^ n10754 ;
  assign n10826 = ( n10754 & n10803 ) | ( n10754 & n10824 ) | ( n10803 & n10824 ) ;
  assign n10827 = ~n6004 & n6791 ;
  assign n10828 = ( ~n6707 & n6788 ) | ( ~n6707 & n10827 ) | ( n6788 & n10827 ) ;
  assign n10829 = n10827 | n10828 ;
  assign n10830 = ( ~n6477 & n6790 ) | ( ~n6477 & n10827 ) | ( n6790 & n10827 ) ;
  assign n10831 = n10829 | n10830 ;
  assign n10832 = n6789 & ~n10200 ;
  assign n10833 = n10831 | n10832 ;
  assign n10834 = ~n6004 & n6901 ;
  assign n10835 = ( ~n6477 & n6906 ) | ( ~n6477 & n10834 ) | ( n6906 & n10834 ) ;
  assign n10836 = n10834 | n10835 ;
  assign n10837 = ( ~n6707 & n6907 ) | ( ~n6707 & n10834 ) | ( n6907 & n10834 ) ;
  assign n10838 = n10836 | n10837 ;
  assign n10839 = n10200 & ~n10838 ;
  assign n10840 = ( n6918 & n10838 ) | ( n6918 & ~n10839 ) | ( n10838 & ~n10839 ) ;
  assign n10841 = n7052 & ~n9912 ;
  assign n10842 = ( n7035 & ~n10241 ) | ( n7035 & n10841 ) | ( ~n10241 & n10841 ) ;
  assign n10843 = n10840 ^ x29 ^ 1'b0 ;
  assign n10844 = n10841 | n10842 ;
  assign n10845 = n10844 ^ x26 ^ 1'b0 ;
  assign n10846 = n10845 ^ n10843 ^ n10734 ;
  assign n10847 = ( n10734 & n10843 ) | ( n10734 & n10845 ) | ( n10843 & n10845 ) ;
  assign n10848 = n7037 & ~n9912 ;
  assign n10849 = ( ~n6707 & n7036 ) | ( ~n6707 & n10848 ) | ( n7036 & n10848 ) ;
  assign n10850 = n10848 | n10849 ;
  assign n10851 = ( ~n6004 & n7052 ) | ( ~n6004 & n10848 ) | ( n7052 & n10848 ) ;
  assign n10852 = n10850 | n10851 ;
  assign n10853 = ( n7035 & ~n10213 ) | ( n7035 & n10852 ) | ( ~n10213 & n10852 ) ;
  assign n10854 = n10852 | n10853 ;
  assign n10855 = n10854 ^ x26 ^ 1'b0 ;
  assign n10856 = ( n10785 & n10804 ) | ( n10785 & n10855 ) | ( n10804 & n10855 ) ;
  assign n10857 = n10855 ^ n10804 ^ n10785 ;
  assign n10858 = n7188 & ~n9912 ;
  assign n10859 = ( ~n6004 & n7190 ) | ( ~n6004 & n10858 ) | ( n7190 & n10858 ) ;
  assign n10860 = n10858 | n10859 ;
  assign n10861 = ( ~n6707 & n7192 ) | ( ~n6707 & n10858 ) | ( n7192 & n10858 ) ;
  assign n10862 = n10860 | n10861 ;
  assign n10863 = ( n7196 & ~n10213 ) | ( n7196 & n10862 ) | ( ~n10213 & n10862 ) ;
  assign n10864 = n10862 | n10863 ;
  assign n10865 = n10864 ^ x23 ^ 1'b0 ;
  assign n10866 = ( n10744 & n10813 ) | ( n10744 & n10865 ) | ( n10813 & n10865 ) ;
  assign n10867 = n10865 ^ n10813 ^ n10744 ;
  assign n10868 = ~n6707 & n6901 ;
  assign n10869 = ( ~n6004 & n6906 ) | ( ~n6004 & n10868 ) | ( n6906 & n10868 ) ;
  assign n10870 = n10868 | n10869 ;
  assign n10871 = ( n6907 & ~n9912 ) | ( n6907 & n10868 ) | ( ~n9912 & n10868 ) ;
  assign n10872 = n10870 | n10871 ;
  assign n10873 = n10792 ^ n10762 ^ n6675 ;
  assign n10874 = ( n6675 & n10762 ) | ( n6675 & n10792 ) | ( n10762 & n10792 ) ;
  assign n10875 = n6918 & ~n10213 ;
  assign n10876 = n10872 | n10875 ;
  assign n10877 = n10876 ^ x29 ^ 1'b0 ;
  assign n10878 = ( n10735 & n10773 ) | ( n10735 & ~n10877 ) | ( n10773 & ~n10877 ) ;
  assign n10879 = n10877 ^ n10773 ^ n10735 ;
  assign n10880 = n6918 & n10251 ;
  assign n10881 = n10874 ^ n6765 ^ n6675 ;
  assign n10882 = ( ~n6675 & n6765 ) | ( ~n6675 & n10874 ) | ( n6765 & n10874 ) ;
  assign n10883 = ( x29 & n6765 ) | ( x29 & ~n6767 ) | ( n6765 & ~n6767 ) ;
  assign n10884 = n6789 & ~n10213 ;
  assign n10885 = ( ~n6004 & n6790 ) | ( ~n6004 & n10884 ) | ( n6790 & n10884 ) ;
  assign n10886 = n6767 ^ n6765 ^ x29 ;
  assign n10887 = ( ~n6707 & n6791 ) | ( ~n6707 & n10884 ) | ( n6791 & n10884 ) ;
  assign n10888 = n10884 | n10887 ;
  assign n10889 = ( n6901 & ~n9912 ) | ( n6901 & n10880 ) | ( ~n9912 & n10880 ) ;
  assign n10890 = n10885 | n10888 ;
  assign n10891 = ( ~n6707 & n6906 ) | ( ~n6707 & n10880 ) | ( n6906 & n10880 ) ;
  assign n10892 = n10880 | n10889 ;
  assign n10893 = n10891 | n10892 ;
  assign n10894 = ( n10882 & n10886 ) | ( n10882 & n10890 ) | ( n10886 & n10890 ) ;
  assign n10895 = n10890 ^ n10886 ^ n10882 ;
  assign n10896 = n10893 ^ x29 ^ 1'b0 ;
  assign n10897 = ( n10774 & n10873 ) | ( n10774 & n10896 ) | ( n10873 & n10896 ) ;
  assign n10898 = n10896 ^ n10873 ^ n10774 ;
  assign n10899 = n7340 & n10251 ;
  assign n10900 = ( n7339 & ~n9912 ) | ( n7339 & n10899 ) | ( ~n9912 & n10899 ) ;
  assign n10901 = n10899 | n10900 ;
  assign n10902 = ( ~n6707 & n7338 ) | ( ~n6707 & n10899 ) | ( n7338 & n10899 ) ;
  assign n10903 = n10901 | n10902 ;
  assign n10904 = n10903 ^ x20 ^ 1'b0 ;
  assign n10905 = ( n10681 & n10793 ) | ( n10681 & n10904 ) | ( n10793 & n10904 ) ;
  assign n10906 = n10904 ^ n10793 ^ n10681 ;
  assign n10907 = n6906 & ~n9912 ;
  assign n10908 = n10907 ^ x29 ^ 1'b0 ;
  assign n10909 = n10906 ^ n10710 ^ n10701 ;
  assign n10910 = ( n10701 & n10710 ) | ( n10701 & n10906 ) | ( n10710 & n10906 ) ;
  assign n10911 = n7036 & ~n9912 ;
  assign n10912 = n10908 ^ n10881 ^ n10833 ;
  assign n10913 = ( n10833 & ~n10881 ) | ( n10833 & n10908 ) | ( ~n10881 & n10908 ) ;
  assign n10914 = ~n6707 & n7190 ;
  assign n10915 = n6789 & n10251 ;
  assign n10916 = ( ~n6707 & n7052 ) | ( ~n6707 & n10911 ) | ( n7052 & n10911 ) ;
  assign n10917 = n10911 | n10916 ;
  assign n10918 = ( n7035 & n10251 ) | ( n7035 & n10911 ) | ( n10251 & n10911 ) ;
  assign n10919 = ( n7196 & n10251 ) | ( n7196 & n10914 ) | ( n10251 & n10914 ) ;
  assign n10920 = n10914 | n10919 ;
  assign n10921 = ( n7192 & ~n9912 ) | ( n7192 & n10914 ) | ( ~n9912 & n10914 ) ;
  assign n10922 = ( n6791 & ~n9912 ) | ( n6791 & n10915 ) | ( ~n9912 & n10915 ) ;
  assign n10923 = n10917 | n10918 ;
  assign n10924 = ( ~n10820 & n10905 ) | ( ~n10820 & n10910 ) | ( n10905 & n10910 ) ;
  assign n10925 = n10920 | n10921 ;
  assign n10926 = n10924 ^ n10867 ^ n10819 ;
  assign n10927 = n10915 | n10922 ;
  assign n10928 = n6709 ^ n6432 ^ 1'b0 ;
  assign n10929 = n6432 & n6709 ;
  assign n10930 = n10910 ^ n10905 ^ n10820 ;
  assign n10931 = n10927 ^ n10883 ^ n6432 ;
  assign n10932 = n10923 ^ x26 ^ 1'b0 ;
  assign n10933 = ( n10819 & n10867 ) | ( n10819 & n10924 ) | ( n10867 & n10924 ) ;
  assign n10934 = n10925 ^ x23 ^ 1'b0 ;
  assign n10935 = n10934 ^ n10755 ^ n10745 ;
  assign n10936 = ( n10866 & n10933 ) | ( n10866 & ~n10935 ) | ( n10933 & ~n10935 ) ;
  assign n10937 = n6432 & ~n6725 ;
  assign n10938 = n10935 ^ n10933 ^ n10866 ;
  assign n10939 = ( n6432 & ~n10883 ) | ( n6432 & n10927 ) | ( ~n10883 & n10927 ) ;
  assign n10940 = ( n10745 & ~n10755 ) | ( n10745 & n10934 ) | ( ~n10755 & n10934 ) ;
  assign n10941 = ( n10825 & n10936 ) | ( n10825 & n10940 ) | ( n10936 & n10940 ) ;
  assign n10942 = ( n10826 & n10857 ) | ( n10826 & n10941 ) | ( n10857 & n10941 ) ;
  assign n10943 = n10932 ^ n10786 ^ n10724 ;
  assign n10944 = n10941 ^ n10857 ^ n10826 ;
  assign n10945 = ( n10856 & n10942 ) | ( n10856 & n10943 ) | ( n10942 & n10943 ) ;
  assign n10946 = ( n10724 & n10786 ) | ( n10724 & n10932 ) | ( n10786 & n10932 ) ;
  assign n10947 = ( n10846 & n10945 ) | ( n10846 & n10946 ) | ( n10945 & n10946 ) ;
  assign n10948 = ( n10847 & n10879 ) | ( n10847 & n10947 ) | ( n10879 & n10947 ) ;
  assign n10949 = ( ~n10878 & n10898 ) | ( ~n10878 & n10948 ) | ( n10898 & n10948 ) ;
  assign n10950 = ( n10897 & ~n10912 ) | ( n10897 & n10949 ) | ( ~n10912 & n10949 ) ;
  assign n10951 = n10950 ^ n10913 ^ n10895 ;
  assign n10952 = n10943 ^ n10942 ^ n10856 ;
  assign n10953 = n6725 ^ n6432 ^ 1'b0 ;
  assign n10954 = n10948 ^ n10898 ^ n10878 ;
  assign n10955 = ( n10895 & n10913 ) | ( n10895 & n10950 ) | ( n10913 & n10950 ) ;
  assign n10956 = n10955 ^ n10931 ^ n10894 ;
  assign n10957 = n10947 ^ n10879 ^ n10847 ;
  assign n10958 = n10937 ^ n10928 ^ 1'b0 ;
  assign n10959 = n10949 ^ n10912 ^ n10897 ;
  assign n10960 = ( n10894 & ~n10931 ) | ( n10894 & n10955 ) | ( ~n10931 & n10955 ) ;
  assign n10961 = ( n10939 & ~n10953 ) | ( n10939 & n10960 ) | ( ~n10953 & n10960 ) ;
  assign n10962 = ( ~n10928 & n10937 ) | ( ~n10928 & n10961 ) | ( n10937 & n10961 ) ;
  assign n10963 = ( n6320 & ~n10929 ) | ( n6320 & n10962 ) | ( ~n10929 & n10962 ) ;
  assign n10964 = n10940 ^ n10936 ^ n10825 ;
  assign n10965 = n10946 ^ n10945 ^ n10846 ;
  assign n10966 = n10929 ^ n6320 ^ 1'b0 ;
  assign n10967 = n10961 ^ n10958 ^ 1'b0 ;
  assign n10968 = n10960 ^ n10953 ^ n10939 ;
  assign n10969 = n10966 ^ n10962 ^ 1'b0 ;
  assign n10970 = ( x2 & ~n8090 ) | ( x2 & n10196 ) | ( ~n8090 & n10196 ) ;
  assign n10971 = ( x2 & ~n8113 ) | ( x2 & n10146 ) | ( ~n8113 & n10146 ) ;
  assign n10972 = ( n10146 & n10196 ) | ( n10146 & ~n10205 ) | ( n10196 & ~n10205 ) ;
  assign n10973 = n10196 ^ n10146 ^ 1'b0 ;
  assign n10974 = n6789 & n10973 ;
  assign n10975 = x2 & n10970 ;
  assign n10976 = n10971 & n10975 ;
  assign n10977 = ( n6788 & ~n10196 ) | ( n6788 & n10974 ) | ( ~n10196 & n10974 ) ;
  assign n10978 = n10146 & ~n10196 ;
  assign n10979 = n10978 ^ n10205 ^ 1'b0 ;
  assign n10980 = n10196 | n10972 ;
  assign n10981 = ( n6791 & ~n10146 ) | ( n6791 & n10974 ) | ( ~n10146 & n10974 ) ;
  assign n10982 = n10974 | n10981 ;
  assign n10983 = n8120 & n10973 ;
  assign n10984 = n10977 | n10982 ;
  assign n10985 = n10980 ^ n10233 ^ n10205 ;
  assign n10986 = n8120 & n10979 ;
  assign n10987 = n8086 & ~n10146 ;
  assign n10988 = ( n10976 & n10983 ) | ( n10976 & ~n10986 ) | ( n10983 & ~n10986 ) ;
  assign n10989 = ~n10983 & n10988 ;
  assign n10990 = ( n8088 & ~n10196 ) | ( n8088 & n10987 ) | ( ~n10196 & n10987 ) ;
  assign n10991 = n10987 | n10990 ;
  assign n10992 = ( n8090 & n10205 ) | ( n8090 & n10987 ) | ( n10205 & n10987 ) ;
  assign n10993 = n10991 | n10992 ;
  assign n10994 = ( x2 & n10986 ) | ( x2 & n10993 ) | ( n10986 & n10993 ) ;
  assign n10995 = n6789 & n10985 ;
  assign n10996 = x0 & ~n10146 ;
  assign n10997 = ( n10989 & n10994 ) | ( n10989 & ~n10996 ) | ( n10994 & ~n10996 ) ;
  assign n10998 = n6791 & ~n10196 ;
  assign n10999 = ~n10994 & n10997 ;
  assign n11000 = ( n6788 & n10205 ) | ( n6788 & n10998 ) | ( n10205 & n10998 ) ;
  assign n11001 = n10998 | n11000 ;
  assign n11002 = ( n6790 & ~n10146 ) | ( n6790 & n10998 ) | ( ~n10146 & n10998 ) ;
  assign n11003 = n11001 | n11002 ;
  assign n11004 = n6789 & ~n10979 ;
  assign n11005 = ( n6789 & n11003 ) | ( n6789 & ~n11004 ) | ( n11003 & ~n11004 ) ;
  assign n11006 = n10984 ^ n6671 ^ 1'b0 ;
  assign n11007 = ~n6671 & n10984 ;
  assign n11008 = ( ~n6712 & n11005 ) | ( ~n6712 & n11007 ) | ( n11005 & n11007 ) ;
  assign n11009 = n11007 ^ n11005 ^ n6712 ;
  assign n11010 = ( n6790 & ~n10196 ) | ( n6790 & n10995 ) | ( ~n10196 & n10995 ) ;
  assign n11011 = ( n6791 & n10205 ) | ( n6791 & n10995 ) | ( n10205 & n10995 ) ;
  assign n11012 = n10995 | n11011 ;
  assign n11013 = n11010 | n11012 ;
  assign n11014 = n8086 & ~n10196 ;
  assign n11015 = ( n8088 & n10205 ) | ( n8088 & n11014 ) | ( n10205 & n11014 ) ;
  assign n11016 = n11014 | n11015 ;
  assign n11017 = ( n8090 & ~n10233 ) | ( n8090 & n11014 ) | ( ~n10233 & n11014 ) ;
  assign n11018 = n11016 | n11017 ;
  assign n11019 = n6788 & ~n10233 ;
  assign n11020 = n11013 | n11019 ;
  assign n11021 = ( n6547 & n11008 ) | ( n6547 & n11020 ) | ( n11008 & n11020 ) ;
  assign n11022 = n11020 ^ n11008 ^ n6547 ;
  assign n11023 = n8029 & ~n10196 ;
  assign n11024 = ( ~n10205 & n10233 ) | ( ~n10205 & n10980 ) | ( n10233 & n10980 ) ;
  assign n11025 = ( n8037 & ~n10146 ) | ( n8037 & n11023 ) | ( ~n10146 & n11023 ) ;
  assign n11026 = n11023 | n11025 ;
  assign n11027 = ( n8033 & n10205 ) | ( n8033 & n11026 ) | ( n10205 & n11026 ) ;
  assign n11028 = n11026 | n11027 ;
  assign n11029 = ( n8034 & n10979 ) | ( n8034 & n11026 ) | ( n10979 & n11026 ) ;
  assign n11030 = n11028 | n11029 ;
  assign n11031 = n11030 ^ x5 ^ 1'b0 ;
  assign n11032 = n8089 & n10985 ;
  assign n11033 = n11018 | n11032 ;
  assign n11034 = n11033 ^ x2 ^ 1'b0 ;
  assign n11035 = n8034 & n10973 ;
  assign n11036 = ( n8029 & ~n10146 ) | ( n8029 & n11035 ) | ( ~n10146 & n11035 ) ;
  assign n11037 = n11024 ^ n10261 ^ n10233 ;
  assign n11038 = n6789 & n11037 ;
  assign n11039 = ( n8033 & ~n10196 ) | ( n8033 & n11035 ) | ( ~n10196 & n11035 ) ;
  assign n11040 = n11035 | n11036 ;
  assign n11041 = n11039 | n11040 ;
  assign n11042 = n6788 & ~n10261 ;
  assign n11043 = ( n6791 & ~n10233 ) | ( n6791 & n11038 ) | ( ~n10233 & n11038 ) ;
  assign n11044 = n11038 | n11043 ;
  assign n11045 = ( n6790 & n10205 ) | ( n6790 & n11038 ) | ( n10205 & n11038 ) ;
  assign n11046 = n11041 ^ x5 ^ 1'b0 ;
  assign n11047 = n11044 | n11045 ;
  assign n11048 = ( n6788 & ~n11042 ) | ( n6788 & n11047 ) | ( ~n11042 & n11047 ) ;
  assign n11049 = n8086 & n10205 ;
  assign n11050 = ( n8088 & ~n10233 ) | ( n8088 & n11049 ) | ( ~n10233 & n11049 ) ;
  assign n11051 = n11049 | n11050 ;
  assign n11052 = ( n8090 & n10261 ) | ( n8090 & n11049 ) | ( n10261 & n11049 ) ;
  assign n11053 = n11051 | n11052 ;
  assign n11054 = ( n8089 & n11037 ) | ( n8089 & n11053 ) | ( n11037 & n11053 ) ;
  assign n11055 = n11053 | n11054 ;
  assign n11056 = n8025 & ~n10146 ;
  assign n11057 = ( n10999 & n11034 ) | ( n10999 & n11056 ) | ( n11034 & n11056 ) ;
  assign n11058 = ( ~n6428 & n11021 ) | ( ~n6428 & n11048 ) | ( n11021 & n11048 ) ;
  assign n11059 = n11048 ^ n11021 ^ n6428 ;
  assign n11060 = n6788 & ~n10283 ;
  assign n11061 = x5 & ~n11056 ;
  assign n11062 = n11046 & n11061 ;
  assign n11063 = n11055 ^ x2 ^ 1'b0 ;
  assign n11064 = ( n10233 & ~n10261 ) | ( n10233 & n11024 ) | ( ~n10261 & n11024 ) ;
  assign n11065 = n11061 ^ n11046 ^ 1'b0 ;
  assign n11066 = ( n10261 & n10283 ) | ( n10261 & ~n11064 ) | ( n10283 & ~n11064 ) ;
  assign n11067 = n11064 ^ n10283 ^ n10261 ;
  assign n11068 = ( n11057 & n11063 ) | ( n11057 & n11065 ) | ( n11063 & n11065 ) ;
  assign n11069 = n6789 & ~n11067 ;
  assign n11070 = ( n6791 & n10261 ) | ( n6791 & n11069 ) | ( n10261 & n11069 ) ;
  assign n11071 = n11069 | n11070 ;
  assign n11072 = ( n6790 & ~n10233 ) | ( n6790 & n11069 ) | ( ~n10233 & n11069 ) ;
  assign n11073 = n11071 | n11072 ;
  assign n11074 = ( n6788 & ~n11060 ) | ( n6788 & n11073 ) | ( ~n11060 & n11073 ) ;
  assign n11075 = n11074 ^ n11058 ^ n6677 ;
  assign n11076 = n8086 & ~n10233 ;
  assign n11077 = ( ~n6677 & n11058 ) | ( ~n6677 & n11074 ) | ( n11058 & n11074 ) ;
  assign n11078 = ( n8088 & n10261 ) | ( n8088 & n11076 ) | ( n10261 & n11076 ) ;
  assign n11079 = n11076 | n11078 ;
  assign n11080 = ( n8090 & n10283 ) | ( n8090 & n11076 ) | ( n10283 & n11076 ) ;
  assign n11081 = n8089 & ~n11067 ;
  assign n11082 = n11079 | n11080 ;
  assign n11083 = n11081 | n11082 ;
  assign n11084 = n11062 ^ n11031 ^ 1'b0 ;
  assign n11085 = n11083 ^ x2 ^ 1'b0 ;
  assign n11086 = ( n11068 & n11084 ) | ( n11068 & n11085 ) | ( n11084 & n11085 ) ;
  assign n11087 = n11066 ^ n10283 ^ n10282 ;
  assign n11088 = n6789 & n11087 ;
  assign n11089 = ( n6791 & n10283 ) | ( n6791 & n11088 ) | ( n10283 & n11088 ) ;
  assign n11090 = n11088 | n11089 ;
  assign n11091 = ( n6790 & n10261 ) | ( n6790 & n11088 ) | ( n10261 & n11088 ) ;
  assign n11092 = ( n10282 & n10283 ) | ( n10282 & n11066 ) | ( n10283 & n11066 ) ;
  assign n11093 = n11090 | n11091 ;
  assign n11094 = n11031 & n11062 ;
  assign n11095 = n6788 & ~n10282 ;
  assign n11096 = ( n6788 & n11093 ) | ( n6788 & ~n11095 ) | ( n11093 & ~n11095 ) ;
  assign n11097 = n11096 ^ n11077 ^ n6768 ;
  assign n11098 = n11092 ^ n10282 ^ n10278 ;
  assign n11099 = ( n6768 & n11077 ) | ( n6768 & n11096 ) | ( n11077 & n11096 ) ;
  assign n11100 = ( n10278 & n10282 ) | ( n10278 & n11092 ) | ( n10282 & n11092 ) ;
  assign n11101 = n6789 & n11098 ;
  assign n11102 = ( n6791 & n10282 ) | ( n6791 & n11101 ) | ( n10282 & n11101 ) ;
  assign n11103 = n11101 | n11102 ;
  assign n11104 = ( n6790 & n10283 ) | ( n6790 & n11101 ) | ( n10283 & n11101 ) ;
  assign n11105 = n11103 | n11104 ;
  assign n11106 = n6788 & ~n10278 ;
  assign n11107 = ( n6788 & n11105 ) | ( n6788 & ~n11106 ) | ( n11105 & ~n11106 ) ;
  assign n11108 = n11107 ^ n11099 ^ n6770 ;
  assign n11109 = ( n6770 & n11099 ) | ( n6770 & n11107 ) | ( n11099 & n11107 ) ;
  assign n11110 = n8086 & n10261 ;
  assign n11111 = n8029 & n10205 ;
  assign n11112 = ( n8088 & n10283 ) | ( n8088 & n11110 ) | ( n10283 & n11110 ) ;
  assign n11113 = n11110 | n11112 ;
  assign n11114 = ( n8089 & n11087 ) | ( n8089 & n11113 ) | ( n11087 & n11113 ) ;
  assign n11115 = ( n8090 & n10282 ) | ( n8090 & n11113 ) | ( n10282 & n11113 ) ;
  assign n11116 = n11113 | n11115 ;
  assign n11117 = n11114 | n11116 ;
  assign n11118 = ( n8033 & ~n10233 ) | ( n8033 & n11111 ) | ( ~n10233 & n11111 ) ;
  assign n11119 = ( n8037 & ~n10196 ) | ( n8037 & n11111 ) | ( ~n10196 & n11111 ) ;
  assign n11120 = n11111 | n11119 ;
  assign n11121 = n11118 | n11120 ;
  assign n11122 = n7927 & ~n10146 ;
  assign n11123 = n8034 & n10985 ;
  assign n11124 = n11121 | n11123 ;
  assign n11125 = n11124 ^ x5 ^ 1'b0 ;
  assign n11126 = n11125 ^ n11122 ^ n11094 ;
  assign n11127 = ( n11094 & n11122 ) | ( n11094 & n11125 ) | ( n11122 & n11125 ) ;
  assign n11128 = n7932 & ~n10146 ;
  assign n11129 = n11117 ^ x2 ^ 1'b0 ;
  assign n11130 = x8 & ~n11122 ;
  assign n11131 = ( n11086 & n11126 ) | ( n11086 & n11129 ) | ( n11126 & n11129 ) ;
  assign n11132 = ( n7930 & n10973 ) | ( n7930 & n11128 ) | ( n10973 & n11128 ) ;
  assign n11133 = ( n7929 & ~n10196 ) | ( n7929 & n11128 ) | ( ~n10196 & n11128 ) ;
  assign n11134 = n11128 | n11132 ;
  assign n11135 = n8029 & ~n10233 ;
  assign n11136 = n11133 | n11134 ;
  assign n11137 = ( n8037 & n10205 ) | ( n8037 & n11135 ) | ( n10205 & n11135 ) ;
  assign n11138 = n11135 | n11137 ;
  assign n11139 = ( n8033 & n10261 ) | ( n8033 & n11135 ) | ( n10261 & n11135 ) ;
  assign n11140 = n11136 ^ x8 ^ 1'b0 ;
  assign n11141 = n11138 | n11139 ;
  assign n11142 = ( n8034 & n11037 ) | ( n8034 & n11141 ) | ( n11037 & n11141 ) ;
  assign n11143 = n11141 | n11142 ;
  assign n11144 = n11140 ^ n11130 ^ 1'b0 ;
  assign n11145 = n11143 ^ x5 ^ 1'b0 ;
  assign n11146 = n11130 & n11140 ;
  assign n11147 = n11145 ^ n11144 ^ n11127 ;
  assign n11148 = ( n11127 & n11144 ) | ( n11127 & n11145 ) | ( n11144 & n11145 ) ;
  assign n11149 = n8086 & n10283 ;
  assign n11150 = ( n8088 & n10282 ) | ( n8088 & n11149 ) | ( n10282 & n11149 ) ;
  assign n11151 = n11149 | n11150 ;
  assign n11152 = ( n8090 & n10278 ) | ( n8090 & n11149 ) | ( n10278 & n11149 ) ;
  assign n11153 = n11151 | n11152 ;
  assign n11154 = n8089 & n11098 ;
  assign n11155 = n11153 | n11154 ;
  assign n11156 = n11155 ^ x2 ^ 1'b0 ;
  assign n11157 = ( n11131 & n11147 ) | ( n11131 & n11156 ) | ( n11147 & n11156 ) ;
  assign n11158 = n11100 ^ n10280 ^ n10278 ;
  assign n11159 = n6789 & ~n11158 ;
  assign n11160 = ( n6791 & n10278 ) | ( n6791 & n11159 ) | ( n10278 & n11159 ) ;
  assign n11161 = n11159 | n11160 ;
  assign n11162 = ( n6790 & n10282 ) | ( n6790 & n11159 ) | ( n10282 & n11159 ) ;
  assign n11163 = n6788 & ~n10280 ;
  assign n11164 = n11161 | n11162 ;
  assign n11165 = n11163 | n11164 ;
  assign n11166 = ( n6824 & n11109 ) | ( n6824 & n11165 ) | ( n11109 & n11165 ) ;
  assign n11167 = n11165 ^ n11109 ^ n6824 ;
  assign n11168 = n7932 & ~n10196 ;
  assign n11169 = ( n7943 & ~n10146 ) | ( n7943 & n11168 ) | ( ~n10146 & n11168 ) ;
  assign n11170 = n11168 | n11169 ;
  assign n11171 = ( n7929 & n10205 ) | ( n7929 & n11170 ) | ( n10205 & n11170 ) ;
  assign n11172 = n8029 & n10261 ;
  assign n11173 = n11170 | n11171 ;
  assign n11174 = ( n7930 & n10979 ) | ( n7930 & n11170 ) | ( n10979 & n11170 ) ;
  assign n11175 = n11173 | n11174 ;
  assign n11176 = n11175 ^ x8 ^ 1'b0 ;
  assign n11177 = n11176 ^ n11146 ^ 1'b0 ;
  assign n11178 = n11146 & n11176 ;
  assign n11179 = ( n8037 & ~n10233 ) | ( n8037 & n11172 ) | ( ~n10233 & n11172 ) ;
  assign n11180 = n11172 | n11179 ;
  assign n11181 = ( n8033 & n10283 ) | ( n8033 & n11172 ) | ( n10283 & n11172 ) ;
  assign n11182 = n11180 | n11181 ;
  assign n11183 = n8034 & ~n11067 ;
  assign n11184 = n11182 | n11183 ;
  assign n11185 = n11184 ^ x5 ^ 1'b0 ;
  assign n11186 = ( n11148 & n11177 ) | ( n11148 & n11185 ) | ( n11177 & n11185 ) ;
  assign n11187 = n11185 ^ n11177 ^ n11148 ;
  assign n11188 = n8086 & n10282 ;
  assign n11189 = ( n10278 & ~n10280 ) | ( n10278 & n11100 ) | ( ~n10280 & n11100 ) ;
  assign n11190 = ( n8088 & n10278 ) | ( n8088 & n11188 ) | ( n10278 & n11188 ) ;
  assign n11191 = n11188 | n11190 ;
  assign n11192 = ( n8090 & ~n10280 ) | ( n8090 & n11188 ) | ( ~n10280 & n11188 ) ;
  assign n11193 = n11191 | n11192 ;
  assign n11194 = n8089 & ~n11158 ;
  assign n11195 = n11193 & ~n11194 ;
  assign n11196 = n11195 ^ n11194 ^ x2 ;
  assign n11197 = ( n11157 & n11187 ) | ( n11157 & n11196 ) | ( n11187 & n11196 ) ;
  assign n11198 = n8029 & n10283 ;
  assign n11199 = ( n8037 & n10261 ) | ( n8037 & n11198 ) | ( n10261 & n11198 ) ;
  assign n11200 = n11198 | n11199 ;
  assign n11201 = ( n8033 & n10282 ) | ( n8033 & n11200 ) | ( n10282 & n11200 ) ;
  assign n11202 = n11200 | n11201 ;
  assign n11203 = ( n8034 & n11087 ) | ( n8034 & n11200 ) | ( n11087 & n11200 ) ;
  assign n11204 = n8086 & n10278 ;
  assign n11205 = ( n8090 & n10306 ) | ( n8090 & n11204 ) | ( n10306 & n11204 ) ;
  assign n11206 = ( n8088 & ~n10280 ) | ( n8088 & n11204 ) | ( ~n10280 & n11204 ) ;
  assign n11207 = n11204 | n11206 ;
  assign n11208 = n11205 | n11207 ;
  assign n11209 = n7932 & n10205 ;
  assign n11210 = n7930 & n10985 ;
  assign n11211 = n11202 | n11203 ;
  assign n11212 = n11211 ^ x5 ^ 1'b0 ;
  assign n11213 = ( n7943 & ~n10196 ) | ( n7943 & n11209 ) | ( ~n10196 & n11209 ) ;
  assign n11214 = n11209 | n11213 ;
  assign n11215 = ( n7929 & ~n10233 ) | ( n7929 & n11209 ) | ( ~n10233 & n11209 ) ;
  assign n11216 = n11214 | n11215 ;
  assign n11217 = n11210 | n11216 ;
  assign n11218 = n11217 ^ x8 ^ 1'b0 ;
  assign n11219 = n7827 & ~n10146 ;
  assign n11220 = n11219 ^ n11218 ^ n11178 ;
  assign n11221 = ( n11186 & n11212 ) | ( n11186 & n11220 ) | ( n11212 & n11220 ) ;
  assign n11222 = n11220 ^ n11212 ^ n11186 ;
  assign n11223 = n11189 ^ n10306 ^ n10280 ;
  assign n11224 = n8089 & ~n11223 ;
  assign n11225 = n11208 & ~n11224 ;
  assign n11226 = n11225 ^ n11224 ^ x2 ;
  assign n11227 = ( ~n10280 & n10306 ) | ( ~n10280 & n11189 ) | ( n10306 & n11189 ) ;
  assign n11228 = n7932 & ~n10233 ;
  assign n11229 = ( n11178 & n11218 ) | ( n11178 & n11219 ) | ( n11218 & n11219 ) ;
  assign n11230 = ( n11197 & n11222 ) | ( n11197 & n11226 ) | ( n11222 & n11226 ) ;
  assign n11231 = n7829 & ~n10146 ;
  assign n11232 = ( n7834 & ~n10196 ) | ( n7834 & n11231 ) | ( ~n10196 & n11231 ) ;
  assign n11233 = ( n7838 & n10973 ) | ( n7838 & n11231 ) | ( n10973 & n11231 ) ;
  assign n11234 = n11231 | n11233 ;
  assign n11235 = ( n7929 & n10261 ) | ( n7929 & n11228 ) | ( n10261 & n11228 ) ;
  assign n11236 = n11232 | n11234 ;
  assign n11237 = n11236 ^ x11 ^ 1'b0 ;
  assign n11238 = x11 & ~n11219 ;
  assign n11239 = ( n7943 & n10205 ) | ( n7943 & n11228 ) | ( n10205 & n11228 ) ;
  assign n11240 = n11228 | n11239 ;
  assign n11241 = n11235 | n11240 ;
  assign n11242 = ( n7930 & n11037 ) | ( n7930 & n11241 ) | ( n11037 & n11241 ) ;
  assign n11243 = n11241 | n11242 ;
  assign n11244 = n11243 ^ x8 ^ 1'b0 ;
  assign n11245 = n8029 & n10282 ;
  assign n11246 = ( n8037 & n10283 ) | ( n8037 & n11245 ) | ( n10283 & n11245 ) ;
  assign n11247 = n11245 | n11246 ;
  assign n11248 = ( n8033 & n10278 ) | ( n8033 & n11245 ) | ( n10278 & n11245 ) ;
  assign n11249 = n11247 | n11248 ;
  assign n11250 = n11238 ^ n11237 ^ 1'b0 ;
  assign n11251 = n11237 & n11238 ;
  assign n11252 = n11250 ^ n11244 ^ n11229 ;
  assign n11253 = ( n11229 & n11244 ) | ( n11229 & n11250 ) | ( n11244 & n11250 ) ;
  assign n11254 = n8034 & n11098 ;
  assign n11255 = n11249 | n11254 ;
  assign n11256 = n8086 & ~n10280 ;
  assign n11257 = ( n8088 & n10306 ) | ( n8088 & n11256 ) | ( n10306 & n11256 ) ;
  assign n11258 = n11256 | n11257 ;
  assign n11259 = ( n8090 & ~n10340 ) | ( n8090 & n11256 ) | ( ~n10340 & n11256 ) ;
  assign n11260 = n11255 ^ x5 ^ 1'b0 ;
  assign n11261 = n11258 | n11259 ;
  assign n11262 = ( n11221 & n11252 ) | ( n11221 & n11260 ) | ( n11252 & n11260 ) ;
  assign n11263 = n11260 ^ n11252 ^ n11221 ;
  assign n11264 = n11227 ^ n10340 ^ n10306 ;
  assign n11265 = ( n10306 & ~n10340 ) | ( n10306 & n11227 ) | ( ~n10340 & n11227 ) ;
  assign n11266 = n8089 & ~n11264 ;
  assign n11267 = n11261 & ~n11266 ;
  assign n11268 = n11267 ^ n11266 ^ x2 ;
  assign n11269 = ( n11230 & n11263 ) | ( n11230 & n11268 ) | ( n11263 & n11268 ) ;
  assign n11270 = n7829 & ~n10196 ;
  assign n11271 = ( n7833 & ~n10146 ) | ( n7833 & n11270 ) | ( ~n10146 & n11270 ) ;
  assign n11272 = n11270 | n11271 ;
  assign n11273 = n6789 & ~n11223 ;
  assign n11274 = ( n7834 & n10205 ) | ( n7834 & n11272 ) | ( n10205 & n11272 ) ;
  assign n11275 = ( n6791 & ~n10280 ) | ( n6791 & n11273 ) | ( ~n10280 & n11273 ) ;
  assign n11276 = n11273 | n11275 ;
  assign n11277 = ( n6790 & n10278 ) | ( n6790 & n11273 ) | ( n10278 & n11273 ) ;
  assign n11278 = n11272 | n11274 ;
  assign n11279 = ( n7838 & n10979 ) | ( n7838 & n11272 ) | ( n10979 & n11272 ) ;
  assign n11280 = n11276 | n11277 ;
  assign n11281 = n6788 & ~n10306 ;
  assign n11282 = ( n6788 & n11280 ) | ( n6788 & ~n11281 ) | ( n11280 & ~n11281 ) ;
  assign n11283 = n11282 ^ n11166 ^ n6773 ;
  assign n11284 = ( n6773 & n11166 ) | ( n6773 & n11282 ) | ( n11166 & n11282 ) ;
  assign n11285 = n7932 & n10261 ;
  assign n11286 = n11278 | n11279 ;
  assign n11287 = ( n7943 & ~n10233 ) | ( n7943 & n11285 ) | ( ~n10233 & n11285 ) ;
  assign n11288 = n11285 | n11287 ;
  assign n11289 = ( n7929 & n10283 ) | ( n7929 & n11285 ) | ( n10283 & n11285 ) ;
  assign n11290 = n11288 | n11289 ;
  assign n11291 = n7930 & ~n11067 ;
  assign n11292 = n11286 ^ x11 ^ 1'b0 ;
  assign n11293 = n11290 | n11291 ;
  assign n11294 = n8029 & n10278 ;
  assign n11295 = ( n8037 & n10282 ) | ( n8037 & n11294 ) | ( n10282 & n11294 ) ;
  assign n11296 = n11294 | n11295 ;
  assign n11297 = ( n8033 & ~n10280 ) | ( n8033 & n11294 ) | ( ~n10280 & n11294 ) ;
  assign n11298 = n11296 | n11297 ;
  assign n11299 = n11292 ^ n11251 ^ 1'b0 ;
  assign n11300 = n11251 & n11292 ;
  assign n11301 = n11293 ^ x8 ^ 1'b0 ;
  assign n11302 = n11301 ^ n11299 ^ n11253 ;
  assign n11303 = ( n11253 & n11299 ) | ( n11253 & n11301 ) | ( n11299 & n11301 ) ;
  assign n11304 = n8086 & n10306 ;
  assign n11305 = ( n8088 & ~n10340 ) | ( n8088 & n11304 ) | ( ~n10340 & n11304 ) ;
  assign n11306 = n11304 | n11305 ;
  assign n11307 = ( n8090 & n10353 ) | ( n8090 & n11304 ) | ( n10353 & n11304 ) ;
  assign n11308 = n11306 | n11307 ;
  assign n11309 = n8034 & ~n11158 ;
  assign n11310 = n11298 & ~n11309 ;
  assign n11311 = n11310 ^ n11309 ^ x5 ;
  assign n11312 = n11311 ^ n11302 ^ n11262 ;
  assign n11313 = ( n11262 & n11302 ) | ( n11262 & n11311 ) | ( n11302 & n11311 ) ;
  assign n11314 = n11265 ^ n10353 ^ n10340 ;
  assign n11315 = ( ~n10340 & n10353 ) | ( ~n10340 & n11265 ) | ( n10353 & n11265 ) ;
  assign n11316 = n8089 & ~n11314 ;
  assign n11317 = n11308 | n11316 ;
  assign n11318 = n6789 & ~n11264 ;
  assign n11319 = n11317 ^ x2 ^ 1'b0 ;
  assign n11320 = ( n11269 & n11312 ) | ( n11269 & n11319 ) | ( n11312 & n11319 ) ;
  assign n11321 = ( n6791 & n10306 ) | ( n6791 & n11318 ) | ( n10306 & n11318 ) ;
  assign n11322 = n11318 | n11321 ;
  assign n11323 = n6788 & ~n10340 ;
  assign n11324 = ( n6790 & ~n10280 ) | ( n6790 & n11318 ) | ( ~n10280 & n11318 ) ;
  assign n11325 = n11322 | n11324 ;
  assign n11326 = n11323 | n11325 ;
  assign n11327 = n11326 ^ n11284 ^ n6703 ;
  assign n11328 = ( n6703 & n11284 ) | ( n6703 & n11326 ) | ( n11284 & n11326 ) ;
  assign n11329 = n7663 & ~n10146 ;
  assign n11330 = n7838 & n10985 ;
  assign n11331 = n7829 & n10205 ;
  assign n11332 = ( n7833 & ~n10196 ) | ( n7833 & n11331 ) | ( ~n10196 & n11331 ) ;
  assign n11333 = n11331 | n11332 ;
  assign n11334 = ( n7834 & ~n10233 ) | ( n7834 & n11331 ) | ( ~n10233 & n11331 ) ;
  assign n11335 = n11333 | n11334 ;
  assign n11336 = n7932 & n10283 ;
  assign n11337 = ( n7943 & n10261 ) | ( n7943 & n11336 ) | ( n10261 & n11336 ) ;
  assign n11338 = n11336 | n11337 ;
  assign n11339 = ( n7929 & n10282 ) | ( n7929 & n11338 ) | ( n10282 & n11338 ) ;
  assign n11340 = n11338 | n11339 ;
  assign n11341 = ( n7930 & n11087 ) | ( n7930 & n11338 ) | ( n11087 & n11338 ) ;
  assign n11342 = n11340 | n11341 ;
  assign n11343 = n11342 ^ x8 ^ 1'b0 ;
  assign n11344 = n11330 | n11335 ;
  assign n11345 = n11344 ^ x11 ^ 1'b0 ;
  assign n11346 = n11345 ^ n11329 ^ n11300 ;
  assign n11347 = ( n11303 & n11343 ) | ( n11303 & n11346 ) | ( n11343 & n11346 ) ;
  assign n11348 = n11346 ^ n11343 ^ n11303 ;
  assign n11349 = n8029 & ~n10280 ;
  assign n11350 = ( n8037 & n10278 ) | ( n8037 & n11349 ) | ( n10278 & n11349 ) ;
  assign n11351 = n11349 | n11350 ;
  assign n11352 = ( n8033 & n10306 ) | ( n8033 & n11349 ) | ( n10306 & n11349 ) ;
  assign n11353 = n11351 | n11352 ;
  assign n11354 = n8034 & ~n11223 ;
  assign n11355 = n11353 & ~n11354 ;
  assign n11356 = n11355 ^ n11354 ^ x5 ;
  assign n11357 = n11356 ^ n11348 ^ n11313 ;
  assign n11358 = ( n11313 & n11348 ) | ( n11313 & n11356 ) | ( n11348 & n11356 ) ;
  assign n11359 = ( n11300 & n11329 ) | ( n11300 & n11345 ) | ( n11329 & n11345 ) ;
  assign n11360 = n8086 & ~n10340 ;
  assign n11361 = ( n8090 & n10372 ) | ( n8090 & n11360 ) | ( n10372 & n11360 ) ;
  assign n11362 = ( n8088 & n10353 ) | ( n8088 & n11360 ) | ( n10353 & n11360 ) ;
  assign n11363 = n11360 | n11362 ;
  assign n11364 = n11361 | n11363 ;
  assign n11365 = n11315 ^ n10372 ^ n10353 ;
  assign n11366 = n8089 & n11365 ;
  assign n11367 = n11364 | n11366 ;
  assign n11368 = n11367 ^ x2 ^ 1'b0 ;
  assign n11369 = ( n11320 & n11357 ) | ( n11320 & n11368 ) | ( n11357 & n11368 ) ;
  assign n11370 = n7829 & ~n10233 ;
  assign n11371 = ( n7833 & n10205 ) | ( n7833 & n11370 ) | ( n10205 & n11370 ) ;
  assign n11372 = n11370 | n11371 ;
  assign n11373 = ( n7834 & n10261 ) | ( n7834 & n11370 ) | ( n10261 & n11370 ) ;
  assign n11374 = n11372 | n11373 ;
  assign n11375 = n7669 & ~n10146 ;
  assign n11376 = ( n7838 & n11037 ) | ( n7838 & n11374 ) | ( n11037 & n11374 ) ;
  assign n11377 = n11374 | n11376 ;
  assign n11378 = ( n7666 & n10973 ) | ( n7666 & n11375 ) | ( n10973 & n11375 ) ;
  assign n11379 = n11375 | n11378 ;
  assign n11380 = n11377 ^ x11 ^ 1'b0 ;
  assign n11381 = ( n7667 & ~n10196 ) | ( n7667 & n11375 ) | ( ~n10196 & n11375 ) ;
  assign n11382 = n11379 | n11381 ;
  assign n11383 = x14 & ~n11329 ;
  assign n11384 = n11382 ^ x14 ^ 1'b0 ;
  assign n11385 = n11383 & n11384 ;
  assign n11386 = n11384 ^ n11383 ^ 1'b0 ;
  assign n11387 = n11386 ^ n11380 ^ n11359 ;
  assign n11388 = ( n11359 & n11380 ) | ( n11359 & n11386 ) | ( n11380 & n11386 ) ;
  assign n11389 = n7932 & n10282 ;
  assign n11390 = ( n7943 & n10283 ) | ( n7943 & n11389 ) | ( n10283 & n11389 ) ;
  assign n11391 = n11389 | n11390 ;
  assign n11392 = ( n7929 & n10278 ) | ( n7929 & n11389 ) | ( n10278 & n11389 ) ;
  assign n11393 = n11391 | n11392 ;
  assign n11394 = n7930 & n11098 ;
  assign n11395 = n11393 | n11394 ;
  assign n11396 = n11395 ^ x8 ^ 1'b0 ;
  assign n11397 = n11396 ^ n11387 ^ n11347 ;
  assign n11398 = ( n11347 & n11387 ) | ( n11347 & n11396 ) | ( n11387 & n11396 ) ;
  assign n11399 = n8029 & n10306 ;
  assign n11400 = ( n8037 & ~n10280 ) | ( n8037 & n11399 ) | ( ~n10280 & n11399 ) ;
  assign n11401 = n11399 | n11400 ;
  assign n11402 = ( n8033 & ~n10340 ) | ( n8033 & n11399 ) | ( ~n10340 & n11399 ) ;
  assign n11403 = n11401 | n11402 ;
  assign n11404 = n8034 & ~n11264 ;
  assign n11405 = n11403 & ~n11404 ;
  assign n11406 = n11405 ^ n11404 ^ x5 ;
  assign n11407 = ( n11358 & n11397 ) | ( n11358 & n11406 ) | ( n11397 & n11406 ) ;
  assign n11408 = n11406 ^ n11397 ^ n11358 ;
  assign n11409 = n7829 & n10261 ;
  assign n11410 = n7838 & ~n11067 ;
  assign n11411 = ( n7833 & ~n10233 ) | ( n7833 & n11409 ) | ( ~n10233 & n11409 ) ;
  assign n11412 = n11409 | n11411 ;
  assign n11413 = ( n7834 & n10283 ) | ( n7834 & n11409 ) | ( n10283 & n11409 ) ;
  assign n11414 = n11412 | n11413 ;
  assign n11415 = n11410 | n11414 ;
  assign n11416 = n7669 & ~n10196 ;
  assign n11417 = ( n7674 & ~n10146 ) | ( n7674 & n11416 ) | ( ~n10146 & n11416 ) ;
  assign n11418 = n11416 | n11417 ;
  assign n11419 = n11415 ^ x11 ^ 1'b0 ;
  assign n11420 = ( n7667 & n10205 ) | ( n7667 & n11418 ) | ( n10205 & n11418 ) ;
  assign n11421 = n11418 | n11420 ;
  assign n11422 = ( n7666 & n10979 ) | ( n7666 & n11418 ) | ( n10979 & n11418 ) ;
  assign n11423 = n11421 | n11422 ;
  assign n11424 = n11423 ^ x14 ^ 1'b0 ;
  assign n11425 = n11385 & n11424 ;
  assign n11426 = n11424 ^ n11385 ^ 1'b0 ;
  assign n11427 = ( n11388 & n11419 ) | ( n11388 & n11426 ) | ( n11419 & n11426 ) ;
  assign n11428 = n11426 ^ n11419 ^ n11388 ;
  assign n11429 = n7932 & n10278 ;
  assign n11430 = ( n7943 & n10282 ) | ( n7943 & n11429 ) | ( n10282 & n11429 ) ;
  assign n11431 = n11429 | n11430 ;
  assign n11432 = ( n7929 & ~n10280 ) | ( n7929 & n11429 ) | ( ~n10280 & n11429 ) ;
  assign n11433 = n11431 | n11432 ;
  assign n11434 = n7930 & ~n11158 ;
  assign n11435 = n11433 & ~n11434 ;
  assign n11436 = n11435 ^ n11434 ^ x8 ;
  assign n11437 = ( n11398 & n11428 ) | ( n11398 & n11436 ) | ( n11428 & n11436 ) ;
  assign n11438 = n11436 ^ n11428 ^ n11398 ;
  assign n11439 = n8029 & ~n10340 ;
  assign n11440 = ( n8037 & n10306 ) | ( n8037 & n11439 ) | ( n10306 & n11439 ) ;
  assign n11441 = n11439 | n11440 ;
  assign n11442 = ( n8033 & n10353 ) | ( n8033 & n11439 ) | ( n10353 & n11439 ) ;
  assign n11443 = n11441 | n11442 ;
  assign n11444 = n8034 & ~n11314 ;
  assign n11445 = n11443 | n11444 ;
  assign n11446 = n11445 ^ x5 ^ 1'b0 ;
  assign n11447 = ( n11407 & n11438 ) | ( n11407 & n11446 ) | ( n11438 & n11446 ) ;
  assign n11448 = n11446 ^ n11438 ^ n11407 ;
  assign n11449 = n7829 & n10283 ;
  assign n11450 = ( n7833 & n10261 ) | ( n7833 & n11449 ) | ( n10261 & n11449 ) ;
  assign n11451 = n11449 | n11450 ;
  assign n11452 = ( n7838 & n11087 ) | ( n7838 & n11451 ) | ( n11087 & n11451 ) ;
  assign n11453 = n7669 & n10205 ;
  assign n11454 = ( n7834 & n10282 ) | ( n7834 & n11451 ) | ( n10282 & n11451 ) ;
  assign n11455 = n11451 | n11454 ;
  assign n11456 = ( n7674 & ~n10196 ) | ( n7674 & n11453 ) | ( ~n10196 & n11453 ) ;
  assign n11457 = n11452 | n11455 ;
  assign n11458 = ( n7667 & ~n10233 ) | ( n7667 & n11453 ) | ( ~n10233 & n11453 ) ;
  assign n11459 = n11453 | n11456 ;
  assign n11460 = n7666 & n10985 ;
  assign n11461 = n11458 | n11459 ;
  assign n11462 = n7483 & ~n10146 ;
  assign n11463 = n11460 | n11461 ;
  assign n11464 = n11463 ^ x14 ^ 1'b0 ;
  assign n11465 = ( n11425 & n11462 ) | ( n11425 & n11464 ) | ( n11462 & n11464 ) ;
  assign n11466 = n11464 ^ n11462 ^ n11425 ;
  assign n11467 = n11457 ^ x11 ^ 1'b0 ;
  assign n11468 = x17 & ~n11462 ;
  assign n11469 = ( n11427 & n11466 ) | ( n11427 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11470 = n11467 ^ n11466 ^ n11427 ;
  assign n11471 = n7932 & ~n10280 ;
  assign n11472 = ( n7943 & n10278 ) | ( n7943 & n11471 ) | ( n10278 & n11471 ) ;
  assign n11473 = n11471 | n11472 ;
  assign n11474 = ( n7929 & n10306 ) | ( n7929 & n11471 ) | ( n10306 & n11471 ) ;
  assign n11475 = n11473 | n11474 ;
  assign n11476 = n7930 & ~n11223 ;
  assign n11477 = n11475 & ~n11476 ;
  assign n11478 = n11477 ^ n11476 ^ x8 ;
  assign n11479 = ( n11437 & n11470 ) | ( n11437 & n11478 ) | ( n11470 & n11478 ) ;
  assign n11480 = n11478 ^ n11470 ^ n11437 ;
  assign n11481 = n8029 & n10353 ;
  assign n11482 = ( n8037 & ~n10340 ) | ( n8037 & n11481 ) | ( ~n10340 & n11481 ) ;
  assign n11483 = n11481 | n11482 ;
  assign n11484 = ( n8033 & n10372 ) | ( n8033 & n11481 ) | ( n10372 & n11481 ) ;
  assign n11485 = n11483 | n11484 ;
  assign n11486 = n8034 & n11365 ;
  assign n11487 = n11485 | n11486 ;
  assign n11488 = n11487 ^ x5 ^ 1'b0 ;
  assign n11489 = n11488 ^ n11480 ^ n11447 ;
  assign n11490 = ( n11447 & n11480 ) | ( n11447 & n11488 ) | ( n11480 & n11488 ) ;
  assign n11491 = n7669 & ~n10233 ;
  assign n11492 = n7485 & ~n10146 ;
  assign n11493 = ( n7674 & n10205 ) | ( n7674 & n11491 ) | ( n10205 & n11491 ) ;
  assign n11494 = n7669 & n10261 ;
  assign n11495 = ( n7486 & ~n10196 ) | ( n7486 & n11492 ) | ( ~n10196 & n11492 ) ;
  assign n11496 = n11491 | n11493 ;
  assign n11497 = ( n7667 & n10283 ) | ( n7667 & n11494 ) | ( n10283 & n11494 ) ;
  assign n11498 = ( n7487 & n10973 ) | ( n7487 & n11492 ) | ( n10973 & n11492 ) ;
  assign n11499 = ( n7667 & n10261 ) | ( n7667 & n11491 ) | ( n10261 & n11491 ) ;
  assign n11500 = n11496 | n11499 ;
  assign n11501 = n11492 | n11498 ;
  assign n11502 = ( n7674 & ~n10233 ) | ( n7674 & n11494 ) | ( ~n10233 & n11494 ) ;
  assign n11503 = n7669 & n10283 ;
  assign n11504 = n11494 | n11502 ;
  assign n11505 = n11495 | n11501 ;
  assign n11506 = ( n7666 & n11037 ) | ( n7666 & n11500 ) | ( n11037 & n11500 ) ;
  assign n11507 = n11505 ^ x17 ^ 1'b0 ;
  assign n11508 = n11500 | n11506 ;
  assign n11509 = n11508 ^ x14 ^ 1'b0 ;
  assign n11510 = n11507 ^ n11468 ^ 1'b0 ;
  assign n11511 = ( n7674 & n10261 ) | ( n7674 & n11503 ) | ( n10261 & n11503 ) ;
  assign n11512 = n11497 | n11504 ;
  assign n11513 = ( n11465 & n11509 ) | ( n11465 & n11510 ) | ( n11509 & n11510 ) ;
  assign n11514 = n11503 | n11511 ;
  assign n11515 = n11468 & n11507 ;
  assign n11516 = ( n7667 & n10282 ) | ( n7667 & n11514 ) | ( n10282 & n11514 ) ;
  assign n11517 = ( n7666 & n11087 ) | ( n7666 & n11514 ) | ( n11087 & n11514 ) ;
  assign n11518 = n11514 | n11516 ;
  assign n11519 = n11517 | n11518 ;
  assign n11520 = n7485 & ~n10196 ;
  assign n11521 = ( n7493 & ~n10146 ) | ( n7493 & n11520 ) | ( ~n10146 & n11520 ) ;
  assign n11522 = n11520 | n11521 ;
  assign n11523 = ( n7486 & n10205 ) | ( n7486 & n11522 ) | ( n10205 & n11522 ) ;
  assign n11524 = n11522 | n11523 ;
  assign n11525 = ( n7487 & n10979 ) | ( n7487 & n11522 ) | ( n10979 & n11522 ) ;
  assign n11526 = n11524 | n11525 ;
  assign n11527 = n11526 ^ x17 ^ 1'b0 ;
  assign n11528 = n11527 ^ n11515 ^ 1'b0 ;
  assign n11529 = n11510 ^ n11509 ^ n11465 ;
  assign n11530 = n11519 ^ x14 ^ 1'b0 ;
  assign n11531 = n7485 & n10205 ;
  assign n11532 = n11515 & n11527 ;
  assign n11533 = ( n7486 & ~n10233 ) | ( n7486 & n11531 ) | ( ~n10233 & n11531 ) ;
  assign n11534 = ( n7493 & ~n10196 ) | ( n7493 & n11531 ) | ( ~n10196 & n11531 ) ;
  assign n11535 = n11531 | n11533 ;
  assign n11536 = n11534 | n11535 ;
  assign n11537 = n7487 & n10985 ;
  assign n11538 = n7666 & ~n11067 ;
  assign n11539 = n11536 | n11537 ;
  assign n11540 = n11512 | n11538 ;
  assign n11541 = n11540 ^ x14 ^ 1'b0 ;
  assign n11542 = n11541 ^ n11528 ^ n11513 ;
  assign n11543 = n11539 ^ x17 ^ 1'b0 ;
  assign n11544 = ( n11513 & n11528 ) | ( n11513 & n11541 ) | ( n11528 & n11541 ) ;
  assign n11545 = n7333 & ~n10146 ;
  assign n11546 = n11545 ^ n11543 ^ n11532 ;
  assign n11547 = n11546 ^ n11544 ^ n11530 ;
  assign n11548 = ( n11532 & n11543 ) | ( n11532 & n11545 ) | ( n11543 & n11545 ) ;
  assign n11549 = n7485 & ~n10233 ;
  assign n11550 = ( n11530 & n11544 ) | ( n11530 & n11546 ) | ( n11544 & n11546 ) ;
  assign n11551 = ( n7486 & n10261 ) | ( n7486 & n11549 ) | ( n10261 & n11549 ) ;
  assign n11552 = n11549 | n11551 ;
  assign n11553 = ( n7493 & n10205 ) | ( n7493 & n11549 ) | ( n10205 & n11549 ) ;
  assign n11554 = n11552 | n11553 ;
  assign n11555 = x20 & ~n11545 ;
  assign n11556 = n7340 & n10973 ;
  assign n11557 = ( n7339 & ~n10146 ) | ( n7339 & n11556 ) | ( ~n10146 & n11556 ) ;
  assign n11558 = n11556 | n11557 ;
  assign n11559 = ( n7337 & ~n10196 ) | ( n7337 & n11556 ) | ( ~n10196 & n11556 ) ;
  assign n11560 = n11558 | n11559 ;
  assign n11561 = n11560 ^ x20 ^ 1'b0 ;
  assign n11562 = ( n7487 & n11037 ) | ( n7487 & n11554 ) | ( n11037 & n11554 ) ;
  assign n11563 = n11554 | n11562 ;
  assign n11564 = n11555 & n11561 ;
  assign n11565 = n11563 ^ x17 ^ 1'b0 ;
  assign n11566 = n11561 ^ n11555 ^ 1'b0 ;
  assign n11567 = n11566 ^ n11565 ^ n11548 ;
  assign n11568 = ( n11548 & n11565 ) | ( n11548 & n11566 ) | ( n11565 & n11566 ) ;
  assign n11569 = n7190 & ~n10146 ;
  assign n11570 = ( n7192 & ~n10196 ) | ( n7192 & n11569 ) | ( ~n10196 & n11569 ) ;
  assign n11571 = n11569 | n11570 ;
  assign n11572 = ( n7196 & n10979 ) | ( n7196 & n11571 ) | ( n10979 & n11571 ) ;
  assign n11573 = ( n7188 & n10205 ) | ( n7188 & n11571 ) | ( n10205 & n11571 ) ;
  assign n11574 = n11571 | n11573 ;
  assign n11575 = n7485 & n10261 ;
  assign n11576 = n7339 & ~n10196 ;
  assign n11577 = ( n7338 & ~n10146 ) | ( n7338 & n11576 ) | ( ~n10146 & n11576 ) ;
  assign n11578 = n11576 | n11577 ;
  assign n11579 = ( n7486 & n10283 ) | ( n7486 & n11575 ) | ( n10283 & n11575 ) ;
  assign n11580 = n11575 | n11579 ;
  assign n11581 = ( n7493 & ~n10233 ) | ( n7493 & n11575 ) | ( ~n10233 & n11575 ) ;
  assign n11582 = n11580 | n11581 ;
  assign n11583 = ( n7337 & n10205 ) | ( n7337 & n11578 ) | ( n10205 & n11578 ) ;
  assign n11584 = n11578 | n11583 ;
  assign n11585 = ( n7340 & n10979 ) | ( n7340 & n11578 ) | ( n10979 & n11578 ) ;
  assign n11586 = n11584 | n11585 ;
  assign n11587 = n7037 & n10205 ;
  assign n11588 = n11572 | n11574 ;
  assign n11589 = ( n7036 & ~n10196 ) | ( n7036 & n11587 ) | ( ~n10196 & n11587 ) ;
  assign n11590 = n11587 | n11589 ;
  assign n11591 = ( n7052 & ~n10146 ) | ( n7052 & n11587 ) | ( ~n10146 & n11587 ) ;
  assign n11592 = n11588 ^ x23 ^ 1'b0 ;
  assign n11593 = n11590 | n11591 ;
  assign n11594 = n7487 & ~n11067 ;
  assign n11595 = n11586 ^ x20 ^ 1'b0 ;
  assign n11596 = n11582 | n11594 ;
  assign n11597 = n11596 ^ x17 ^ 1'b0 ;
  assign n11598 = ~n7035 & n10979 ;
  assign n11599 = ( n10979 & n11593 ) | ( n10979 & ~n11598 ) | ( n11593 & ~n11598 ) ;
  assign n11600 = n11564 & n11595 ;
  assign n11601 = n11599 ^ x26 ^ 1'b0 ;
  assign n11602 = n11595 ^ n11564 ^ 1'b0 ;
  assign n11603 = n11602 ^ n11597 ^ n11568 ;
  assign n11604 = ( n11568 & n11597 ) | ( n11568 & n11602 ) | ( n11597 & n11602 ) ;
  assign n11605 = n6901 & ~n10196 ;
  assign n11606 = ( n6906 & ~n10146 ) | ( n6906 & n11605 ) | ( ~n10146 & n11605 ) ;
  assign n11607 = n11605 | n11606 ;
  assign n11608 = ( n6907 & n10205 ) | ( n6907 & n11607 ) | ( n10205 & n11607 ) ;
  assign n11609 = n11607 | n11608 ;
  assign n11610 = ( n6918 & n10979 ) | ( n6918 & n11607 ) | ( n10979 & n11607 ) ;
  assign n11611 = n11609 | n11610 ;
  assign n11612 = n7339 & n10205 ;
  assign n11613 = ( n7338 & ~n10196 ) | ( n7338 & n11612 ) | ( ~n10196 & n11612 ) ;
  assign n11614 = ( n7337 & ~n10233 ) | ( n7337 & n11612 ) | ( ~n10233 & n11612 ) ;
  assign n11615 = n11612 | n11614 ;
  assign n11616 = n7188 & ~n10196 ;
  assign n11617 = n11613 | n11615 ;
  assign n11618 = n7340 & n10985 ;
  assign n11619 = n11617 | n11618 ;
  assign n11620 = n7187 & ~n10146 ;
  assign n11621 = n11619 ^ x20 ^ 1'b0 ;
  assign n11622 = ( n7196 & n10973 ) | ( n7196 & n11616 ) | ( n10973 & n11616 ) ;
  assign n11623 = n11616 | n11622 ;
  assign n11624 = ( n11600 & n11620 ) | ( n11600 & n11621 ) | ( n11620 & n11621 ) ;
  assign n11625 = n11621 ^ n11620 ^ n11600 ;
  assign n11626 = x23 & ~n11620 ;
  assign n11627 = ( n7192 & ~n10146 ) | ( n7192 & n11616 ) | ( ~n10146 & n11616 ) ;
  assign n11628 = n7339 & ~n10233 ;
  assign n11629 = n11623 | n11627 ;
  assign n11630 = n11629 ^ x23 ^ 1'b0 ;
  assign n11631 = ( n7337 & n10261 ) | ( n7337 & n11628 ) | ( n10261 & n11628 ) ;
  assign n11632 = n11628 | n11631 ;
  assign n11633 = ( n7338 & n10205 ) | ( n7338 & n11628 ) | ( n10205 & n11628 ) ;
  assign n11634 = n11632 | n11633 ;
  assign n11635 = ( n7340 & n11037 ) | ( n7340 & n11634 ) | ( n11037 & n11634 ) ;
  assign n11636 = n11634 | n11635 ;
  assign n11637 = n11626 & n11630 ;
  assign n11638 = n11630 ^ n11626 ^ 1'b0 ;
  assign n11639 = n11636 ^ x20 ^ 1'b0 ;
  assign n11640 = ( n11624 & n11638 ) | ( n11624 & n11639 ) | ( n11638 & n11639 ) ;
  assign n11641 = n11639 ^ n11638 ^ n11624 ;
  assign n11642 = n7485 & n10283 ;
  assign n11643 = ( n7493 & n10261 ) | ( n7493 & n11642 ) | ( n10261 & n11642 ) ;
  assign n11644 = n11642 | n11643 ;
  assign n11645 = n11637 ^ n11592 ^ 1'b0 ;
  assign n11646 = n11592 & n11637 ;
  assign n11647 = ( n7486 & n10282 ) | ( n7486 & n11644 ) | ( n10282 & n11644 ) ;
  assign n11648 = n11644 | n11647 ;
  assign n11649 = ( n7487 & n11087 ) | ( n7487 & n11644 ) | ( n11087 & n11644 ) ;
  assign n11650 = n11648 | n11649 ;
  assign n11651 = n11650 ^ x17 ^ 1'b0 ;
  assign n11652 = n11651 ^ n11625 ^ n11604 ;
  assign n11653 = ( n11604 & n11625 ) | ( n11604 & n11651 ) | ( n11625 & n11651 ) ;
  assign n11654 = n7339 & n10261 ;
  assign n11655 = ( n7337 & n10283 ) | ( n7337 & n11654 ) | ( n10283 & n11654 ) ;
  assign n11656 = n11654 | n11655 ;
  assign n11657 = ( n7338 & ~n10233 ) | ( n7338 & n11654 ) | ( ~n10233 & n11654 ) ;
  assign n11658 = n11656 | n11657 ;
  assign n11659 = n7340 & ~n11067 ;
  assign n11660 = n11658 | n11659 ;
  assign n11661 = n11660 ^ x20 ^ 1'b0 ;
  assign n11662 = n11661 ^ n11645 ^ n11640 ;
  assign n11663 = ( n11640 & n11645 ) | ( n11640 & n11661 ) | ( n11645 & n11661 ) ;
  assign n11664 = n7037 & ~n10233 ;
  assign n11665 = n7188 & ~n10233 ;
  assign n11666 = ( n7190 & ~n10196 ) | ( n7190 & n11665 ) | ( ~n10196 & n11665 ) ;
  assign n11667 = n11665 | n11666 ;
  assign n11668 = ( n7036 & n10205 ) | ( n7036 & n11664 ) | ( n10205 & n11664 ) ;
  assign n11669 = n11664 | n11668 ;
  assign n11670 = ( n7192 & n10205 ) | ( n7192 & n11665 ) | ( n10205 & n11665 ) ;
  assign n11671 = n11667 | n11670 ;
  assign n11672 = ( n7052 & ~n10196 ) | ( n7052 & n11664 ) | ( ~n10196 & n11664 ) ;
  assign n11673 = n7037 & ~n10196 ;
  assign n11674 = ( n7036 & ~n10146 ) | ( n7036 & n11673 ) | ( ~n10146 & n11673 ) ;
  assign n11675 = n11673 | n11674 ;
  assign n11676 = ( n7035 & n10973 ) | ( n7035 & n11673 ) | ( n10973 & n11673 ) ;
  assign n11677 = n6918 & n10973 ;
  assign n11678 = n11669 | n11672 ;
  assign n11679 = ( n6901 & ~n10146 ) | ( n6901 & n11677 ) | ( ~n10146 & n11677 ) ;
  assign n11680 = n11677 | n11679 ;
  assign n11681 = ( n6907 & ~n10196 ) | ( n6907 & n11677 ) | ( ~n10196 & n11677 ) ;
  assign n11682 = n11680 | n11681 ;
  assign n11683 = n7035 & n10985 ;
  assign n11684 = n11678 | n11683 ;
  assign n11685 = n7196 & n10985 ;
  assign n11686 = n11684 ^ x26 ^ 1'b0 ;
  assign n11687 = n11671 | n11685 ;
  assign n11688 = n6901 & n10205 ;
  assign n11689 = ( n6906 & ~n10196 ) | ( n6906 & n11688 ) | ( ~n10196 & n11688 ) ;
  assign n11690 = n11688 | n11689 ;
  assign n11691 = n11675 | n11676 ;
  assign n11692 = ( n6907 & ~n10233 ) | ( n6907 & n11688 ) | ( ~n10233 & n11688 ) ;
  assign n11693 = n6787 & ~n10146 ;
  assign n11694 = n11690 | n11692 ;
  assign n11695 = n11687 ^ x23 ^ 1'b0 ;
  assign n11696 = n11691 ^ x26 ^ 1'b0 ;
  assign n11697 = n6898 & ~n10146 ;
  assign n11698 = n7030 & ~n10146 ;
  assign n11699 = n11611 ^ x29 ^ 1'b0 ;
  assign n11700 = n6918 & n10985 ;
  assign n11701 = n11682 ^ x29 ^ 1'b0 ;
  assign n11702 = n11694 | n11700 ;
  assign n11703 = n11702 ^ x29 ^ 1'b0 ;
  assign n11704 = n11698 ^ n11695 ^ n11646 ;
  assign n11705 = ( n11646 & n11695 ) | ( n11646 & n11698 ) | ( n11695 & n11698 ) ;
  assign n11706 = x26 & ~n11698 ;
  assign n11707 = n11706 ^ n11696 ^ 1'b0 ;
  assign n11708 = n11696 & n11706 ;
  assign n11709 = n11601 & n11708 ;
  assign n11710 = n11708 ^ n11601 ^ 1'b0 ;
  assign n11711 = ( n11686 & n11697 ) | ( n11686 & n11709 ) | ( n11697 & n11709 ) ;
  assign n11712 = n11709 ^ n11697 ^ n11686 ;
  assign n11713 = x29 & ~n11697 ;
  assign n11714 = n11713 ^ n11701 ^ 1'b0 ;
  assign n11715 = n11701 & n11713 ;
  assign n11716 = n11715 ^ n11699 ^ 1'b0 ;
  assign n11717 = n11699 & n11715 ;
  assign n11718 = ( n11693 & n11703 ) | ( n11693 & n11717 ) | ( n11703 & n11717 ) ;
  assign n11719 = n11717 ^ n11703 ^ n11693 ;
  assign n11720 = n6901 & ~n10233 ;
  assign n11721 = ( n6906 & n10205 ) | ( n6906 & n11720 ) | ( n10205 & n11720 ) ;
  assign n11722 = n11720 | n11721 ;
  assign n11723 = ( n6907 & n10261 ) | ( n6907 & n11720 ) | ( n10261 & n11720 ) ;
  assign n11724 = n11722 | n11723 ;
  assign n11725 = n6918 & n11037 ;
  assign n11726 = n11724 | n11725 ;
  assign n11727 = n11726 ^ x29 ^ 1'b0 ;
  assign n11728 = n11727 ^ n11718 ^ n11006 ;
  assign n11729 = ( ~n11006 & n11718 ) | ( ~n11006 & n11727 ) | ( n11718 & n11727 ) ;
  assign n11730 = n6901 & n10261 ;
  assign n11731 = ( n6906 & ~n10233 ) | ( n6906 & n11730 ) | ( ~n10233 & n11730 ) ;
  assign n11732 = n11730 | n11731 ;
  assign n11733 = ( n6907 & n10283 ) | ( n6907 & n11730 ) | ( n10283 & n11730 ) ;
  assign n11734 = n11732 | n11733 ;
  assign n11735 = n6918 & ~n11067 ;
  assign n11736 = n11734 | n11735 ;
  assign n11737 = n11736 ^ x29 ^ 1'b0 ;
  assign n11738 = ( ~n11009 & n11729 ) | ( ~n11009 & n11737 ) | ( n11729 & n11737 ) ;
  assign n11739 = n11737 ^ n11729 ^ n11009 ;
  assign n11740 = n7037 & n10261 ;
  assign n11741 = ( n7036 & ~n10233 ) | ( n7036 & n11740 ) | ( ~n10233 & n11740 ) ;
  assign n11742 = n11740 | n11741 ;
  assign n11743 = ( n7052 & n10205 ) | ( n7052 & n11740 ) | ( n10205 & n11740 ) ;
  assign n11744 = n11742 | n11743 ;
  assign n11745 = ( n7035 & n11037 ) | ( n7035 & n11744 ) | ( n11037 & n11744 ) ;
  assign n11746 = n11744 | n11745 ;
  assign n11747 = n11746 ^ x26 ^ 1'b0 ;
  assign n11748 = ( n11711 & n11714 ) | ( n11711 & n11747 ) | ( n11714 & n11747 ) ;
  assign n11749 = n11747 ^ n11714 ^ n11711 ;
  assign n11750 = n7196 & ~n11067 ;
  assign n11751 = n7188 & n10261 ;
  assign n11752 = ( n7190 & n10205 ) | ( n7190 & n11751 ) | ( n10205 & n11751 ) ;
  assign n11753 = n11751 | n11752 ;
  assign n11754 = ( n7192 & ~n10233 ) | ( n7192 & n11751 ) | ( ~n10233 & n11751 ) ;
  assign n11755 = n11753 | n11754 ;
  assign n11756 = n7037 & n10283 ;
  assign n11757 = ( n7196 & n11037 ) | ( n7196 & n11755 ) | ( n11037 & n11755 ) ;
  assign n11758 = n11755 | n11757 ;
  assign n11759 = n11758 ^ x23 ^ 1'b0 ;
  assign n11760 = n11759 ^ n11707 ^ n11705 ;
  assign n11761 = ( n11705 & n11707 ) | ( n11705 & n11759 ) | ( n11707 & n11759 ) ;
  assign n11762 = n7188 & n10283 ;
  assign n11763 = ( n7190 & ~n10233 ) | ( n7190 & n11762 ) | ( ~n10233 & n11762 ) ;
  assign n11764 = n11762 | n11763 ;
  assign n11765 = ( n7192 & n10261 ) | ( n7192 & n11762 ) | ( n10261 & n11762 ) ;
  assign n11766 = ( n7052 & ~n10233 ) | ( n7052 & n11756 ) | ( ~n10233 & n11756 ) ;
  assign n11767 = n11764 | n11765 ;
  assign n11768 = ( n7036 & n10261 ) | ( n7036 & n11756 ) | ( n10261 & n11756 ) ;
  assign n11769 = n11756 | n11768 ;
  assign n11770 = n11766 | n11769 ;
  assign n11771 = n11750 | n11767 ;
  assign n11772 = n7035 & ~n11067 ;
  assign n11773 = n11770 | n11772 ;
  assign n11774 = n11773 ^ x26 ^ 1'b0 ;
  assign n11775 = ( n11716 & n11748 ) | ( n11716 & n11774 ) | ( n11748 & n11774 ) ;
  assign n11776 = n11774 ^ n11748 ^ n11716 ;
  assign n11777 = n11771 ^ x23 ^ 1'b0 ;
  assign n11778 = ( n11710 & n11761 ) | ( n11710 & n11777 ) | ( n11761 & n11777 ) ;
  assign n11779 = n11777 ^ n11761 ^ n11710 ;
  assign n11780 = n7339 & n10283 ;
  assign n11781 = ( n7338 & n10261 ) | ( n7338 & n11780 ) | ( n10261 & n11780 ) ;
  assign n11782 = n11780 | n11781 ;
  assign n11783 = ( n7337 & n10282 ) | ( n7337 & n11782 ) | ( n10282 & n11782 ) ;
  assign n11784 = n11782 | n11783 ;
  assign n11785 = ( n7340 & n11087 ) | ( n7340 & n11782 ) | ( n11087 & n11782 ) ;
  assign n11786 = n11784 | n11785 ;
  assign n11787 = n11786 ^ x20 ^ 1'b0 ;
  assign n11788 = n11787 ^ n11704 ^ n11663 ;
  assign n11789 = ( n11663 & n11704 ) | ( n11663 & n11787 ) | ( n11704 & n11787 ) ;
  assign n11790 = n7190 & n10261 ;
  assign n11791 = ( n7192 & n10283 ) | ( n7192 & n11790 ) | ( n10283 & n11790 ) ;
  assign n11792 = n11790 | n11791 ;
  assign n11793 = ( n7188 & n10282 ) | ( n7188 & n11792 ) | ( n10282 & n11792 ) ;
  assign n11794 = n11792 | n11793 ;
  assign n11795 = ( n7196 & n11087 ) | ( n7196 & n11792 ) | ( n11087 & n11792 ) ;
  assign n11796 = n11794 | n11795 ;
  assign n11797 = n11796 ^ x23 ^ 1'b0 ;
  assign n11798 = ( n11712 & n11778 ) | ( n11712 & n11797 ) | ( n11778 & n11797 ) ;
  assign n11799 = n11797 ^ n11778 ^ n11712 ;
  assign n11800 = n7037 & n10282 ;
  assign n11801 = ( n7036 & n10283 ) | ( n7036 & n11800 ) | ( n10283 & n11800 ) ;
  assign n11802 = n11800 | n11801 ;
  assign n11803 = ( n7052 & n10261 ) | ( n7052 & n11800 ) | ( n10261 & n11800 ) ;
  assign n11804 = n11802 | n11803 ;
  assign n11805 = n7035 & n11087 ;
  assign n11806 = n11804 | n11805 ;
  assign n11807 = n11806 ^ x26 ^ 1'b0 ;
  assign n11808 = n11807 ^ n11775 ^ n11719 ;
  assign n11809 = ( n11719 & n11775 ) | ( n11719 & n11807 ) | ( n11775 & n11807 ) ;
  assign n11810 = n6901 & n10283 ;
  assign n11811 = ( n6906 & n10261 ) | ( n6906 & n11810 ) | ( n10261 & n11810 ) ;
  assign n11812 = n11810 | n11811 ;
  assign n11813 = ( n6907 & n10282 ) | ( n6907 & n11810 ) | ( n10282 & n11810 ) ;
  assign n11814 = n11812 | n11813 ;
  assign n11815 = n6918 & n11087 ;
  assign n11816 = n11814 | n11815 ;
  assign n11817 = n11816 ^ x29 ^ 1'b0 ;
  assign n11818 = ( n11022 & n11738 ) | ( n11022 & n11817 ) | ( n11738 & n11817 ) ;
  assign n11819 = n11817 ^ n11738 ^ n11022 ;
  assign n11820 = n7339 & n10282 ;
  assign n11821 = ( n7337 & n10278 ) | ( n7337 & n11820 ) | ( n10278 & n11820 ) ;
  assign n11822 = n11820 | n11821 ;
  assign n11823 = ( n7338 & n10283 ) | ( n7338 & n11820 ) | ( n10283 & n11820 ) ;
  assign n11824 = n11822 | n11823 ;
  assign n11825 = n7340 & n11098 ;
  assign n11826 = n11824 | n11825 ;
  assign n11827 = n11826 ^ x20 ^ 1'b0 ;
  assign n11828 = ( n11760 & n11789 ) | ( n11760 & n11827 ) | ( n11789 & n11827 ) ;
  assign n11829 = n11827 ^ n11789 ^ n11760 ;
  assign n11830 = n7339 & n10278 ;
  assign n11831 = ( n7337 & ~n10280 ) | ( n7337 & n11830 ) | ( ~n10280 & n11830 ) ;
  assign n11832 = n11830 | n11831 ;
  assign n11833 = ( n7338 & n10282 ) | ( n7338 & n11830 ) | ( n10282 & n11830 ) ;
  assign n11834 = n11832 | n11833 ;
  assign n11835 = n7340 & ~n11158 ;
  assign n11836 = n11834 & ~n11835 ;
  assign n11837 = n11836 ^ n11835 ^ x20 ;
  assign n11838 = n11837 ^ n11828 ^ n11779 ;
  assign n11839 = ( n11779 & n11828 ) | ( n11779 & n11837 ) | ( n11828 & n11837 ) ;
  assign n11840 = n7339 & ~n10280 ;
  assign n11841 = ( n7337 & n10306 ) | ( n7337 & n11840 ) | ( n10306 & n11840 ) ;
  assign n11842 = n11840 | n11841 ;
  assign n11843 = ( n7338 & n10278 ) | ( n7338 & n11840 ) | ( n10278 & n11840 ) ;
  assign n11844 = n11842 | n11843 ;
  assign n11845 = n7340 & ~n11223 ;
  assign n11846 = n11844 & ~n11845 ;
  assign n11847 = n11846 ^ n11845 ^ x20 ;
  assign n11848 = n11847 ^ n11839 ^ n11799 ;
  assign n11849 = ( n11799 & n11839 ) | ( n11799 & n11847 ) | ( n11839 & n11847 ) ;
  assign n11850 = n7188 & n10278 ;
  assign n11851 = ( n7190 & n10283 ) | ( n7190 & n11850 ) | ( n10283 & n11850 ) ;
  assign n11852 = n11850 | n11851 ;
  assign n11853 = ( n7192 & n10282 ) | ( n7192 & n11850 ) | ( n10282 & n11850 ) ;
  assign n11854 = n11852 | n11853 ;
  assign n11855 = n7196 & n11098 ;
  assign n11856 = n11854 | n11855 ;
  assign n11857 = n11856 ^ x23 ^ 1'b0 ;
  assign n11858 = ( n11749 & n11798 ) | ( n11749 & n11857 ) | ( n11798 & n11857 ) ;
  assign n11859 = n11857 ^ n11798 ^ n11749 ;
  assign n11860 = n7339 & n10306 ;
  assign n11861 = ( n7337 & ~n10340 ) | ( n7337 & n11860 ) | ( ~n10340 & n11860 ) ;
  assign n11862 = n11860 | n11861 ;
  assign n11863 = ( n7338 & ~n10280 ) | ( n7338 & n11860 ) | ( ~n10280 & n11860 ) ;
  assign n11864 = n11862 | n11863 ;
  assign n11865 = n7340 & ~n11264 ;
  assign n11866 = n11864 & ~n11865 ;
  assign n11867 = n11866 ^ n11865 ^ x20 ;
  assign n11868 = ( n11849 & n11859 ) | ( n11849 & n11867 ) | ( n11859 & n11867 ) ;
  assign n11869 = n11867 ^ n11859 ^ n11849 ;
  assign n11870 = n7485 & n10282 ;
  assign n11871 = ( n7486 & n10278 ) | ( n7486 & n11870 ) | ( n10278 & n11870 ) ;
  assign n11872 = n11870 | n11871 ;
  assign n11873 = ( n7493 & n10283 ) | ( n7493 & n11870 ) | ( n10283 & n11870 ) ;
  assign n11874 = n11872 | n11873 ;
  assign n11875 = n7487 & n11098 ;
  assign n11876 = n11874 | n11875 ;
  assign n11877 = n11876 ^ x17 ^ 1'b0 ;
  assign n11878 = n7669 & n10282 ;
  assign n11879 = ( n11641 & n11653 ) | ( n11641 & n11877 ) | ( n11653 & n11877 ) ;
  assign n11880 = n11877 ^ n11653 ^ n11641 ;
  assign n11881 = n7829 & n10282 ;
  assign n11882 = ( n7833 & n10283 ) | ( n7833 & n11881 ) | ( n10283 & n11881 ) ;
  assign n11883 = n11881 | n11882 ;
  assign n11884 = ( n7834 & n10278 ) | ( n7834 & n11881 ) | ( n10278 & n11881 ) ;
  assign n11885 = n11883 | n11884 ;
  assign n11886 = ( n7674 & n10283 ) | ( n7674 & n11878 ) | ( n10283 & n11878 ) ;
  assign n11887 = n11878 | n11886 ;
  assign n11888 = ( n7667 & n10278 ) | ( n7667 & n11878 ) | ( n10278 & n11878 ) ;
  assign n11889 = n11887 | n11888 ;
  assign n11890 = n7666 & n11098 ;
  assign n11891 = n11889 | n11890 ;
  assign n11892 = n7838 & n11098 ;
  assign n11893 = n11891 ^ x14 ^ 1'b0 ;
  assign n11894 = n11885 | n11892 ;
  assign n11895 = ( n11550 & n11567 ) | ( n11550 & n11893 ) | ( n11567 & n11893 ) ;
  assign n11896 = n11893 ^ n11567 ^ n11550 ;
  assign n11897 = n7669 & n10278 ;
  assign n11898 = ( n7674 & n10282 ) | ( n7674 & n11897 ) | ( n10282 & n11897 ) ;
  assign n11899 = n11897 | n11898 ;
  assign n11900 = ( n7667 & ~n10280 ) | ( n7667 & n11897 ) | ( ~n10280 & n11897 ) ;
  assign n11901 = n11899 | n11900 ;
  assign n11902 = n7666 & ~n11158 ;
  assign n11903 = n11901 & ~n11902 ;
  assign n11904 = n11894 ^ x11 ^ 1'b0 ;
  assign n11905 = n11903 ^ n11902 ^ x14 ;
  assign n11906 = n11905 ^ n11895 ^ n11603 ;
  assign n11907 = ( n11603 & n11895 ) | ( n11603 & n11905 ) | ( n11895 & n11905 ) ;
  assign n11908 = n7037 & n10278 ;
  assign n11909 = ( n7036 & n10282 ) | ( n7036 & n11908 ) | ( n10282 & n11908 ) ;
  assign n11910 = n11908 | n11909 ;
  assign n11911 = ( n7052 & n10283 ) | ( n7052 & n11908 ) | ( n10283 & n11908 ) ;
  assign n11912 = n11910 | n11911 ;
  assign n11913 = ( n7035 & n11098 ) | ( n7035 & n11912 ) | ( n11098 & n11912 ) ;
  assign n11914 = n11912 | n11913 ;
  assign n11915 = n11914 ^ x26 ^ 1'b0 ;
  assign n11916 = n11915 ^ n11809 ^ n11728 ;
  assign n11917 = ( ~n11728 & n11809 ) | ( ~n11728 & n11915 ) | ( n11809 & n11915 ) ;
  assign n11918 = n11904 ^ n11529 ^ n11469 ;
  assign n11919 = n7485 & n10278 ;
  assign n11920 = n6918 & n11098 ;
  assign n11921 = ( n11469 & n11529 ) | ( n11469 & n11904 ) | ( n11529 & n11904 ) ;
  assign n11922 = n6901 & n10282 ;
  assign n11923 = ( n6906 & n10283 ) | ( n6906 & n11922 ) | ( n10283 & n11922 ) ;
  assign n11924 = ( n7486 & ~n10280 ) | ( n7486 & n11919 ) | ( ~n10280 & n11919 ) ;
  assign n11925 = n11922 | n11923 ;
  assign n11926 = n11919 | n11924 ;
  assign n11927 = ( n7493 & n10282 ) | ( n7493 & n11919 ) | ( n10282 & n11919 ) ;
  assign n11928 = ( n6907 & n10278 ) | ( n6907 & n11922 ) | ( n10278 & n11922 ) ;
  assign n11929 = n11925 | n11928 ;
  assign n11930 = n11920 | n11929 ;
  assign n11931 = n11926 | n11927 ;
  assign n11932 = n11930 ^ x29 ^ 1'b0 ;
  assign n11933 = n7829 & n10278 ;
  assign n11934 = ( n7833 & n10282 ) | ( n7833 & n11933 ) | ( n10282 & n11933 ) ;
  assign n11935 = n11933 | n11934 ;
  assign n11936 = ( n7834 & ~n10280 ) | ( n7834 & n11933 ) | ( ~n10280 & n11933 ) ;
  assign n11937 = n11935 | n11936 ;
  assign n11938 = n7838 & ~n11158 ;
  assign n11939 = n11932 ^ n11818 ^ n11059 ;
  assign n11940 = n11937 & ~n11938 ;
  assign n11941 = ( ~n11059 & n11818 ) | ( ~n11059 & n11932 ) | ( n11818 & n11932 ) ;
  assign n11942 = n7487 & ~n11158 ;
  assign n11943 = n11931 & ~n11942 ;
  assign n11944 = n11940 ^ n11938 ^ x11 ;
  assign n11945 = ( n11542 & n11921 ) | ( n11542 & n11944 ) | ( n11921 & n11944 ) ;
  assign n11946 = n11943 ^ n11942 ^ x17 ;
  assign n11947 = ( n11662 & n11879 ) | ( n11662 & n11946 ) | ( n11879 & n11946 ) ;
  assign n11948 = n11944 ^ n11921 ^ n11542 ;
  assign n11949 = n11946 ^ n11879 ^ n11662 ;
  assign n11950 = n6901 & n10278 ;
  assign n11951 = ( n6906 & n10282 ) | ( n6906 & n11950 ) | ( n10282 & n11950 ) ;
  assign n11952 = n11950 | n11951 ;
  assign n11953 = ( n6907 & ~n10280 ) | ( n6907 & n11950 ) | ( ~n10280 & n11950 ) ;
  assign n11954 = n11952 | n11953 ;
  assign n11955 = n6918 & ~n11158 ;
  assign n11956 = n11954 | n11955 ;
  assign n11957 = n11956 ^ x29 ^ 1'b0 ;
  assign n11958 = ( ~n11075 & n11941 ) | ( ~n11075 & n11957 ) | ( n11941 & n11957 ) ;
  assign n11959 = n11957 ^ n11941 ^ n11075 ;
  assign n11960 = n6901 & ~n10280 ;
  assign n11961 = ( n6906 & n10278 ) | ( n6906 & n11960 ) | ( n10278 & n11960 ) ;
  assign n11962 = n11960 | n11961 ;
  assign n11963 = ( n6907 & n10306 ) | ( n6907 & n11960 ) | ( n10306 & n11960 ) ;
  assign n11964 = n11962 | n11963 ;
  assign n11965 = n6918 & ~n11223 ;
  assign n11966 = n11964 & ~n11965 ;
  assign n11967 = n11966 ^ n11965 ^ x29 ;
  assign n11968 = ( n11097 & n11958 ) | ( n11097 & n11967 ) | ( n11958 & n11967 ) ;
  assign n11969 = n11967 ^ n11958 ^ n11097 ;
  assign n11970 = n7037 & ~n10280 ;
  assign n11971 = ( n7036 & n10278 ) | ( n7036 & n11970 ) | ( n10278 & n11970 ) ;
  assign n11972 = n11970 | n11971 ;
  assign n11973 = ( n7052 & n10282 ) | ( n7052 & n11970 ) | ( n10282 & n11970 ) ;
  assign n11974 = n11972 | n11973 ;
  assign n11975 = n7188 & ~n10280 ;
  assign n11976 = ( n7190 & n10282 ) | ( n7190 & n11975 ) | ( n10282 & n11975 ) ;
  assign n11977 = n11975 | n11976 ;
  assign n11978 = ( n7192 & n10278 ) | ( n7192 & n11975 ) | ( n10278 & n11975 ) ;
  assign n11979 = n11977 | n11978 ;
  assign n11980 = n7196 & ~n11158 ;
  assign n11981 = n11979 & ~n11980 ;
  assign n11982 = n11981 ^ n11980 ^ x23 ;
  assign n11983 = n11982 ^ n11858 ^ n11776 ;
  assign n11984 = n7035 & ~n11158 ;
  assign n11985 = ( n11776 & n11858 ) | ( n11776 & n11982 ) | ( n11858 & n11982 ) ;
  assign n11986 = n11974 & ~n11984 ;
  assign n11987 = n7829 & ~n10280 ;
  assign n11988 = n11986 ^ n11984 ^ x26 ;
  assign n11989 = ( ~n11739 & n11917 ) | ( ~n11739 & n11988 ) | ( n11917 & n11988 ) ;
  assign n11990 = n11988 ^ n11917 ^ n11739 ;
  assign n11991 = ( n7833 & n10278 ) | ( n7833 & n11987 ) | ( n10278 & n11987 ) ;
  assign n11992 = n11987 | n11991 ;
  assign n11993 = ( n7834 & n10306 ) | ( n7834 & n11987 ) | ( n10306 & n11987 ) ;
  assign n11994 = n11992 | n11993 ;
  assign n11995 = n7838 & ~n11223 ;
  assign n11996 = n11994 & ~n11995 ;
  assign n11997 = n11996 ^ n11995 ^ x11 ;
  assign n11998 = ( n11547 & n11945 ) | ( n11547 & n11997 ) | ( n11945 & n11997 ) ;
  assign n11999 = n11997 ^ n11945 ^ n11547 ;
  assign n12000 = n7669 & ~n10280 ;
  assign n12001 = ( n7674 & n10278 ) | ( n7674 & n12000 ) | ( n10278 & n12000 ) ;
  assign n12002 = n12000 | n12001 ;
  assign n12003 = ( n7667 & n10306 ) | ( n7667 & n12000 ) | ( n10306 & n12000 ) ;
  assign n12004 = n12002 | n12003 ;
  assign n12005 = n7666 & ~n11223 ;
  assign n12006 = n12004 & ~n12005 ;
  assign n12007 = n12006 ^ n12005 ^ x14 ;
  assign n12008 = n12007 ^ n11907 ^ n11652 ;
  assign n12009 = ( n11652 & n11907 ) | ( n11652 & n12007 ) | ( n11907 & n12007 ) ;
  assign n12010 = n7188 & n10306 ;
  assign n12011 = ( n7190 & n10278 ) | ( n7190 & n12010 ) | ( n10278 & n12010 ) ;
  assign n12012 = n12010 | n12011 ;
  assign n12013 = ( n7192 & ~n10280 ) | ( n7192 & n12010 ) | ( ~n10280 & n12010 ) ;
  assign n12014 = n12012 | n12013 ;
  assign n12015 = n7196 & ~n11223 ;
  assign n12016 = n12014 & ~n12015 ;
  assign n12017 = n12016 ^ n12015 ^ x23 ;
  assign n12018 = ( n11808 & n11985 ) | ( n11808 & n12017 ) | ( n11985 & n12017 ) ;
  assign n12019 = n12017 ^ n11985 ^ n11808 ;
  assign n12020 = n7037 & n10306 ;
  assign n12021 = ( n7036 & ~n10280 ) | ( n7036 & n12020 ) | ( ~n10280 & n12020 ) ;
  assign n12022 = n12020 | n12021 ;
  assign n12023 = ( n7052 & n10278 ) | ( n7052 & n12020 ) | ( n10278 & n12020 ) ;
  assign n12024 = n12022 | n12023 ;
  assign n12025 = n7487 & ~n11223 ;
  assign n12026 = n7035 & ~n11223 ;
  assign n12027 = n12024 & ~n12026 ;
  assign n12028 = n12027 ^ n12026 ^ x26 ;
  assign n12029 = ( n11819 & n11989 ) | ( n11819 & n12028 ) | ( n11989 & n12028 ) ;
  assign n12030 = n12028 ^ n11989 ^ n11819 ;
  assign n12031 = n7485 & ~n10280 ;
  assign n12032 = ( n7486 & n10306 ) | ( n7486 & n12031 ) | ( n10306 & n12031 ) ;
  assign n12033 = ( n7493 & n10278 ) | ( n7493 & n12031 ) | ( n10278 & n12031 ) ;
  assign n12034 = n12031 | n12032 ;
  assign n12035 = n12033 | n12034 ;
  assign n12036 = ~n12025 & n12035 ;
  assign n12037 = n12036 ^ n12025 ^ x17 ;
  assign n12038 = n12037 ^ n11947 ^ n11788 ;
  assign n12039 = ( n11788 & n11947 ) | ( n11788 & n12037 ) | ( n11947 & n12037 ) ;
  assign n12040 = n7485 & n10306 ;
  assign n12041 = n7932 & n10306 ;
  assign n12042 = ( n7943 & ~n10280 ) | ( n7943 & n12041 ) | ( ~n10280 & n12041 ) ;
  assign n12043 = n12041 | n12042 ;
  assign n12044 = ( n7929 & ~n10340 ) | ( n7929 & n12041 ) | ( ~n10340 & n12041 ) ;
  assign n12045 = n7930 & ~n11264 ;
  assign n12046 = n12043 | n12044 ;
  assign n12047 = ~n12045 & n12046 ;
  assign n12048 = n12047 ^ n12045 ^ x8 ;
  assign n12049 = n12048 ^ n11918 ^ n11479 ;
  assign n12050 = n7829 & n10306 ;
  assign n12051 = ( n11479 & n11918 ) | ( n11479 & n12048 ) | ( n11918 & n12048 ) ;
  assign n12052 = ( n7834 & ~n10340 ) | ( n7834 & n12050 ) | ( ~n10340 & n12050 ) ;
  assign n12053 = ( n7833 & ~n10280 ) | ( n7833 & n12050 ) | ( ~n10280 & n12050 ) ;
  assign n12054 = n12050 | n12053 ;
  assign n12055 = n12052 | n12054 ;
  assign n12056 = ( n7486 & ~n10340 ) | ( n7486 & n12040 ) | ( ~n10340 & n12040 ) ;
  assign n12057 = ( n7493 & ~n10280 ) | ( n7493 & n12040 ) | ( ~n10280 & n12040 ) ;
  assign n12058 = n12040 | n12056 ;
  assign n12059 = n12057 | n12058 ;
  assign n12060 = n7669 & n10306 ;
  assign n12061 = ( n7674 & ~n10280 ) | ( n7674 & n12060 ) | ( ~n10280 & n12060 ) ;
  assign n12062 = n12060 | n12061 ;
  assign n12063 = ( n7667 & ~n10340 ) | ( n7667 & n12060 ) | ( ~n10340 & n12060 ) ;
  assign n12064 = n12062 | n12063 ;
  assign n12065 = n7487 & ~n11264 ;
  assign n12066 = n12059 & ~n12065 ;
  assign n12067 = n12066 ^ n12065 ^ x17 ;
  assign n12068 = ( n11829 & n12039 ) | ( n11829 & n12067 ) | ( n12039 & n12067 ) ;
  assign n12069 = n12067 ^ n12039 ^ n11829 ;
  assign n12070 = n7838 & ~n11264 ;
  assign n12071 = n12055 & ~n12070 ;
  assign n12072 = n6901 & ~n10340 ;
  assign n12073 = n12071 ^ n12070 ^ x11 ;
  assign n12074 = n7666 & ~n11264 ;
  assign n12075 = n12064 & ~n12074 ;
  assign n12076 = n12075 ^ n12074 ^ x14 ;
  assign n12077 = n12076 ^ n12009 ^ n11880 ;
  assign n12078 = ( n11880 & n12009 ) | ( n11880 & n12076 ) | ( n12009 & n12076 ) ;
  assign n12079 = ( n6906 & n10306 ) | ( n6906 & n12072 ) | ( n10306 & n12072 ) ;
  assign n12080 = ( n6907 & n10353 ) | ( n6907 & n12072 ) | ( n10353 & n12072 ) ;
  assign n12081 = n12072 | n12079 ;
  assign n12082 = n7188 & ~n10340 ;
  assign n12083 = n12080 | n12081 ;
  assign n12084 = n6918 & ~n11314 ;
  assign n12085 = n12083 & ~n12084 ;
  assign n12086 = n12085 ^ n12084 ^ x29 ;
  assign n12087 = ( n7190 & ~n10280 ) | ( n7190 & n12082 ) | ( ~n10280 & n12082 ) ;
  assign n12088 = n12082 | n12087 ;
  assign n12089 = ( n7192 & n10306 ) | ( n7192 & n12082 ) | ( n10306 & n12082 ) ;
  assign n12090 = n12088 | n12089 ;
  assign n12091 = n12073 ^ n11998 ^ n11896 ;
  assign n12092 = ( n11896 & n11998 ) | ( n11896 & n12073 ) | ( n11998 & n12073 ) ;
  assign n12093 = n7037 & ~n10340 ;
  assign n12094 = n7196 & ~n11264 ;
  assign n12095 = n12090 | n12094 ;
  assign n12096 = ( n7036 & n10306 ) | ( n7036 & n12093 ) | ( n10306 & n12093 ) ;
  assign n12097 = n12093 | n12096 ;
  assign n12098 = ( n7052 & ~n10280 ) | ( n7052 & n12093 ) | ( ~n10280 & n12093 ) ;
  assign n12099 = n12097 | n12098 ;
  assign n12100 = n6918 & ~n11264 ;
  assign n12101 = n7035 & ~n11264 ;
  assign n12102 = n12099 & ~n12101 ;
  assign n12103 = n12102 ^ n12101 ^ x26 ;
  assign n12104 = n12103 ^ n12029 ^ n11939 ;
  assign n12105 = ( ~n11939 & n12029 ) | ( ~n11939 & n12103 ) | ( n12029 & n12103 ) ;
  assign n12106 = n12095 ^ x23 ^ 1'b0 ;
  assign n12107 = ( ~n11916 & n12018 ) | ( ~n11916 & n12106 ) | ( n12018 & n12106 ) ;
  assign n12108 = n6901 & n10306 ;
  assign n12109 = ( n6906 & ~n10280 ) | ( n6906 & n12108 ) | ( ~n10280 & n12108 ) ;
  assign n12110 = n12108 | n12109 ;
  assign n12111 = ( n6907 & ~n10340 ) | ( n6907 & n12108 ) | ( ~n10340 & n12108 ) ;
  assign n12112 = n12110 | n12111 ;
  assign n12113 = ~n12100 & n12112 ;
  assign n12114 = n12113 ^ n12100 ^ x29 ;
  assign n12115 = n12114 ^ n11968 ^ n11108 ;
  assign n12116 = ( n11108 & n11968 ) | ( n11108 & n12114 ) | ( n11968 & n12114 ) ;
  assign n12117 = n12106 ^ n12018 ^ n11916 ;
  assign n12118 = ( n11167 & n12086 ) | ( n11167 & n12116 ) | ( n12086 & n12116 ) ;
  assign n12119 = n12116 ^ n12086 ^ n11167 ;
  assign n12120 = n7932 & ~n10340 ;
  assign n12121 = ( n7943 & n10306 ) | ( n7943 & n12120 ) | ( n10306 & n12120 ) ;
  assign n12122 = ( n7929 & n10353 ) | ( n7929 & n12120 ) | ( n10353 & n12120 ) ;
  assign n12123 = n12120 | n12121 ;
  assign n12124 = n7485 & ~n10340 ;
  assign n12125 = ( n7486 & n10353 ) | ( n7486 & n12124 ) | ( n10353 & n12124 ) ;
  assign n12126 = n12122 | n12123 ;
  assign n12127 = n7487 & ~n11314 ;
  assign n12128 = n12124 | n12125 ;
  assign n12129 = ( n7493 & n10306 ) | ( n7493 & n12124 ) | ( n10306 & n12124 ) ;
  assign n12130 = n12128 | n12129 ;
  assign n12131 = n12127 | n12130 ;
  assign n12132 = n7037 & n10353 ;
  assign n12133 = ( n7036 & ~n10340 ) | ( n7036 & n12132 ) | ( ~n10340 & n12132 ) ;
  assign n12134 = n12131 ^ x17 ^ 1'b0 ;
  assign n12135 = n12132 | n12133 ;
  assign n12136 = ( n7052 & n10306 ) | ( n7052 & n12132 ) | ( n10306 & n12132 ) ;
  assign n12137 = n12135 | n12136 ;
  assign n12138 = n12134 ^ n12068 ^ n11838 ;
  assign n12139 = ( n11838 & n12068 ) | ( n11838 & n12134 ) | ( n12068 & n12134 ) ;
  assign n12140 = n7035 & ~n11314 ;
  assign n12141 = n12137 & ~n12140 ;
  assign n12142 = n12141 ^ n12140 ^ x26 ;
  assign n12143 = n7188 & n10353 ;
  assign n12144 = ( n7190 & n10306 ) | ( n7190 & n12143 ) | ( n10306 & n12143 ) ;
  assign n12145 = n12143 | n12144 ;
  assign n12146 = ( n7192 & ~n10340 ) | ( n7192 & n12143 ) | ( ~n10340 & n12143 ) ;
  assign n12147 = n12145 | n12146 ;
  assign n12148 = n12142 ^ n12105 ^ n11959 ;
  assign n12149 = ( ~n11959 & n12105 ) | ( ~n11959 & n12142 ) | ( n12105 & n12142 ) ;
  assign n12150 = n7196 & ~n11314 ;
  assign n12151 = n12147 | n12150 ;
  assign n12152 = n7669 & ~n10340 ;
  assign n12153 = n12151 ^ x23 ^ 1'b0 ;
  assign n12154 = ( n7674 & n10306 ) | ( n7674 & n12152 ) | ( n10306 & n12152 ) ;
  assign n12155 = n12152 | n12154 ;
  assign n12156 = ( n7667 & n10353 ) | ( n7667 & n12152 ) | ( n10353 & n12152 ) ;
  assign n12157 = n12155 | n12156 ;
  assign n12158 = ( ~n11990 & n12107 ) | ( ~n11990 & n12153 ) | ( n12107 & n12153 ) ;
  assign n12159 = n12153 ^ n12107 ^ n11990 ;
  assign n12160 = n7930 & ~n11314 ;
  assign n12161 = n6791 & ~n10340 ;
  assign n12162 = n12126 | n12160 ;
  assign n12163 = ( n6788 & n10353 ) | ( n6788 & n12161 ) | ( n10353 & n12161 ) ;
  assign n12164 = n12161 | n12163 ;
  assign n12165 = ( n6790 & n10306 ) | ( n6790 & n12161 ) | ( n10306 & n12161 ) ;
  assign n12166 = n12164 | n12165 ;
  assign n12167 = n6789 & ~n11314 ;
  assign n12168 = n12166 | n12167 ;
  assign n12169 = n7666 & ~n11314 ;
  assign n12170 = n12157 | n12169 ;
  assign n12171 = n12162 ^ x8 ^ 1'b0 ;
  assign n12172 = ( n11948 & n12051 ) | ( n11948 & n12171 ) | ( n12051 & n12171 ) ;
  assign n12173 = n12171 ^ n12051 ^ n11948 ;
  assign n12174 = n7339 & ~n10340 ;
  assign n12175 = ( n7337 & n10353 ) | ( n7337 & n12174 ) | ( n10353 & n12174 ) ;
  assign n12176 = n12174 | n12175 ;
  assign n12177 = ( n7338 & n10306 ) | ( n7338 & n12174 ) | ( n10306 & n12174 ) ;
  assign n12178 = n12176 | n12177 ;
  assign n12179 = n7340 & ~n11314 ;
  assign n12180 = n12178 | n12179 ;
  assign n12181 = n7829 & ~n10340 ;
  assign n12182 = n7838 & ~n11314 ;
  assign n12183 = ( n7833 & n10306 ) | ( n7833 & n12181 ) | ( n10306 & n12181 ) ;
  assign n12184 = n12180 ^ x20 ^ 1'b0 ;
  assign n12185 = n12181 | n12183 ;
  assign n12186 = ( n7834 & n10353 ) | ( n7834 & n12181 ) | ( n10353 & n12181 ) ;
  assign n12187 = n12185 | n12186 ;
  assign n12188 = n12182 | n12187 ;
  assign n12189 = n12188 ^ x11 ^ 1'b0 ;
  assign n12190 = n12189 ^ n12092 ^ n11906 ;
  assign n12191 = n12170 ^ x14 ^ 1'b0 ;
  assign n12192 = ( n11949 & n12078 ) | ( n11949 & n12191 ) | ( n12078 & n12191 ) ;
  assign n12193 = ( n11906 & n12092 ) | ( n11906 & n12189 ) | ( n12092 & n12189 ) ;
  assign n12194 = n12191 ^ n12078 ^ n11949 ;
  assign n12195 = ( n11868 & n11983 ) | ( n11868 & n12184 ) | ( n11983 & n12184 ) ;
  assign n12196 = n12184 ^ n11983 ^ n11868 ;
  assign n12197 = n7339 & n10353 ;
  assign n12198 = ( n7337 & n10372 ) | ( n7337 & n12197 ) | ( n10372 & n12197 ) ;
  assign n12199 = n12197 | n12198 ;
  assign n12200 = ( n7338 & ~n10340 ) | ( n7338 & n12197 ) | ( ~n10340 & n12197 ) ;
  assign n12201 = n12199 | n12200 ;
  assign n12202 = n7340 & n11365 ;
  assign n12203 = n12201 | n12202 ;
  assign n12204 = n12203 ^ x20 ^ 1'b0 ;
  assign n12205 = ( n12019 & n12195 ) | ( n12019 & n12204 ) | ( n12195 & n12204 ) ;
  assign n12206 = n12204 ^ n12195 ^ n12019 ;
  assign n12207 = n7485 & n10353 ;
  assign n12208 = ( n7486 & n10372 ) | ( n7486 & n12207 ) | ( n10372 & n12207 ) ;
  assign n12209 = n12207 | n12208 ;
  assign n12210 = ( n7493 & ~n10340 ) | ( n7493 & n12207 ) | ( ~n10340 & n12207 ) ;
  assign n12211 = n12209 | n12210 ;
  assign n12212 = n7487 & n11365 ;
  assign n12213 = n12211 | n12212 ;
  assign n12214 = n12213 ^ x17 ^ 1'b0 ;
  assign n12215 = ( n11848 & n12139 ) | ( n11848 & n12214 ) | ( n12139 & n12214 ) ;
  assign n12216 = n12214 ^ n12139 ^ n11848 ;
  assign n12217 = n7188 & n10372 ;
  assign n12218 = ( n7190 & ~n10340 ) | ( n7190 & n12217 ) | ( ~n10340 & n12217 ) ;
  assign n12219 = n12217 | n12218 ;
  assign n12220 = ( n7192 & n10353 ) | ( n7192 & n12217 ) | ( n10353 & n12217 ) ;
  assign n12221 = n12219 | n12220 ;
  assign n12222 = n7196 & n11365 ;
  assign n12223 = n12221 | n12222 ;
  assign n12224 = n12223 ^ x23 ^ 1'b0 ;
  assign n12225 = ( n12030 & n12158 ) | ( n12030 & n12224 ) | ( n12158 & n12224 ) ;
  assign n12226 = n12224 ^ n12158 ^ n12030 ;
  assign n12227 = n7669 & n10353 ;
  assign n12228 = ( n7674 & ~n10340 ) | ( n7674 & n12227 ) | ( ~n10340 & n12227 ) ;
  assign n12229 = n12227 | n12228 ;
  assign n12230 = ( n7667 & n10372 ) | ( n7667 & n12227 ) | ( n10372 & n12227 ) ;
  assign n12231 = n12229 | n12230 ;
  assign n12232 = n7666 & n11365 ;
  assign n12233 = n12231 | n12232 ;
  assign n12234 = n12233 ^ x14 ^ 1'b0 ;
  assign n12235 = ( n12038 & n12192 ) | ( n12038 & n12234 ) | ( n12192 & n12234 ) ;
  assign n12236 = n12234 ^ n12192 ^ n12038 ;
  assign n12237 = n7829 & n10353 ;
  assign n12238 = ( n7833 & ~n10340 ) | ( n7833 & n12237 ) | ( ~n10340 & n12237 ) ;
  assign n12239 = n12237 | n12238 ;
  assign n12240 = ( n7834 & n10372 ) | ( n7834 & n12237 ) | ( n10372 & n12237 ) ;
  assign n12241 = n12239 | n12240 ;
  assign n12242 = n7838 & n11365 ;
  assign n12243 = n12241 | n12242 ;
  assign n12244 = n12243 ^ x11 ^ 1'b0 ;
  assign n12245 = ( n12008 & n12193 ) | ( n12008 & n12244 ) | ( n12193 & n12244 ) ;
  assign n12246 = n12244 ^ n12193 ^ n12008 ;
  assign n12247 = n7037 & n10372 ;
  assign n12248 = ( n7036 & n10353 ) | ( n7036 & n12247 ) | ( n10353 & n12247 ) ;
  assign n12249 = n12247 | n12248 ;
  assign n12250 = ( n7052 & ~n10340 ) | ( n7052 & n12247 ) | ( ~n10340 & n12247 ) ;
  assign n12251 = n12249 | n12250 ;
  assign n12252 = ( n7035 & n11365 ) | ( n7035 & n12251 ) | ( n11365 & n12251 ) ;
  assign n12253 = n12251 | n12252 ;
  assign n12254 = n12253 ^ x26 ^ 1'b0 ;
  assign n12255 = n12254 ^ n12149 ^ n11969 ;
  assign n12256 = ( n11969 & n12149 ) | ( n11969 & n12254 ) | ( n12149 & n12254 ) ;
  assign n12257 = ( ~x2 & n8085 ) | ( ~x2 & n8090 ) | ( n8085 & n8090 ) ;
  assign n12258 = n7932 & n10353 ;
  assign n12259 = ( n7943 & ~n10340 ) | ( n7943 & n12258 ) | ( ~n10340 & n12258 ) ;
  assign n12260 = n12258 | n12259 ;
  assign n12261 = ( n7929 & n10372 ) | ( n7929 & n12258 ) | ( n10372 & n12258 ) ;
  assign n12262 = n12260 | n12261 ;
  assign n12263 = n7930 & n11365 ;
  assign n12264 = n12262 | n12263 ;
  assign n12265 = n12264 ^ x8 ^ 1'b0 ;
  assign n12266 = ( n11999 & n12172 ) | ( n11999 & n12265 ) | ( n12172 & n12265 ) ;
  assign n12267 = n12265 ^ n12172 ^ n11999 ;
  assign n12268 = ( ~n6633 & n12168 ) | ( ~n6633 & n12257 ) | ( n12168 & n12257 ) ;
  assign n12269 = n6791 & n10353 ;
  assign n12270 = n12257 ^ n12168 ^ n6633 ;
  assign n12271 = ( n6788 & n10372 ) | ( n6788 & n12269 ) | ( n10372 & n12269 ) ;
  assign n12272 = n12269 | n12271 ;
  assign n12273 = ( n6790 & ~n10340 ) | ( n6790 & n12269 ) | ( ~n10340 & n12269 ) ;
  assign n12274 = n12272 | n12273 ;
  assign n12275 = n6901 & n10353 ;
  assign n12276 = ( n6906 & ~n10340 ) | ( n6906 & n12275 ) | ( ~n10340 & n12275 ) ;
  assign n12277 = n12275 | n12276 ;
  assign n12278 = ( n6907 & n10372 ) | ( n6907 & n12275 ) | ( n10372 & n12275 ) ;
  assign n12279 = n12277 | n12278 ;
  assign n12280 = ( n6918 & n11365 ) | ( n6918 & n12279 ) | ( n11365 & n12279 ) ;
  assign n12281 = n12279 | n12280 ;
  assign n12282 = n6789 & ~n11365 ;
  assign n12283 = ( n6789 & n12274 ) | ( n6789 & ~n12282 ) | ( n12274 & ~n12282 ) ;
  assign n12284 = n12281 ^ x29 ^ 1'b0 ;
  assign n12285 = n12284 ^ n12118 ^ n11283 ;
  assign n12286 = ( n10353 & n10372 ) | ( n10353 & n11315 ) | ( n10372 & n11315 ) ;
  assign n12287 = ( n11283 & n12118 ) | ( n11283 & n12284 ) | ( n12118 & n12284 ) ;
  assign n12288 = n8086 & n10353 ;
  assign n12289 = ( n6710 & n12257 ) | ( n6710 & n12268 ) | ( n12257 & n12268 ) ;
  assign n12290 = ( n8088 & n10372 ) | ( n8088 & n12288 ) | ( n10372 & n12288 ) ;
  assign n12291 = n12268 ^ n12257 ^ n6710 ;
  assign n12292 = ( n8090 & n10408 ) | ( n8090 & n12288 ) | ( n10408 & n12288 ) ;
  assign n12293 = n12288 | n12290 ;
  assign n12294 = n12292 | n12293 ;
  assign n12295 = n12286 ^ n10408 ^ n10372 ;
  assign n12296 = n8089 & n12295 ;
  assign n12297 = n12294 | n12296 ;
  assign n12298 = n12297 ^ x2 ^ 1'b0 ;
  assign n12299 = ( n11369 & n11408 ) | ( n11369 & n12298 ) | ( n11408 & n12298 ) ;
  assign n12300 = n7669 & n10372 ;
  assign n12301 = ( n7674 & n10353 ) | ( n7674 & n12300 ) | ( n10353 & n12300 ) ;
  assign n12302 = n12300 | n12301 ;
  assign n12303 = n7932 & n10372 ;
  assign n12304 = ( n7667 & n10408 ) | ( n7667 & n12300 ) | ( n10408 & n12300 ) ;
  assign n12305 = n12302 | n12304 ;
  assign n12306 = ( n7943 & n10353 ) | ( n7943 & n12303 ) | ( n10353 & n12303 ) ;
  assign n12307 = n12303 | n12306 ;
  assign n12308 = ( n7929 & n10408 ) | ( n7929 & n12303 ) | ( n10408 & n12303 ) ;
  assign n12309 = n12307 | n12308 ;
  assign n12310 = n7930 & n12295 ;
  assign n12311 = n12309 | n12310 ;
  assign n12312 = n7666 & n12295 ;
  assign n12313 = n12305 | n12312 ;
  assign n12314 = n12313 ^ x14 ^ 1'b0 ;
  assign n12315 = ( n12069 & n12235 ) | ( n12069 & n12314 ) | ( n12235 & n12314 ) ;
  assign n12316 = n12314 ^ n12235 ^ n12069 ;
  assign n12317 = n8086 & n10372 ;
  assign n12318 = ( n8088 & n10408 ) | ( n8088 & n12317 ) | ( n10408 & n12317 ) ;
  assign n12319 = n12317 | n12318 ;
  assign n12320 = ( n8090 & n10419 ) | ( n8090 & n12317 ) | ( n10419 & n12317 ) ;
  assign n12321 = ( n10372 & n10408 ) | ( n10372 & n12286 ) | ( n10408 & n12286 ) ;
  assign n12322 = n12319 | n12320 ;
  assign n12323 = n12311 ^ x8 ^ 1'b0 ;
  assign n12324 = ( n12091 & n12266 ) | ( n12091 & n12323 ) | ( n12266 & n12323 ) ;
  assign n12325 = n12323 ^ n12266 ^ n12091 ;
  assign n12326 = n12321 ^ n10419 ^ n10408 ;
  assign n12327 = ( n8089 & n12322 ) | ( n8089 & n12326 ) | ( n12322 & n12326 ) ;
  assign n12328 = n12322 | n12327 ;
  assign n12329 = n12328 ^ x2 ^ 1'b0 ;
  assign n12330 = ( n11448 & n12299 ) | ( n11448 & n12329 ) | ( n12299 & n12329 ) ;
  assign n12331 = n6901 & n10408 ;
  assign n12332 = ( n6906 & n10372 ) | ( n6906 & n12331 ) | ( n10372 & n12331 ) ;
  assign n12333 = n12331 | n12332 ;
  assign n12334 = ( n6907 & n10419 ) | ( n6907 & n12331 ) | ( n10419 & n12331 ) ;
  assign n12335 = n12333 | n12334 ;
  assign n12336 = n7669 & n10408 ;
  assign n12337 = ( n7674 & n10372 ) | ( n7674 & n12336 ) | ( n10372 & n12336 ) ;
  assign n12338 = n12336 | n12337 ;
  assign n12339 = ( n7667 & n10419 ) | ( n7667 & n12336 ) | ( n10419 & n12336 ) ;
  assign n12340 = n12338 | n12339 ;
  assign n12341 = ( n7666 & n12326 ) | ( n7666 & n12340 ) | ( n12326 & n12340 ) ;
  assign n12342 = n12340 | n12341 ;
  assign n12343 = n12342 ^ x14 ^ 1'b0 ;
  assign n12344 = ( n12138 & n12315 ) | ( n12138 & n12343 ) | ( n12315 & n12343 ) ;
  assign n12345 = n12343 ^ n12315 ^ n12138 ;
  assign n12346 = ( n6918 & n12326 ) | ( n6918 & n12335 ) | ( n12326 & n12335 ) ;
  assign n12347 = n12335 | n12346 ;
  assign n12348 = n12347 ^ x29 ^ 1'b0 ;
  assign n12349 = n12348 ^ n12270 ^ n11328 ;
  assign n12350 = ( n11328 & ~n12270 ) | ( n11328 & n12348 ) | ( ~n12270 & n12348 ) ;
  assign n12351 = ( n12283 & n12291 ) | ( n12283 & n12350 ) | ( n12291 & n12350 ) ;
  assign n12352 = n7932 & n10408 ;
  assign n12353 = ( n7943 & n10372 ) | ( n7943 & n12352 ) | ( n10372 & n12352 ) ;
  assign n12354 = n12352 | n12353 ;
  assign n12355 = ( n7929 & n10419 ) | ( n7929 & n12352 ) | ( n10419 & n12352 ) ;
  assign n12356 = n12354 | n12355 ;
  assign n12357 = ( n7930 & n12326 ) | ( n7930 & n12356 ) | ( n12326 & n12356 ) ;
  assign n12358 = n12356 | n12357 ;
  assign n12359 = n12358 ^ x8 ^ 1'b0 ;
  assign n12360 = n12350 ^ n12291 ^ n12283 ;
  assign n12361 = n12359 ^ n12324 ^ n12190 ;
  assign n12362 = ( n12190 & n12324 ) | ( n12190 & n12359 ) | ( n12324 & n12359 ) ;
  assign n12363 = n6901 & n10372 ;
  assign n12364 = ( n6906 & n10353 ) | ( n6906 & n12363 ) | ( n10353 & n12363 ) ;
  assign n12365 = n12363 | n12364 ;
  assign n12366 = ( n6907 & n10408 ) | ( n6907 & n12363 ) | ( n10408 & n12363 ) ;
  assign n12367 = n12365 | n12366 ;
  assign n12368 = ( n6918 & n12295 ) | ( n6918 & n12367 ) | ( n12295 & n12367 ) ;
  assign n12369 = n12367 | n12368 ;
  assign n12370 = n12369 ^ x29 ^ 1'b0 ;
  assign n12371 = ( n11327 & n12287 ) | ( n11327 & n12370 ) | ( n12287 & n12370 ) ;
  assign n12372 = n12370 ^ n12287 ^ n11327 ;
  assign n12373 = n8029 & n10372 ;
  assign n12374 = ( n8037 & n10353 ) | ( n8037 & n12373 ) | ( n10353 & n12373 ) ;
  assign n12375 = n12373 | n12374 ;
  assign n12376 = ( n8033 & n10408 ) | ( n8033 & n12373 ) | ( n10408 & n12373 ) ;
  assign n12377 = n12375 | n12376 ;
  assign n12378 = n8034 & n12295 ;
  assign n12379 = n12377 | n12378 ;
  assign n12380 = n12379 ^ x5 ^ 1'b0 ;
  assign n12381 = n12380 ^ n12049 ^ n11490 ;
  assign n12382 = ( n11490 & n12049 ) | ( n11490 & n12380 ) | ( n12049 & n12380 ) ;
  assign n12383 = n7485 & n10372 ;
  assign n12384 = ( n7486 & n10408 ) | ( n7486 & n12383 ) | ( n10408 & n12383 ) ;
  assign n12385 = n12383 | n12384 ;
  assign n12386 = ( n7493 & n10353 ) | ( n7493 & n12383 ) | ( n10353 & n12383 ) ;
  assign n12387 = n12385 | n12386 ;
  assign n12388 = n7487 & n12295 ;
  assign n12389 = n12387 | n12388 ;
  assign n12390 = n12389 ^ x17 ^ 1'b0 ;
  assign n12391 = n12390 ^ n12215 ^ n11869 ;
  assign n12392 = ( n11869 & n12215 ) | ( n11869 & n12390 ) | ( n12215 & n12390 ) ;
  assign n12393 = n7829 & n10372 ;
  assign n12394 = ( n7833 & n10353 ) | ( n7833 & n12393 ) | ( n10353 & n12393 ) ;
  assign n12395 = n12393 | n12394 ;
  assign n12396 = ( n7834 & n10408 ) | ( n7834 & n12393 ) | ( n10408 & n12393 ) ;
  assign n12397 = n12395 | n12396 ;
  assign n12398 = n7838 & n12295 ;
  assign n12399 = n12397 | n12398 ;
  assign n12400 = n12399 ^ x11 ^ 1'b0 ;
  assign n12401 = ( n12077 & n12245 ) | ( n12077 & n12400 ) | ( n12245 & n12400 ) ;
  assign n12402 = n12400 ^ n12245 ^ n12077 ;
  assign n12403 = n7188 & n10408 ;
  assign n12404 = ( n7190 & n10353 ) | ( n7190 & n12403 ) | ( n10353 & n12403 ) ;
  assign n12405 = n12403 | n12404 ;
  assign n12406 = ( n7192 & n10372 ) | ( n7192 & n12403 ) | ( n10372 & n12403 ) ;
  assign n12407 = n12405 | n12406 ;
  assign n12408 = n7196 & n12295 ;
  assign n12409 = n12407 | n12408 ;
  assign n12410 = n12289 ^ n12257 ^ n6775 ;
  assign n12411 = ( ~n6775 & n12257 ) | ( ~n6775 & n12289 ) | ( n12257 & n12289 ) ;
  assign n12412 = n12409 ^ x23 ^ 1'b0 ;
  assign n12413 = n12412 ^ n12225 ^ n12104 ;
  assign n12414 = ( ~n12104 & n12225 ) | ( ~n12104 & n12412 ) | ( n12225 & n12412 ) ;
  assign n12415 = n7339 & n10372 ;
  assign n12416 = ( n7337 & n10408 ) | ( n7337 & n12415 ) | ( n10408 & n12415 ) ;
  assign n12417 = n12415 | n12416 ;
  assign n12418 = ( n7338 & n10353 ) | ( n7338 & n12415 ) | ( n10353 & n12415 ) ;
  assign n12419 = n12417 | n12418 ;
  assign n12420 = ( n7340 & n12295 ) | ( n7340 & n12419 ) | ( n12295 & n12419 ) ;
  assign n12421 = n12419 | n12420 ;
  assign n12422 = n12421 ^ x20 ^ 1'b0 ;
  assign n12423 = n12422 ^ n12205 ^ n12117 ;
  assign n12424 = ( ~n12117 & n12205 ) | ( ~n12117 & n12422 ) | ( n12205 & n12422 ) ;
  assign n12425 = n6791 & n10372 ;
  assign n12426 = ( n6788 & n10408 ) | ( n6788 & n12425 ) | ( n10408 & n12425 ) ;
  assign n12427 = n12425 | n12426 ;
  assign n12428 = ( n6790 & n10353 ) | ( n6790 & n12425 ) | ( n10353 & n12425 ) ;
  assign n12429 = n12427 | n12428 ;
  assign n12430 = n6789 & ~n12295 ;
  assign n12431 = ( n6789 & n12429 ) | ( n6789 & ~n12430 ) | ( n12429 & ~n12430 ) ;
  assign n12432 = ( n12351 & ~n12410 ) | ( n12351 & n12431 ) | ( ~n12410 & n12431 ) ;
  assign n12433 = n12431 ^ n12410 ^ n12351 ;
  assign n12434 = n7037 & n10408 ;
  assign n12435 = ( n7036 & n10372 ) | ( n7036 & n12434 ) | ( n10372 & n12434 ) ;
  assign n12436 = n12434 | n12435 ;
  assign n12437 = ( n7052 & n10353 ) | ( n7052 & n12434 ) | ( n10353 & n12434 ) ;
  assign n12438 = n12436 | n12437 ;
  assign n12439 = ( n7035 & n12295 ) | ( n7035 & n12438 ) | ( n12295 & n12438 ) ;
  assign n12440 = n12438 | n12439 ;
  assign n12441 = n12440 ^ x26 ^ 1'b0 ;
  assign n12442 = n12441 ^ n12256 ^ n12115 ;
  assign n12443 = ( n12115 & n12256 ) | ( n12115 & n12441 ) | ( n12256 & n12441 ) ;
  assign n12444 = n7339 & n10408 ;
  assign n12445 = ( n7338 & n10372 ) | ( n7338 & n12444 ) | ( n10372 & n12444 ) ;
  assign n12446 = ( n7337 & n10419 ) | ( n7337 & n12444 ) | ( n10419 & n12444 ) ;
  assign n12447 = n12444 | n12446 ;
  assign n12448 = n12445 | n12447 ;
  assign n12449 = ( n7340 & n12326 ) | ( n7340 & n12448 ) | ( n12326 & n12448 ) ;
  assign n12450 = n12448 | n12449 ;
  assign n12451 = n12450 ^ x20 ^ 1'b0 ;
  assign n12452 = ( ~n12159 & n12424 ) | ( ~n12159 & n12451 ) | ( n12424 & n12451 ) ;
  assign n12453 = n7485 & n10408 ;
  assign n12454 = ( n7493 & n10372 ) | ( n7493 & n12453 ) | ( n10372 & n12453 ) ;
  assign n12455 = ( n7486 & n10419 ) | ( n7486 & n12453 ) | ( n10419 & n12453 ) ;
  assign n12456 = n12453 | n12455 ;
  assign n12457 = n12454 | n12456 ;
  assign n12458 = ( n7487 & n12326 ) | ( n7487 & n12457 ) | ( n12326 & n12457 ) ;
  assign n12459 = n12457 | n12458 ;
  assign n12460 = n12459 ^ x17 ^ 1'b0 ;
  assign n12461 = ( n12196 & n12392 ) | ( n12196 & n12460 ) | ( n12392 & n12460 ) ;
  assign n12462 = n12460 ^ n12392 ^ n12196 ;
  assign n12463 = n7829 & n10408 ;
  assign n12464 = ( n7834 & n10419 ) | ( n7834 & n12463 ) | ( n10419 & n12463 ) ;
  assign n12465 = ( n7833 & n10372 ) | ( n7833 & n12463 ) | ( n10372 & n12463 ) ;
  assign n12466 = n12451 ^ n12424 ^ n12159 ;
  assign n12467 = n12463 | n12465 ;
  assign n12468 = n12464 | n12467 ;
  assign n12469 = ( n7838 & n12326 ) | ( n7838 & n12468 ) | ( n12326 & n12468 ) ;
  assign n12470 = n12468 | n12469 ;
  assign n12471 = n12470 ^ x11 ^ 1'b0 ;
  assign n12472 = ( n12194 & n12401 ) | ( n12194 & n12471 ) | ( n12401 & n12471 ) ;
  assign n12473 = n12471 ^ n12401 ^ n12194 ;
  assign n12474 = n8029 & n10408 ;
  assign n12475 = ( n8033 & n10419 ) | ( n8033 & n12474 ) | ( n10419 & n12474 ) ;
  assign n12476 = ( n8037 & n10372 ) | ( n8037 & n12474 ) | ( n10372 & n12474 ) ;
  assign n12477 = n12474 | n12476 ;
  assign n12478 = n12475 | n12477 ;
  assign n12479 = ( n8034 & n12326 ) | ( n8034 & n12478 ) | ( n12326 & n12478 ) ;
  assign n12480 = n12478 | n12479 ;
  assign n12481 = n12480 ^ x5 ^ 1'b0 ;
  assign n12482 = ( n12173 & n12382 ) | ( n12173 & n12481 ) | ( n12382 & n12481 ) ;
  assign n12483 = n12481 ^ n12382 ^ n12173 ;
  assign n12484 = n7196 & n12326 ;
  assign n12485 = n7188 & n10419 ;
  assign n12486 = ( n7192 & n10408 ) | ( n7192 & n12485 ) | ( n10408 & n12485 ) ;
  assign n12487 = ( n7190 & n10372 ) | ( n7190 & n12485 ) | ( n10372 & n12485 ) ;
  assign n12488 = n12485 | n12487 ;
  assign n12489 = n12486 | n12488 ;
  assign n12490 = n12484 | n12489 ;
  assign n12491 = n12490 ^ x23 ^ 1'b0 ;
  assign n12492 = n12491 ^ n12414 ^ n12148 ;
  assign n12493 = ( ~n12148 & n12414 ) | ( ~n12148 & n12491 ) | ( n12414 & n12491 ) ;
  assign n12494 = n7037 & n10419 ;
  assign n12495 = ( n7052 & n10372 ) | ( n7052 & n12494 ) | ( n10372 & n12494 ) ;
  assign n12496 = ( n7036 & n10408 ) | ( n7036 & n12494 ) | ( n10408 & n12494 ) ;
  assign n12497 = n12494 | n12496 ;
  assign n12498 = n12495 | n12497 ;
  assign n12499 = ( n7035 & n12326 ) | ( n7035 & n12498 ) | ( n12326 & n12498 ) ;
  assign n12500 = n12498 | n12499 ;
  assign n12501 = n12500 ^ x26 ^ 1'b0 ;
  assign n12502 = n12501 ^ n12443 ^ n12119 ;
  assign n12503 = ( n12119 & n12443 ) | ( n12119 & n12501 ) | ( n12443 & n12501 ) ;
  assign n12504 = n6789 & ~n12326 ;
  assign n12505 = n6791 & n10408 ;
  assign n12506 = ( n6790 & n10372 ) | ( n6790 & n12505 ) | ( n10372 & n12505 ) ;
  assign n12507 = ( n6788 & n10419 ) | ( n6788 & n12505 ) | ( n10419 & n12505 ) ;
  assign n12508 = n12505 | n12507 ;
  assign n12509 = n12506 | n12508 ;
  assign n12510 = ( n6789 & ~n12504 ) | ( n6789 & n12509 ) | ( ~n12504 & n12509 ) ;
  assign n12511 = n7188 & n10425 ;
  assign n12512 = ( n7190 & n10408 ) | ( n7190 & n12511 ) | ( n10408 & n12511 ) ;
  assign n12513 = ( n10408 & n10419 ) | ( n10408 & n12321 ) | ( n10419 & n12321 ) ;
  assign n12514 = n12513 ^ n10425 ^ n10419 ;
  assign n12515 = n12511 | n12512 ;
  assign n12516 = ( n7192 & n10419 ) | ( n7192 & n12511 ) | ( n10419 & n12511 ) ;
  assign n12517 = n12515 | n12516 ;
  assign n12518 = n7196 & n12514 ;
  assign n12519 = n12517 | n12518 ;
  assign n12520 = n12519 ^ x23 ^ 1'b0 ;
  assign n12521 = n12520 ^ n12493 ^ n12255 ;
  assign n12522 = ( n12255 & n12493 ) | ( n12255 & n12520 ) | ( n12493 & n12520 ) ;
  assign n12523 = n8086 & n10408 ;
  assign n12524 = ( n8088 & n10419 ) | ( n8088 & n12523 ) | ( n10419 & n12523 ) ;
  assign n12525 = n12523 | n12524 ;
  assign n12526 = ( n8090 & n10425 ) | ( n8090 & n12523 ) | ( n10425 & n12523 ) ;
  assign n12527 = n12525 | n12526 ;
  assign n12528 = ( n8089 & n12514 ) | ( n8089 & n12527 ) | ( n12514 & n12527 ) ;
  assign n12529 = n12527 | n12528 ;
  assign n12530 = n12529 ^ x2 ^ 1'b0 ;
  assign n12531 = ( n11489 & n12330 ) | ( n11489 & n12530 ) | ( n12330 & n12530 ) ;
  assign n12532 = n8086 & n10419 ;
  assign n12533 = ( n8090 & n10491 ) | ( n8090 & n12532 ) | ( n10491 & n12532 ) ;
  assign n12534 = ( n8088 & n10425 ) | ( n8088 & n12532 ) | ( n10425 & n12532 ) ;
  assign n12535 = n12532 | n12534 ;
  assign n12536 = n7037 & n10425 ;
  assign n12537 = n12533 | n12535 ;
  assign n12538 = ( n7036 & n10419 ) | ( n7036 & n12536 ) | ( n10419 & n12536 ) ;
  assign n12539 = n12536 | n12538 ;
  assign n12540 = ( n7052 & n10408 ) | ( n7052 & n12536 ) | ( n10408 & n12536 ) ;
  assign n12541 = n12539 | n12540 ;
  assign n12542 = ( n7035 & n12514 ) | ( n7035 & n12541 ) | ( n12514 & n12541 ) ;
  assign n12543 = n12541 | n12542 ;
  assign n12544 = n12543 ^ x26 ^ 1'b0 ;
  assign n12545 = n12544 ^ n12503 ^ n12285 ;
  assign n12546 = ( n12285 & n12503 ) | ( n12285 & n12544 ) | ( n12503 & n12544 ) ;
  assign n12547 = n8029 & n10419 ;
  assign n12548 = ( n8037 & n10408 ) | ( n8037 & n12547 ) | ( n10408 & n12547 ) ;
  assign n12549 = n12547 | n12548 ;
  assign n12550 = ( n8033 & n10425 ) | ( n8033 & n12547 ) | ( n10425 & n12547 ) ;
  assign n12551 = n12549 | n12550 ;
  assign n12552 = ( n8034 & n12514 ) | ( n8034 & n12551 ) | ( n12514 & n12551 ) ;
  assign n12553 = n12551 | n12552 ;
  assign n12554 = n12553 ^ x5 ^ 1'b0 ;
  assign n12555 = ( n12267 & n12482 ) | ( n12267 & n12554 ) | ( n12482 & n12554 ) ;
  assign n12556 = ( n10419 & n10425 ) | ( n10419 & n12513 ) | ( n10425 & n12513 ) ;
  assign n12557 = n12554 ^ n12482 ^ n12267 ;
  assign n12558 = n12556 ^ n10491 ^ n10425 ;
  assign n12559 = ( n8089 & n12537 ) | ( n8089 & n12558 ) | ( n12537 & n12558 ) ;
  assign n12560 = n12537 | n12559 ;
  assign n12561 = n12560 ^ x2 ^ 1'b0 ;
  assign n12562 = ( n12381 & n12531 ) | ( n12381 & n12561 ) | ( n12531 & n12561 ) ;
  assign n12563 = n8029 & n10425 ;
  assign n12564 = ( n8037 & n10419 ) | ( n8037 & n12563 ) | ( n10419 & n12563 ) ;
  assign n12565 = n12563 | n12564 ;
  assign n12566 = ( n8033 & n10491 ) | ( n8033 & n12563 ) | ( n10491 & n12563 ) ;
  assign n12567 = n12565 | n12566 ;
  assign n12568 = ( n8034 & n12558 ) | ( n8034 & n12567 ) | ( n12558 & n12567 ) ;
  assign n12569 = n12567 | n12568 ;
  assign n12570 = n12569 ^ x5 ^ 1'b0 ;
  assign n12571 = n12570 ^ n12555 ^ n12325 ;
  assign n12572 = ( n12325 & n12555 ) | ( n12325 & n12570 ) | ( n12555 & n12570 ) ;
  assign n12573 = n7037 & n10491 ;
  assign n12574 = ( n7052 & n10419 ) | ( n7052 & n12573 ) | ( n10419 & n12573 ) ;
  assign n12575 = ( n7036 & n10425 ) | ( n7036 & n12573 ) | ( n10425 & n12573 ) ;
  assign n12576 = n12573 | n12575 ;
  assign n12577 = n12574 | n12576 ;
  assign n12578 = ( n7035 & n12558 ) | ( n7035 & n12577 ) | ( n12558 & n12577 ) ;
  assign n12579 = n12577 | n12578 ;
  assign n12580 = n12579 ^ x26 ^ 1'b0 ;
  assign n12581 = ( n12372 & n12546 ) | ( n12372 & n12580 ) | ( n12546 & n12580 ) ;
  assign n12582 = n12580 ^ n12546 ^ n12372 ;
  assign n12583 = n7829 & n10419 ;
  assign n12584 = n7669 & n10419 ;
  assign n12585 = ( n7667 & n10425 ) | ( n7667 & n12584 ) | ( n10425 & n12584 ) ;
  assign n12586 = ( n7674 & n10408 ) | ( n7674 & n12584 ) | ( n10408 & n12584 ) ;
  assign n12587 = n12584 | n12586 ;
  assign n12588 = n7339 & n10419 ;
  assign n12589 = n12585 | n12587 ;
  assign n12590 = ( n7337 & n10425 ) | ( n7337 & n12588 ) | ( n10425 & n12588 ) ;
  assign n12591 = n12588 | n12590 ;
  assign n12592 = ( n7338 & n10408 ) | ( n7338 & n12588 ) | ( n10408 & n12588 ) ;
  assign n12593 = n12591 | n12592 ;
  assign n12594 = ( n7666 & n12514 ) | ( n7666 & n12589 ) | ( n12514 & n12589 ) ;
  assign n12595 = n12589 | n12594 ;
  assign n12596 = ( n7833 & n10408 ) | ( n7833 & n12583 ) | ( n10408 & n12583 ) ;
  assign n12597 = n12583 | n12596 ;
  assign n12598 = n12595 ^ x14 ^ 1'b0 ;
  assign n12599 = ( n7834 & n10425 ) | ( n7834 & n12583 ) | ( n10425 & n12583 ) ;
  assign n12600 = n12597 | n12599 ;
  assign n12601 = ( n12216 & n12344 ) | ( n12216 & n12598 ) | ( n12344 & n12598 ) ;
  assign n12602 = n12598 ^ n12344 ^ n12216 ;
  assign n12603 = ( n7340 & n12514 ) | ( n7340 & n12593 ) | ( n12514 & n12593 ) ;
  assign n12604 = n12593 | n12603 ;
  assign n12605 = n12604 ^ x20 ^ 1'b0 ;
  assign n12606 = ( n12226 & n12452 ) | ( n12226 & n12605 ) | ( n12452 & n12605 ) ;
  assign n12607 = ( n7838 & n12514 ) | ( n7838 & n12600 ) | ( n12514 & n12600 ) ;
  assign n12608 = n12600 | n12607 ;
  assign n12609 = n7485 & n10419 ;
  assign n12610 = n12605 ^ n12452 ^ n12226 ;
  assign n12611 = ( n7493 & n10408 ) | ( n7493 & n12609 ) | ( n10408 & n12609 ) ;
  assign n12612 = ( n7486 & n10425 ) | ( n7486 & n12609 ) | ( n10425 & n12609 ) ;
  assign n12613 = n12609 | n12612 ;
  assign n12614 = n6901 & n10419 ;
  assign n12615 = n12611 | n12613 ;
  assign n12616 = ( n6906 & n10408 ) | ( n6906 & n12614 ) | ( n10408 & n12614 ) ;
  assign n12617 = n12614 | n12616 ;
  assign n12618 = n12608 ^ x11 ^ 1'b0 ;
  assign n12619 = ( n6907 & n10425 ) | ( n6907 & n12614 ) | ( n10425 & n12614 ) ;
  assign n12620 = n12617 | n12619 ;
  assign n12621 = n12618 ^ n12472 ^ n12236 ;
  assign n12622 = ( n12236 & n12472 ) | ( n12236 & n12618 ) | ( n12472 & n12618 ) ;
  assign n12623 = ( n7487 & n12514 ) | ( n7487 & n12615 ) | ( n12514 & n12615 ) ;
  assign n12624 = n12615 | n12623 ;
  assign n12625 = n7932 & n10419 ;
  assign n12626 = ( n7943 & n10408 ) | ( n7943 & n12625 ) | ( n10408 & n12625 ) ;
  assign n12627 = n12625 | n12626 ;
  assign n12628 = ( n7929 & n10425 ) | ( n7929 & n12625 ) | ( n10425 & n12625 ) ;
  assign n12629 = n12624 ^ x17 ^ 1'b0 ;
  assign n12630 = n12627 | n12628 ;
  assign n12631 = n12629 ^ n12461 ^ n12206 ;
  assign n12632 = ( n12206 & n12461 ) | ( n12206 & n12629 ) | ( n12461 & n12629 ) ;
  assign n12633 = n6789 & n12514 ;
  assign n12634 = n6918 & n12514 ;
  assign n12635 = n12620 | n12634 ;
  assign n12636 = n7932 & n10425 ;
  assign n12637 = ( n6790 & n10408 ) | ( n6790 & n12633 ) | ( n10408 & n12633 ) ;
  assign n12638 = ( n7930 & n12514 ) | ( n7930 & n12630 ) | ( n12514 & n12630 ) ;
  assign n12639 = n12630 | n12638 ;
  assign n12640 = ( n6791 & n10419 ) | ( n6791 & n12633 ) | ( n10419 & n12633 ) ;
  assign n12641 = n12633 | n12640 ;
  assign n12642 = n12639 ^ x8 ^ 1'b0 ;
  assign n12643 = ( n7943 & n10419 ) | ( n7943 & n12636 ) | ( n10419 & n12636 ) ;
  assign n12644 = n12636 | n12643 ;
  assign n12645 = ( n7929 & n10491 ) | ( n7929 & n12636 ) | ( n10491 & n12636 ) ;
  assign n12646 = n12644 | n12645 ;
  assign n12647 = ( n7930 & n12558 ) | ( n7930 & n12646 ) | ( n12558 & n12646 ) ;
  assign n12648 = n12646 | n12647 ;
  assign n12649 = n12637 | n12641 ;
  assign n12650 = n12648 ^ x8 ^ 1'b0 ;
  assign n12651 = ( n12246 & n12362 ) | ( n12246 & n12642 ) | ( n12362 & n12642 ) ;
  assign n12652 = n12651 ^ n12650 ^ n12402 ;
  assign n12653 = ( n12402 & n12650 ) | ( n12402 & n12651 ) | ( n12650 & n12651 ) ;
  assign n12654 = n12642 ^ n12362 ^ n12246 ;
  assign n12655 = n8030 ^ x5 ^ 1'b0 ;
  assign n12656 = n12655 ^ n12257 ^ n6684 ;
  assign n12657 = ( n6684 & n12257 ) | ( n6684 & n12655 ) | ( n12257 & n12655 ) ;
  assign n12658 = ( n10425 & n10491 ) | ( n10425 & n12556 ) | ( n10491 & n12556 ) ;
  assign n12659 = n8086 & n10425 ;
  assign n12660 = ( n8088 & n10491 ) | ( n8088 & n12659 ) | ( n10491 & n12659 ) ;
  assign n12661 = n12659 | n12660 ;
  assign n12662 = ( n8090 & n10492 ) | ( n8090 & n12659 ) | ( n10492 & n12659 ) ;
  assign n12663 = n12661 | n12662 ;
  assign n12664 = ( n12411 & n12510 ) | ( n12411 & ~n12656 ) | ( n12510 & ~n12656 ) ;
  assign n12665 = n12656 ^ n12510 ^ n12411 ;
  assign n12666 = n7669 & n10425 ;
  assign n12667 = ( n7674 & n10419 ) | ( n7674 & n12666 ) | ( n10419 & n12666 ) ;
  assign n12668 = n12666 | n12667 ;
  assign n12669 = ( n7667 & n10491 ) | ( n7667 & n12666 ) | ( n10491 & n12666 ) ;
  assign n12670 = n12668 | n12669 ;
  assign n12671 = ( n7666 & n12558 ) | ( n7666 & n12670 ) | ( n12558 & n12670 ) ;
  assign n12672 = n12670 | n12671 ;
  assign n12673 = n12672 ^ x14 ^ 1'b0 ;
  assign n12674 = ( n12391 & n12601 ) | ( n12391 & n12673 ) | ( n12601 & n12673 ) ;
  assign n12675 = n12673 ^ n12601 ^ n12391 ;
  assign n12676 = ( n10491 & n10492 ) | ( n10491 & n12658 ) | ( n10492 & n12658 ) ;
  assign n12677 = n12658 ^ n10492 ^ n10491 ;
  assign n12678 = n8089 & n12677 ;
  assign n12679 = n12663 | n12678 ;
  assign n12680 = n12679 ^ x2 ^ 1'b0 ;
  assign n12681 = ( n12483 & n12562 ) | ( n12483 & n12680 ) | ( n12562 & n12680 ) ;
  assign n12682 = n6788 & ~n10425 ;
  assign n12683 = ( n6788 & n12649 ) | ( n6788 & ~n12682 ) | ( n12649 & ~n12682 ) ;
  assign n12684 = ( n6714 & n12657 ) | ( n6714 & ~n12683 ) | ( n12657 & ~n12683 ) ;
  assign n12685 = n7339 & n10425 ;
  assign n12686 = ( n7337 & n10491 ) | ( n7337 & n12685 ) | ( n10491 & n12685 ) ;
  assign n12687 = n12685 | n12686 ;
  assign n12688 = n12683 ^ n12657 ^ n6714 ;
  assign n12689 = ( n7338 & n10419 ) | ( n7338 & n12685 ) | ( n10419 & n12685 ) ;
  assign n12690 = n12687 | n12689 ;
  assign n12691 = ( n7340 & n12558 ) | ( n7340 & n12690 ) | ( n12558 & n12690 ) ;
  assign n12692 = ( n6711 & n6714 ) | ( n6711 & n12684 ) | ( n6714 & n12684 ) ;
  assign n12693 = n12690 | n12691 ;
  assign n12694 = n12693 ^ x20 ^ 1'b0 ;
  assign n12695 = n12694 ^ n12606 ^ n12413 ;
  assign n12696 = ( ~n12413 & n12606 ) | ( ~n12413 & n12694 ) | ( n12606 & n12694 ) ;
  assign n12697 = n12684 ^ n6714 ^ n6711 ;
  assign n12698 = n8086 & n10491 ;
  assign n12699 = ( n8088 & n10492 ) | ( n8088 & n12698 ) | ( n10492 & n12698 ) ;
  assign n12700 = ( n8090 & ~n10539 ) | ( n8090 & n12698 ) | ( ~n10539 & n12698 ) ;
  assign n12701 = n12698 | n12699 ;
  assign n12702 = n12700 | n12701 ;
  assign n12703 = n12676 ^ n10539 ^ n10492 ;
  assign n12704 = n8089 & ~n12703 ;
  assign n12705 = n12702 | n12704 ;
  assign n12706 = n12705 ^ x2 ^ 1'b0 ;
  assign n12707 = ( n12557 & n12681 ) | ( n12557 & n12706 ) | ( n12681 & n12706 ) ;
  assign n12708 = n7487 & n12558 ;
  assign n12709 = n7485 & n10425 ;
  assign n12710 = ( n7486 & n10491 ) | ( n7486 & n12709 ) | ( n10491 & n12709 ) ;
  assign n12711 = n12709 | n12710 ;
  assign n12712 = ( n7493 & n10419 ) | ( n7493 & n12709 ) | ( n10419 & n12709 ) ;
  assign n12713 = n12711 | n12712 ;
  assign n12714 = n12708 | n12713 ;
  assign n12715 = n12714 ^ x17 ^ 1'b0 ;
  assign n12716 = n6791 & n10425 ;
  assign n12717 = ( ~n12423 & n12632 ) | ( ~n12423 & n12715 ) | ( n12632 & n12715 ) ;
  assign n12718 = n12715 ^ n12632 ^ n12423 ;
  assign n12719 = ( n6788 & n10491 ) | ( n6788 & n12716 ) | ( n10491 & n12716 ) ;
  assign n12720 = n12716 | n12719 ;
  assign n12721 = n6901 & n10492 ;
  assign n12722 = ( n6790 & n10419 ) | ( n6790 & n12716 ) | ( n10419 & n12716 ) ;
  assign n12723 = n12720 | n12722 ;
  assign n12724 = ( n6906 & n10491 ) | ( n6906 & n12721 ) | ( n10491 & n12721 ) ;
  assign n12725 = n12721 | n12724 ;
  assign n12726 = ( n6907 & ~n10539 ) | ( n6907 & n12721 ) | ( ~n10539 & n12721 ) ;
  assign n12727 = n12725 | n12726 ;
  assign n12728 = n6918 & ~n12703 ;
  assign n12729 = n12727 & ~n12728 ;
  assign n12730 = n12729 ^ n12728 ^ x29 ;
  assign n12731 = n12730 ^ n12688 ^ n12664 ;
  assign n12732 = ( n12664 & n12688 ) | ( n12664 & n12730 ) | ( n12688 & n12730 ) ;
  assign n12733 = n6789 & ~n12558 ;
  assign n12734 = ( n6789 & n12723 ) | ( n6789 & ~n12733 ) | ( n12723 & ~n12733 ) ;
  assign n12735 = ( ~n12697 & n12732 ) | ( ~n12697 & n12734 ) | ( n12732 & n12734 ) ;
  assign n12736 = n12734 ^ n12732 ^ n12697 ;
  assign n12737 = n7829 & n10425 ;
  assign n12738 = ( n7834 & n10491 ) | ( n7834 & n12737 ) | ( n10491 & n12737 ) ;
  assign n12739 = ( n7833 & n10419 ) | ( n7833 & n12737 ) | ( n10419 & n12737 ) ;
  assign n12740 = n12737 | n12739 ;
  assign n12741 = n12738 | n12740 ;
  assign n12742 = n8086 & n10492 ;
  assign n12743 = ( n7838 & n12558 ) | ( n7838 & n12741 ) | ( n12558 & n12741 ) ;
  assign n12744 = n12741 | n12743 ;
  assign n12745 = ( n8088 & ~n10539 ) | ( n8088 & n12742 ) | ( ~n10539 & n12742 ) ;
  assign n12746 = ( n10492 & ~n10539 ) | ( n10492 & n12676 ) | ( ~n10539 & n12676 ) ;
  assign n12747 = n12742 | n12745 ;
  assign n12748 = ( n8090 & n10555 ) | ( n8090 & n12742 ) | ( n10555 & n12742 ) ;
  assign n12749 = n12747 | n12748 ;
  assign n12750 = n12744 ^ x11 ^ 1'b0 ;
  assign n12751 = n12750 ^ n12622 ^ n12316 ;
  assign n12752 = ( n12316 & n12622 ) | ( n12316 & n12750 ) | ( n12622 & n12750 ) ;
  assign n12753 = n12746 ^ n10555 ^ n10539 ;
  assign n12754 = n8089 & ~n12753 ;
  assign n12755 = n12749 | n12754 ;
  assign n12756 = n12755 ^ x2 ^ 1'b0 ;
  assign n12757 = ( n12571 & n12707 ) | ( n12571 & n12756 ) | ( n12707 & n12756 ) ;
  assign n12758 = n7188 & n10491 ;
  assign n12759 = ( n7190 & n10419 ) | ( n7190 & n12758 ) | ( n10419 & n12758 ) ;
  assign n12760 = n12758 | n12759 ;
  assign n12761 = n6901 & n10425 ;
  assign n12762 = ( n6906 & n10419 ) | ( n6906 & n12761 ) | ( n10419 & n12761 ) ;
  assign n12763 = n12761 | n12762 ;
  assign n12764 = ( n6907 & n10491 ) | ( n6907 & n12761 ) | ( n10491 & n12761 ) ;
  assign n12765 = ( n7192 & n10425 ) | ( n7192 & n12758 ) | ( n10425 & n12758 ) ;
  assign n12766 = n12760 | n12765 ;
  assign n12767 = n7196 & n12558 ;
  assign n12768 = n12763 | n12764 ;
  assign n12769 = n7188 & n10492 ;
  assign n12770 = n12766 | n12767 ;
  assign n12771 = ( n7190 & n10425 ) | ( n7190 & n12769 ) | ( n10425 & n12769 ) ;
  assign n12772 = n12769 | n12771 ;
  assign n12773 = ( n7192 & n10491 ) | ( n7192 & n12769 ) | ( n10491 & n12769 ) ;
  assign n12774 = n6918 & n12558 ;
  assign n12775 = n12768 | n12774 ;
  assign n12776 = n7188 & n10555 ;
  assign n12777 = n12772 | n12773 ;
  assign n12778 = ( n7190 & n10492 ) | ( n7190 & n12776 ) | ( n10492 & n12776 ) ;
  assign n12779 = n12776 | n12778 ;
  assign n12780 = ( n7192 & ~n10539 ) | ( n7192 & n12776 ) | ( ~n10539 & n12776 ) ;
  assign n12781 = n12779 | n12780 ;
  assign n12782 = n12770 ^ x23 ^ 1'b0 ;
  assign n12783 = ( n12442 & n12522 ) | ( n12442 & n12782 ) | ( n12522 & n12782 ) ;
  assign n12784 = n12782 ^ n12522 ^ n12442 ;
  assign n12785 = n7196 & n12677 ;
  assign n12786 = n12777 | n12785 ;
  assign n12787 = n7196 & ~n12753 ;
  assign n12788 = n12781 | n12787 ;
  assign n12789 = n12786 ^ x23 ^ 1'b0 ;
  assign n12790 = ( ~n10539 & n10555 ) | ( ~n10539 & n12746 ) | ( n10555 & n12746 ) ;
  assign n12791 = ( n12502 & n12783 ) | ( n12502 & n12789 ) | ( n12783 & n12789 ) ;
  assign n12792 = n12789 ^ n12783 ^ n12502 ;
  assign n12793 = n7188 & ~n10539 ;
  assign n12794 = ( n7190 & n10491 ) | ( n7190 & n12793 ) | ( n10491 & n12793 ) ;
  assign n12795 = n12788 ^ x23 ^ 1'b0 ;
  assign n12796 = n12793 | n12794 ;
  assign n12797 = ( n7192 & n10492 ) | ( n7192 & n12793 ) | ( n10492 & n12793 ) ;
  assign n12798 = n12796 | n12797 ;
  assign n12799 = n7196 & ~n12703 ;
  assign n12800 = n12798 | n12799 ;
  assign n12801 = n12800 ^ x23 ^ 1'b0 ;
  assign n12802 = ( n12545 & n12791 ) | ( n12545 & n12801 ) | ( n12791 & n12801 ) ;
  assign n12803 = n12802 ^ n12795 ^ n12582 ;
  assign n12804 = n12801 ^ n12791 ^ n12545 ;
  assign n12805 = ( n12582 & n12795 ) | ( n12582 & n12802 ) | ( n12795 & n12802 ) ;
  assign n12806 = n7829 & n10491 ;
  assign n12807 = ( n7833 & n10425 ) | ( n7833 & n12806 ) | ( n10425 & n12806 ) ;
  assign n12808 = n12806 | n12807 ;
  assign n12809 = ( n7834 & n10492 ) | ( n7834 & n12806 ) | ( n10492 & n12806 ) ;
  assign n12810 = n12808 | n12809 ;
  assign n12811 = n7838 & n12677 ;
  assign n12812 = n12810 | n12811 ;
  assign n12813 = n12812 ^ x11 ^ 1'b0 ;
  assign n12814 = n12813 ^ n12752 ^ n12345 ;
  assign n12815 = ( n12345 & n12752 ) | ( n12345 & n12813 ) | ( n12752 & n12813 ) ;
  assign n12816 = n7669 & n10491 ;
  assign n12817 = ( n7674 & n10425 ) | ( n7674 & n12816 ) | ( n10425 & n12816 ) ;
  assign n12818 = n12816 | n12817 ;
  assign n12819 = ( n7667 & n10492 ) | ( n7667 & n12816 ) | ( n10492 & n12816 ) ;
  assign n12820 = n12818 | n12819 ;
  assign n12821 = n7666 & n12677 ;
  assign n12822 = n12820 | n12821 ;
  assign n12823 = n12822 ^ x14 ^ 1'b0 ;
  assign n12824 = ( n12462 & n12674 ) | ( n12462 & n12823 ) | ( n12674 & n12823 ) ;
  assign n12825 = n12823 ^ n12674 ^ n12462 ;
  assign n12826 = n7339 & n10491 ;
  assign n12827 = ( n7337 & n10492 ) | ( n7337 & n12826 ) | ( n10492 & n12826 ) ;
  assign n12828 = n12826 | n12827 ;
  assign n12829 = ( n7338 & n10425 ) | ( n7338 & n12826 ) | ( n10425 & n12826 ) ;
  assign n12830 = n12828 | n12829 ;
  assign n12831 = ( n7340 & n12677 ) | ( n7340 & n12830 ) | ( n12677 & n12830 ) ;
  assign n12832 = n12830 | n12831 ;
  assign n12833 = n12832 ^ x20 ^ 1'b0 ;
  assign n12834 = n12833 ^ n12696 ^ n12492 ;
  assign n12835 = ( ~n12492 & n12696 ) | ( ~n12492 & n12833 ) | ( n12696 & n12833 ) ;
  assign n12836 = n8029 & n10491 ;
  assign n12837 = ( n8037 & n10425 ) | ( n8037 & n12836 ) | ( n10425 & n12836 ) ;
  assign n12838 = n12836 | n12837 ;
  assign n12839 = ( n8033 & n10492 ) | ( n8033 & n12836 ) | ( n10492 & n12836 ) ;
  assign n12840 = n12838 | n12839 ;
  assign n12841 = n8034 & n12677 ;
  assign n12842 = n12840 | n12841 ;
  assign n12843 = n12842 ^ x5 ^ 1'b0 ;
  assign n12844 = ( n12361 & n12572 ) | ( n12361 & n12843 ) | ( n12572 & n12843 ) ;
  assign n12845 = n12843 ^ n12572 ^ n12361 ;
  assign n12846 = n7485 & n10491 ;
  assign n12847 = ( n7486 & n10492 ) | ( n7486 & n12846 ) | ( n10492 & n12846 ) ;
  assign n12848 = n12846 | n12847 ;
  assign n12849 = ( n7493 & n10425 ) | ( n7493 & n12846 ) | ( n10425 & n12846 ) ;
  assign n12850 = n12848 | n12849 ;
  assign n12851 = n7487 & n12677 ;
  assign n12852 = n12850 | n12851 ;
  assign n12853 = n12852 ^ x17 ^ 1'b0 ;
  assign n12854 = n12853 ^ n12717 ^ n12466 ;
  assign n12855 = ( ~n12466 & n12717 ) | ( ~n12466 & n12853 ) | ( n12717 & n12853 ) ;
  assign n12856 = n7932 & n10491 ;
  assign n12857 = ( n7943 & n10425 ) | ( n7943 & n12856 ) | ( n10425 & n12856 ) ;
  assign n12858 = n12856 | n12857 ;
  assign n12859 = ( n7929 & n10492 ) | ( n7929 & n12856 ) | ( n10492 & n12856 ) ;
  assign n12860 = n12858 | n12859 ;
  assign n12861 = n7930 & n12677 ;
  assign n12862 = n12860 | n12861 ;
  assign n12863 = n12862 ^ x8 ^ 1'b0 ;
  assign n12864 = n12863 ^ n12653 ^ n12473 ;
  assign n12865 = ( n12473 & n12653 ) | ( n12473 & n12863 ) | ( n12653 & n12863 ) ;
  assign n12866 = n7829 & n10492 ;
  assign n12867 = ( n7833 & n10491 ) | ( n7833 & n12866 ) | ( n10491 & n12866 ) ;
  assign n12868 = n12866 | n12867 ;
  assign n12869 = ( n7834 & ~n10539 ) | ( n7834 & n12866 ) | ( ~n10539 & n12866 ) ;
  assign n12870 = n12868 | n12869 ;
  assign n12871 = n7838 & ~n12703 ;
  assign n12872 = n12870 | n12871 ;
  assign n12873 = n12872 ^ x11 ^ 1'b0 ;
  assign n12874 = ( n12602 & n12815 ) | ( n12602 & n12873 ) | ( n12815 & n12873 ) ;
  assign n12875 = n12873 ^ n12815 ^ n12602 ;
  assign n12876 = n6791 & n10491 ;
  assign n12877 = ( n6788 & n10492 ) | ( n6788 & n12876 ) | ( n10492 & n12876 ) ;
  assign n12878 = n12876 | n12877 ;
  assign n12879 = ( n6790 & n10425 ) | ( n6790 & n12876 ) | ( n10425 & n12876 ) ;
  assign n12880 = n12878 | n12879 ;
  assign n12881 = n6789 & ~n12677 ;
  assign n12882 = ( n6789 & n12880 ) | ( n6789 & ~n12881 ) | ( n12880 & ~n12881 ) ;
  assign n12883 = n7942 ^ x8 ^ 1'b0 ;
  assign n12884 = ( n6566 & ~n6714 ) | ( n6566 & n12883 ) | ( ~n6714 & n12883 ) ;
  assign n12885 = n12883 ^ n6714 ^ n6566 ;
  assign n12886 = n12885 ^ n12882 ^ n12692 ;
  assign n12887 = ( ~n12692 & n12882 ) | ( ~n12692 & n12885 ) | ( n12882 & n12885 ) ;
  assign n12888 = n7037 & n10492 ;
  assign n12889 = ( n7036 & n10491 ) | ( n7036 & n12888 ) | ( n10491 & n12888 ) ;
  assign n12890 = n12888 | n12889 ;
  assign n12891 = ( n7052 & n10425 ) | ( n7052 & n12888 ) | ( n10425 & n12888 ) ;
  assign n12892 = n12890 | n12891 ;
  assign n12893 = n6918 & n12677 ;
  assign n12894 = n7035 & n12677 ;
  assign n12895 = n12892 | n12894 ;
  assign n12896 = n12895 ^ x26 ^ 1'b0 ;
  assign n12897 = n12896 ^ n12371 ^ n12349 ;
  assign n12898 = ( ~n12349 & n12371 ) | ( ~n12349 & n12896 ) | ( n12371 & n12896 ) ;
  assign n12899 = n7339 & n10492 ;
  assign n12900 = ( n7337 & ~n10539 ) | ( n7337 & n12899 ) | ( ~n10539 & n12899 ) ;
  assign n12901 = n12899 | n12900 ;
  assign n12902 = ( n7338 & n10491 ) | ( n7338 & n12899 ) | ( n10491 & n12899 ) ;
  assign n12903 = n12901 | n12902 ;
  assign n12904 = n7340 & ~n12703 ;
  assign n12905 = n12903 & ~n12904 ;
  assign n12906 = n12905 ^ n12904 ^ x20 ;
  assign n12907 = ( n12521 & n12835 ) | ( n12521 & n12906 ) | ( n12835 & n12906 ) ;
  assign n12908 = n12906 ^ n12835 ^ n12521 ;
  assign n12909 = n6901 & n10491 ;
  assign n12910 = ( n6906 & n10425 ) | ( n6906 & n12909 ) | ( n10425 & n12909 ) ;
  assign n12911 = n12909 | n12910 ;
  assign n12912 = ( n6907 & n10492 ) | ( n6907 & n12909 ) | ( n10492 & n12909 ) ;
  assign n12913 = n12911 | n12912 ;
  assign n12914 = n12893 | n12913 ;
  assign n12915 = n12914 ^ x29 ^ 1'b0 ;
  assign n12916 = n12915 ^ n12665 ^ n12432 ;
  assign n12917 = ( n12432 & ~n12665 ) | ( n12432 & n12915 ) | ( ~n12665 & n12915 ) ;
  assign n12918 = n7485 & n10492 ;
  assign n12919 = ( n7486 & ~n10539 ) | ( n7486 & n12918 ) | ( ~n10539 & n12918 ) ;
  assign n12920 = n12918 | n12919 ;
  assign n12921 = ( n7493 & n10491 ) | ( n7493 & n12918 ) | ( n10491 & n12918 ) ;
  assign n12922 = n12920 | n12921 ;
  assign n12923 = n7487 & ~n12703 ;
  assign n12924 = n12922 | n12923 ;
  assign n12925 = n12924 ^ x17 ^ 1'b0 ;
  assign n12926 = n12925 ^ n12855 ^ n12610 ;
  assign n12927 = ( n12610 & n12855 ) | ( n12610 & n12925 ) | ( n12855 & n12925 ) ;
  assign n12928 = n8029 & n10492 ;
  assign n12929 = ( n8037 & n10491 ) | ( n8037 & n12928 ) | ( n10491 & n12928 ) ;
  assign n12930 = n12928 | n12929 ;
  assign n12931 = ( n8033 & ~n10539 ) | ( n8033 & n12928 ) | ( ~n10539 & n12928 ) ;
  assign n12932 = n12930 | n12931 ;
  assign n12933 = n8034 & ~n12703 ;
  assign n12934 = n12932 | n12933 ;
  assign n12935 = n12934 ^ x5 ^ 1'b0 ;
  assign n12936 = n12935 ^ n12844 ^ n12654 ;
  assign n12937 = ( n12654 & n12844 ) | ( n12654 & n12935 ) | ( n12844 & n12935 ) ;
  assign n12938 = n7037 & ~n10539 ;
  assign n12939 = ( n7036 & n10492 ) | ( n7036 & n12938 ) | ( n10492 & n12938 ) ;
  assign n12940 = n12938 | n12939 ;
  assign n12941 = ( n7052 & n10491 ) | ( n7052 & n12938 ) | ( n10491 & n12938 ) ;
  assign n12942 = n12940 | n12941 ;
  assign n12943 = n7035 & ~n12703 ;
  assign n12944 = n12942 | n12943 ;
  assign n12945 = n12944 ^ x26 ^ 1'b0 ;
  assign n12946 = n12635 ^ x29 ^ 1'b0 ;
  assign n12947 = ( n12360 & n12945 ) | ( n12360 & n12946 ) | ( n12945 & n12946 ) ;
  assign n12948 = n12946 ^ n12945 ^ n12360 ;
  assign n12949 = n7669 & n10492 ;
  assign n12950 = ( n7674 & n10491 ) | ( n7674 & n12949 ) | ( n10491 & n12949 ) ;
  assign n12951 = n12949 | n12950 ;
  assign n12952 = ( n7667 & ~n10539 ) | ( n7667 & n12949 ) | ( ~n10539 & n12949 ) ;
  assign n12953 = n12951 | n12952 ;
  assign n12954 = n7666 & ~n12703 ;
  assign n12955 = n12953 | n12954 ;
  assign n12956 = n12955 ^ x14 ^ 1'b0 ;
  assign n12957 = ( n12631 & n12824 ) | ( n12631 & n12956 ) | ( n12824 & n12956 ) ;
  assign n12958 = n12956 ^ n12824 ^ n12631 ;
  assign n12959 = n7932 & n10492 ;
  assign n12960 = ( n7943 & n10491 ) | ( n7943 & n12959 ) | ( n10491 & n12959 ) ;
  assign n12961 = n12959 | n12960 ;
  assign n12962 = ( n7929 & ~n10539 ) | ( n7929 & n12959 ) | ( ~n10539 & n12959 ) ;
  assign n12963 = n12961 | n12962 ;
  assign n12964 = n6789 & ~n12703 ;
  assign n12965 = n7930 & ~n12703 ;
  assign n12966 = ( n6790 & n10491 ) | ( n6790 & n12964 ) | ( n10491 & n12964 ) ;
  assign n12967 = n12963 | n12965 ;
  assign n12968 = ( n6791 & n10492 ) | ( n6791 & n12964 ) | ( n10492 & n12964 ) ;
  assign n12969 = n12964 | n12968 ;
  assign n12970 = n12967 ^ x8 ^ 1'b0 ;
  assign n12971 = ( n12621 & n12865 ) | ( n12621 & n12970 ) | ( n12865 & n12970 ) ;
  assign n12972 = n12970 ^ n12865 ^ n12621 ;
  assign n12973 = n8034 & ~n12753 ;
  assign n12974 = n8029 & ~n10539 ;
  assign n12975 = n12966 | n12969 ;
  assign n12976 = ( n8037 & n10492 ) | ( n8037 & n12974 ) | ( n10492 & n12974 ) ;
  assign n12977 = n12974 | n12976 ;
  assign n12978 = ( n8033 & n10555 ) | ( n8033 & n12974 ) | ( n10555 & n12974 ) ;
  assign n12979 = n12977 | n12978 ;
  assign n12980 = n12973 | n12979 ;
  assign n12981 = n12980 ^ x5 ^ 1'b0 ;
  assign n12982 = n12981 ^ n12937 ^ n12652 ;
  assign n12983 = ( n12652 & n12937 ) | ( n12652 & n12981 ) | ( n12937 & n12981 ) ;
  assign n12984 = n7932 & ~n10539 ;
  assign n12985 = n7930 & ~n12753 ;
  assign n12986 = ( n7943 & n10492 ) | ( n7943 & n12984 ) | ( n10492 & n12984 ) ;
  assign n12987 = n12984 | n12986 ;
  assign n12988 = ( n7929 & n10555 ) | ( n7929 & n12984 ) | ( n10555 & n12984 ) ;
  assign n12989 = n12987 | n12988 ;
  assign n12990 = n12985 | n12989 ;
  assign n12991 = n8086 & ~n10539 ;
  assign n12992 = n12990 ^ x8 ^ 1'b0 ;
  assign n12993 = ( n12751 & n12971 ) | ( n12751 & n12992 ) | ( n12971 & n12992 ) ;
  assign n12994 = n12992 ^ n12971 ^ n12751 ;
  assign n12995 = ( n8090 & ~n10669 ) | ( n8090 & n12991 ) | ( ~n10669 & n12991 ) ;
  assign n12996 = ( n8088 & n10555 ) | ( n8088 & n12991 ) | ( n10555 & n12991 ) ;
  assign n12997 = n12991 | n12996 ;
  assign n12998 = n12995 | n12997 ;
  assign n12999 = n7829 & ~n10539 ;
  assign n13000 = ( n7833 & n10492 ) | ( n7833 & n12999 ) | ( n10492 & n12999 ) ;
  assign n13001 = n12999 | n13000 ;
  assign n13002 = ( n7834 & n10555 ) | ( n7834 & n12999 ) | ( n10555 & n12999 ) ;
  assign n13003 = n13001 | n13002 ;
  assign n13004 = n7838 & ~n12753 ;
  assign n13005 = n13003 | n13004 ;
  assign n13006 = n13005 ^ x11 ^ 1'b0 ;
  assign n13007 = n13006 ^ n12874 ^ n12675 ;
  assign n13008 = ( n12675 & n12874 ) | ( n12675 & n13006 ) | ( n12874 & n13006 ) ;
  assign n13009 = n12790 ^ n10669 ^ n10555 ;
  assign n13010 = n8089 & ~n13009 ;
  assign n13011 = n12998 & ~n13010 ;
  assign n13012 = n13011 ^ n13010 ^ x2 ;
  assign n13013 = ( n12757 & n12845 ) | ( n12757 & n13012 ) | ( n12845 & n13012 ) ;
  assign n13014 = n7829 & n10555 ;
  assign n13015 = n7932 & n10555 ;
  assign n13016 = ( n7833 & ~n10539 ) | ( n7833 & n13014 ) | ( ~n10539 & n13014 ) ;
  assign n13017 = n13014 | n13016 ;
  assign n13018 = ( n7834 & ~n10669 ) | ( n7834 & n13014 ) | ( ~n10669 & n13014 ) ;
  assign n13019 = n13017 | n13018 ;
  assign n13020 = n7838 & ~n13009 ;
  assign n13021 = n13019 & ~n13020 ;
  assign n13022 = n13021 ^ n13020 ^ x11 ;
  assign n13023 = n13022 ^ n13008 ^ n12825 ;
  assign n13024 = ( n12825 & n13008 ) | ( n12825 & n13022 ) | ( n13008 & n13022 ) ;
  assign n13025 = ( n7943 & ~n10539 ) | ( n7943 & n13015 ) | ( ~n10539 & n13015 ) ;
  assign n13026 = n13015 | n13025 ;
  assign n13027 = n7669 & ~n10539 ;
  assign n13028 = ( n7929 & ~n10669 ) | ( n7929 & n13015 ) | ( ~n10669 & n13015 ) ;
  assign n13029 = n13026 | n13028 ;
  assign n13030 = n7930 & ~n13009 ;
  assign n13031 = n13029 & ~n13030 ;
  assign n13032 = n13031 ^ n13030 ^ x8 ;
  assign n13033 = n13032 ^ n12993 ^ n12814 ;
  assign n13034 = ( n12814 & n12993 ) | ( n12814 & n13032 ) | ( n12993 & n13032 ) ;
  assign n13035 = ( n7674 & n10492 ) | ( n7674 & n13027 ) | ( n10492 & n13027 ) ;
  assign n13036 = n13027 | n13035 ;
  assign n13037 = ( n7667 & n10555 ) | ( n7667 & n13027 ) | ( n10555 & n13027 ) ;
  assign n13038 = n13036 | n13037 ;
  assign n13039 = n7666 & ~n12753 ;
  assign n13040 = n13038 & ~n13039 ;
  assign n13041 = n13040 ^ n13039 ^ x14 ;
  assign n13042 = ( ~n12718 & n12957 ) | ( ~n12718 & n13041 ) | ( n12957 & n13041 ) ;
  assign n13043 = n13041 ^ n12957 ^ n12718 ;
  assign n13044 = n7037 & ~n10669 ;
  assign n13045 = ( n7036 & n10555 ) | ( n7036 & n13044 ) | ( n10555 & n13044 ) ;
  assign n13046 = n12775 ^ x29 ^ 1'b0 ;
  assign n13047 = n7188 & ~n10669 ;
  assign n13048 = n13044 | n13045 ;
  assign n13049 = ( n7052 & ~n10539 ) | ( n7052 & n13044 ) | ( ~n10539 & n13044 ) ;
  assign n13050 = n13048 | n13049 ;
  assign n13051 = ( n7190 & ~n10539 ) | ( n7190 & n13047 ) | ( ~n10539 & n13047 ) ;
  assign n13052 = n13047 | n13051 ;
  assign n13053 = ( n7192 & n10555 ) | ( n7192 & n13047 ) | ( n10555 & n13047 ) ;
  assign n13054 = n13052 | n13053 ;
  assign n13055 = n7196 & ~n13009 ;
  assign n13056 = n13054 | n13055 ;
  assign n13057 = n13056 ^ x23 ^ 1'b0 ;
  assign n13058 = n13057 ^ n12897 ^ n12581 ;
  assign n13059 = ( n12581 & ~n12897 ) | ( n12581 & n13057 ) | ( ~n12897 & n13057 ) ;
  assign n13060 = n7037 & n10555 ;
  assign n13061 = ( n7036 & ~n10539 ) | ( n7036 & n13060 ) | ( ~n10539 & n13060 ) ;
  assign n13062 = n13060 | n13061 ;
  assign n13063 = ( n7052 & n10492 ) | ( n7052 & n13060 ) | ( n10492 & n13060 ) ;
  assign n13064 = n13062 | n13063 ;
  assign n13065 = n7035 & ~n12753 ;
  assign n13066 = n13064 | n13065 ;
  assign n13067 = n13066 ^ x26 ^ 1'b0 ;
  assign n13068 = n6788 & ~n10539 ;
  assign n13069 = n12975 | n13068 ;
  assign n13070 = ( ~n12433 & n13046 ) | ( ~n12433 & n13067 ) | ( n13046 & n13067 ) ;
  assign n13071 = n13067 ^ n13046 ^ n12433 ;
  assign n13072 = n7035 & ~n13009 ;
  assign n13073 = n7485 & ~n10539 ;
  assign n13074 = n13050 | n13072 ;
  assign n13075 = ( n7486 & n10555 ) | ( n7486 & n13073 ) | ( n10555 & n13073 ) ;
  assign n13076 = n13073 | n13075 ;
  assign n13077 = ( n7493 & n10492 ) | ( n7493 & n13073 ) | ( n10492 & n13073 ) ;
  assign n13078 = n13076 | n13077 ;
  assign n13079 = n13074 ^ x26 ^ 1'b0 ;
  assign n13080 = n7487 & ~n12753 ;
  assign n13081 = n13078 | n13080 ;
  assign n13082 = n13081 ^ x17 ^ 1'b0 ;
  assign n13083 = ( ~n12695 & n12927 ) | ( ~n12695 & n13082 ) | ( n12927 & n13082 ) ;
  assign n13084 = n13082 ^ n12927 ^ n12695 ;
  assign n13085 = n13079 ^ n13070 ^ n12916 ;
  assign n13086 = ( ~n12916 & n13070 ) | ( ~n12916 & n13079 ) | ( n13070 & n13079 ) ;
  assign n13087 = n7339 & ~n10539 ;
  assign n13088 = ( n7337 & n10555 ) | ( n7337 & n13087 ) | ( n10555 & n13087 ) ;
  assign n13089 = n7340 & ~n12753 ;
  assign n13090 = n13087 | n13088 ;
  assign n13091 = ( n7338 & n10492 ) | ( n7338 & n13087 ) | ( n10492 & n13087 ) ;
  assign n13092 = n13090 | n13091 ;
  assign n13093 = ( n6777 & ~n12884 ) | ( n6777 & n13069 ) | ( ~n12884 & n13069 ) ;
  assign n13094 = ~n13089 & n13092 ;
  assign n13095 = n13094 ^ n13089 ^ x20 ;
  assign n13096 = n13095 ^ n12907 ^ n12784 ;
  assign n13097 = ( n12784 & n12907 ) | ( n12784 & n13095 ) | ( n12907 & n13095 ) ;
  assign n13098 = n7485 & n10555 ;
  assign n13099 = ( n7486 & ~n10669 ) | ( n7486 & n13098 ) | ( ~n10669 & n13098 ) ;
  assign n13100 = n13069 ^ n12884 ^ n6777 ;
  assign n13101 = ( n7493 & ~n10539 ) | ( n7493 & n13098 ) | ( ~n10539 & n13098 ) ;
  assign n13102 = n13098 | n13099 ;
  assign n13103 = n7487 & ~n13009 ;
  assign n13104 = n13101 | n13102 ;
  assign n13105 = n13103 | n13104 ;
  assign n13106 = n13105 ^ x17 ^ 1'b0 ;
  assign n13107 = n13106 ^ n13083 ^ n12834 ;
  assign n13108 = ( ~n12834 & n13083 ) | ( ~n12834 & n13106 ) | ( n13083 & n13106 ) ;
  assign n13109 = n7669 & n10555 ;
  assign n13110 = ( n7674 & ~n10539 ) | ( n7674 & n13109 ) | ( ~n10539 & n13109 ) ;
  assign n13111 = n13109 | n13110 ;
  assign n13112 = ( n7667 & ~n10669 ) | ( n7667 & n13109 ) | ( ~n10669 & n13109 ) ;
  assign n13113 = n13111 | n13112 ;
  assign n13114 = n7666 & ~n13009 ;
  assign n13115 = n13113 & ~n13114 ;
  assign n13116 = n13115 ^ n13114 ^ x14 ;
  assign n13117 = n13116 ^ n13042 ^ n12854 ;
  assign n13118 = ( ~n12854 & n13042 ) | ( ~n12854 & n13116 ) | ( n13042 & n13116 ) ;
  assign n13119 = n8029 & n10555 ;
  assign n13120 = ( n8037 & ~n10539 ) | ( n8037 & n13119 ) | ( ~n10539 & n13119 ) ;
  assign n13121 = n13119 | n13120 ;
  assign n13122 = ( n8033 & ~n10669 ) | ( n8033 & n13119 ) | ( ~n10669 & n13119 ) ;
  assign n13123 = n13121 | n13122 ;
  assign n13124 = n8034 & ~n13009 ;
  assign n13125 = n13123 & ~n13124 ;
  assign n13126 = n13125 ^ n13124 ^ x5 ;
  assign n13127 = ( n12864 & n12983 ) | ( n12864 & n13126 ) | ( n12983 & n13126 ) ;
  assign n13128 = n13126 ^ n12983 ^ n12864 ;
  assign n13129 = n6901 & n10555 ;
  assign n13130 = ( n6906 & ~n10539 ) | ( n6906 & n13129 ) | ( ~n10539 & n13129 ) ;
  assign n13131 = n13129 | n13130 ;
  assign n13132 = ( n6907 & ~n10669 ) | ( n6907 & n13129 ) | ( ~n10669 & n13129 ) ;
  assign n13133 = n13131 | n13132 ;
  assign n13134 = n6918 & ~n13009 ;
  assign n13135 = n13133 | n13134 ;
  assign n13136 = n13135 ^ x29 ^ 1'b0 ;
  assign n13137 = ( n12735 & ~n12886 ) | ( n12735 & n13136 ) | ( ~n12886 & n13136 ) ;
  assign n13138 = n13136 ^ n12886 ^ n12735 ;
  assign n13139 = n7339 & n10555 ;
  assign n13140 = ( n7337 & ~n10669 ) | ( n7337 & n13139 ) | ( ~n10669 & n13139 ) ;
  assign n13141 = n13139 | n13140 ;
  assign n13142 = ( n7338 & ~n10539 ) | ( n7338 & n13139 ) | ( ~n10539 & n13139 ) ;
  assign n13143 = n13141 | n13142 ;
  assign n13144 = n7340 & ~n13009 ;
  assign n13145 = n13143 & ~n13144 ;
  assign n13146 = n13145 ^ n13144 ^ x20 ;
  assign n13147 = n13146 ^ n13097 ^ n12792 ;
  assign n13148 = ( n12792 & n13097 ) | ( n12792 & n13146 ) | ( n13097 & n13146 ) ;
  assign n13149 = n6791 & ~n10539 ;
  assign n13150 = ( n6788 & n10555 ) | ( n6788 & n13149 ) | ( n10555 & n13149 ) ;
  assign n13151 = n13149 | n13150 ;
  assign n13152 = ( n6790 & n10492 ) | ( n6790 & n13149 ) | ( n10492 & n13149 ) ;
  assign n13153 = n13151 | n13152 ;
  assign n13154 = n6789 & ~n12753 ;
  assign n13155 = n13153 | n13154 ;
  assign n13156 = n6901 & ~n10539 ;
  assign n13157 = ( n6906 & n10492 ) | ( n6906 & n13156 ) | ( n10492 & n13156 ) ;
  assign n13158 = n13156 | n13157 ;
  assign n13159 = n7832 ^ x11 ^ 1'b0 ;
  assign n13160 = ( n6907 & n10555 ) | ( n6907 & n13156 ) | ( n10555 & n13156 ) ;
  assign n13161 = n6918 & ~n12753 ;
  assign n13162 = n6789 & ~n13009 ;
  assign n13163 = n13158 | n13160 ;
  assign n13164 = n13093 ^ n6777 ^ n6686 ;
  assign n13165 = ( ~n6686 & n6777 ) | ( ~n6686 & n13093 ) | ( n6777 & n13093 ) ;
  assign n13166 = n6791 & n10555 ;
  assign n13167 = n13161 | n13163 ;
  assign n13168 = ( n6788 & ~n10669 ) | ( n6788 & n13166 ) | ( ~n10669 & n13166 ) ;
  assign n13169 = n13166 | n13168 ;
  assign n13170 = ( n6790 & ~n10539 ) | ( n6790 & n13166 ) | ( ~n10539 & n13166 ) ;
  assign n13171 = n13159 ^ n6777 ^ n6393 ;
  assign n13172 = n13169 | n13170 ;
  assign n13173 = n13162 | n13172 ;
  assign n13174 = ( n6393 & n6777 ) | ( n6393 & n13159 ) | ( n6777 & n13159 ) ;
  assign n13175 = n13173 ^ n13171 ^ n13165 ;
  assign n13176 = ( n13165 & ~n13171 ) | ( n13165 & n13173 ) | ( ~n13171 & n13173 ) ;
  assign n13177 = n7932 & ~n10669 ;
  assign n13178 = ( n7943 & n10555 ) | ( n7943 & n13177 ) | ( n10555 & n13177 ) ;
  assign n13179 = ( n10555 & ~n10669 ) | ( n10555 & n12790 ) | ( ~n10669 & n12790 ) ;
  assign n13180 = n13177 | n13178 ;
  assign n13181 = n13179 ^ n10711 ^ n10669 ;
  assign n13182 = ( n7929 & n10711 ) | ( n7929 & n13177 ) | ( n10711 & n13177 ) ;
  assign n13183 = n13180 | n13182 ;
  assign n13184 = n7930 & ~n13181 ;
  assign n13185 = n13183 & ~n13184 ;
  assign n13186 = n13185 ^ n13184 ^ x8 ;
  assign n13187 = n13186 ^ n13034 ^ n12875 ;
  assign n13188 = ( n12875 & n13034 ) | ( n12875 & n13186 ) | ( n13034 & n13186 ) ;
  assign n13189 = n8086 & n10555 ;
  assign n13190 = ( n8088 & ~n10669 ) | ( n8088 & n13189 ) | ( ~n10669 & n13189 ) ;
  assign n13191 = n13189 | n13190 ;
  assign n13192 = ( n8090 & n10711 ) | ( n8090 & n13189 ) | ( n10711 & n13189 ) ;
  assign n13193 = n13191 | n13192 ;
  assign n13194 = n8089 & ~n13181 ;
  assign n13195 = n13193 & ~n13194 ;
  assign n13196 = n13195 ^ n13194 ^ x2 ;
  assign n13197 = ( n12936 & n13013 ) | ( n12936 & n13196 ) | ( n13013 & n13196 ) ;
  assign n13198 = n7037 & n10711 ;
  assign n13199 = n8029 & ~n10669 ;
  assign n13200 = ( n8037 & n10555 ) | ( n8037 & n13199 ) | ( n10555 & n13199 ) ;
  assign n13201 = n13199 | n13200 ;
  assign n13202 = ( n8033 & n10711 ) | ( n8033 & n13199 ) | ( n10711 & n13199 ) ;
  assign n13203 = n13201 | n13202 ;
  assign n13204 = n8034 & ~n13181 ;
  assign n13205 = n13203 & ~n13204 ;
  assign n13206 = n13205 ^ n13204 ^ x5 ;
  assign n13207 = ( n7036 & ~n10669 ) | ( n7036 & n13198 ) | ( ~n10669 & n13198 ) ;
  assign n13208 = n13198 | n13207 ;
  assign n13209 = ( n7052 & n10555 ) | ( n7052 & n13198 ) | ( n10555 & n13198 ) ;
  assign n13210 = n13208 | n13209 ;
  assign n13211 = n7035 & ~n13181 ;
  assign n13212 = n13210 | n13211 ;
  assign n13213 = n13206 ^ n13127 ^ n12972 ;
  assign n13214 = ( n12972 & n13127 ) | ( n12972 & n13206 ) | ( n13127 & n13206 ) ;
  assign n13215 = n13212 ^ x26 ^ 1'b0 ;
  assign n13216 = n13215 ^ n12917 ^ n12731 ;
  assign n13217 = ( ~n10669 & n10711 ) | ( ~n10669 & n13179 ) | ( n10711 & n13179 ) ;
  assign n13218 = ( n12731 & n12917 ) | ( n12731 & n13215 ) | ( n12917 & n13215 ) ;
  assign n13219 = n8086 & ~n10669 ;
  assign n13220 = ( n8088 & n10711 ) | ( n8088 & n13219 ) | ( n10711 & n13219 ) ;
  assign n13221 = n13219 | n13220 ;
  assign n13222 = ( n8090 & n10909 ) | ( n8090 & n13219 ) | ( n10909 & n13219 ) ;
  assign n13223 = n13221 | n13222 ;
  assign n13224 = n13217 ^ n10909 ^ n10711 ;
  assign n13225 = ( n8089 & n13223 ) | ( n8089 & n13224 ) | ( n13223 & n13224 ) ;
  assign n13226 = n13223 | n13225 ;
  assign n13227 = n13226 ^ x2 ^ 1'b0 ;
  assign n13228 = ( n12982 & n13197 ) | ( n12982 & n13227 ) | ( n13197 & n13227 ) ;
  assign n13229 = n7339 & ~n10669 ;
  assign n13230 = ( n7337 & n10711 ) | ( n7337 & n13229 ) | ( n10711 & n13229 ) ;
  assign n13231 = n13229 | n13230 ;
  assign n13232 = ( n7338 & n10555 ) | ( n7338 & n13229 ) | ( n10555 & n13229 ) ;
  assign n13233 = n7340 & ~n13181 ;
  assign n13234 = n13231 | n13232 ;
  assign n13235 = ~n13233 & n13234 ;
  assign n13236 = n7485 & ~n10669 ;
  assign n13237 = n13235 ^ n13233 ^ x20 ;
  assign n13238 = ( n12804 & n13148 ) | ( n12804 & n13237 ) | ( n13148 & n13237 ) ;
  assign n13239 = n13237 ^ n13148 ^ n12804 ;
  assign n13240 = ( n7486 & n10711 ) | ( n7486 & n13236 ) | ( n10711 & n13236 ) ;
  assign n13241 = n13236 | n13240 ;
  assign n13242 = ( n10711 & n10909 ) | ( n10711 & n13217 ) | ( n10909 & n13217 ) ;
  assign n13243 = n7487 & ~n13181 ;
  assign n13244 = ( n7493 & n10555 ) | ( n7493 & n13236 ) | ( n10555 & n13236 ) ;
  assign n13245 = n13241 | n13244 ;
  assign n13246 = n13243 | n13245 ;
  assign n13247 = n13246 ^ x17 ^ 1'b0 ;
  assign n13248 = n13247 ^ n13108 ^ n12908 ;
  assign n13249 = ( n12908 & n13108 ) | ( n12908 & n13247 ) | ( n13108 & n13247 ) ;
  assign n13250 = n7669 & ~n10669 ;
  assign n13251 = ( n7674 & n10555 ) | ( n7674 & n13250 ) | ( n10555 & n13250 ) ;
  assign n13252 = ( n7667 & n10711 ) | ( n7667 & n13250 ) | ( n10711 & n13250 ) ;
  assign n13253 = n13250 | n13251 ;
  assign n13254 = n13252 | n13253 ;
  assign n13255 = n7666 & ~n13181 ;
  assign n13256 = n13254 & ~n13255 ;
  assign n13257 = n13256 ^ n13255 ^ x14 ;
  assign n13258 = ( n12926 & n13118 ) | ( n12926 & n13257 ) | ( n13118 & n13257 ) ;
  assign n13259 = n8086 & n10711 ;
  assign n13260 = n13257 ^ n13118 ^ n12926 ;
  assign n13261 = ( n8088 & n10909 ) | ( n8088 & n13259 ) | ( n10909 & n13259 ) ;
  assign n13262 = ( n8090 & ~n10930 ) | ( n8090 & n13259 ) | ( ~n10930 & n13259 ) ;
  assign n13263 = n13259 | n13261 ;
  assign n13264 = n13262 | n13263 ;
  assign n13265 = n13242 ^ n10930 ^ n10909 ;
  assign n13266 = n8089 & ~n13265 ;
  assign n13267 = n13264 | n13266 ;
  assign n13268 = n6918 & ~n13181 ;
  assign n13269 = n13267 ^ x2 ^ 1'b0 ;
  assign n13270 = ( n13128 & n13228 ) | ( n13128 & n13269 ) | ( n13228 & n13269 ) ;
  assign n13271 = n6901 & ~n10669 ;
  assign n13272 = ( n6906 & n10555 ) | ( n6906 & n13271 ) | ( n10555 & n13271 ) ;
  assign n13273 = n13271 | n13272 ;
  assign n13274 = ( n6907 & n10711 ) | ( n6907 & n13271 ) | ( n10711 & n13271 ) ;
  assign n13275 = n13273 | n13274 ;
  assign n13276 = ~n13268 & n13275 ;
  assign n13277 = n13276 ^ n13268 ^ x29 ;
  assign n13278 = n7188 & n10711 ;
  assign n13279 = ( n7190 & n10555 ) | ( n7190 & n13278 ) | ( n10555 & n13278 ) ;
  assign n13280 = n13278 | n13279 ;
  assign n13281 = ( n7192 & ~n10669 ) | ( n7192 & n13278 ) | ( ~n10669 & n13278 ) ;
  assign n13282 = n13280 | n13281 ;
  assign n13283 = n13277 ^ n13100 ^ n12887 ;
  assign n13284 = ( n12887 & ~n13100 ) | ( n12887 & n13277 ) | ( ~n13100 & n13277 ) ;
  assign n13285 = n6789 & ~n13181 ;
  assign n13286 = ( n6791 & ~n10669 ) | ( n6791 & n13285 ) | ( ~n10669 & n13285 ) ;
  assign n13287 = n13285 | n13286 ;
  assign n13288 = ( n6790 & n10555 ) | ( n6790 & n13285 ) | ( n10555 & n13285 ) ;
  assign n13289 = n13287 | n13288 ;
  assign n13290 = n7838 & ~n13181 ;
  assign n13291 = n7196 & ~n13181 ;
  assign n13292 = n13282 | n13291 ;
  assign n13293 = n13292 ^ x23 ^ 1'b0 ;
  assign n13294 = ( n12898 & n12948 ) | ( n12898 & n13293 ) | ( n12948 & n13293 ) ;
  assign n13295 = n13293 ^ n12948 ^ n12898 ;
  assign n13296 = n6788 & ~n10711 ;
  assign n13297 = ( n6788 & n13289 ) | ( n6788 & ~n13296 ) | ( n13289 & ~n13296 ) ;
  assign n13298 = ( n10909 & ~n10930 ) | ( n10909 & n13242 ) | ( ~n10930 & n13242 ) ;
  assign n13299 = n7829 & ~n10669 ;
  assign n13300 = ( n7833 & n10555 ) | ( n7833 & n13299 ) | ( n10555 & n13299 ) ;
  assign n13301 = n13299 | n13300 ;
  assign n13302 = ( n7834 & n10711 ) | ( n7834 & n13299 ) | ( n10711 & n13299 ) ;
  assign n13303 = n13301 | n13302 ;
  assign n13304 = n8086 & n10909 ;
  assign n13305 = ~n13290 & n13303 ;
  assign n13306 = n13298 ^ n10930 ^ n10926 ;
  assign n13307 = n13305 ^ n13290 ^ x11 ;
  assign n13308 = ( n8088 & ~n10930 ) | ( n8088 & n13304 ) | ( ~n10930 & n13304 ) ;
  assign n13309 = n13304 | n13308 ;
  assign n13310 = ( n8090 & n10926 ) | ( n8090 & n13304 ) | ( n10926 & n13304 ) ;
  assign n13311 = n13309 | n13310 ;
  assign n13312 = n13307 ^ n13024 ^ n12958 ;
  assign n13313 = ( n12958 & n13024 ) | ( n12958 & n13307 ) | ( n13024 & n13307 ) ;
  assign n13314 = n8089 & ~n13306 ;
  assign n13315 = n13311 | n13314 ;
  assign n13316 = n13315 ^ x2 ^ 1'b0 ;
  assign n13317 = ( n13213 & n13270 ) | ( n13213 & n13316 ) | ( n13270 & n13316 ) ;
  assign n13318 = n7829 & n10711 ;
  assign n13319 = ( n7833 & ~n10669 ) | ( n7833 & n13318 ) | ( ~n10669 & n13318 ) ;
  assign n13320 = n13318 | n13319 ;
  assign n13321 = ( n7834 & n10909 ) | ( n7834 & n13318 ) | ( n10909 & n13318 ) ;
  assign n13322 = n13320 | n13321 ;
  assign n13323 = n7838 & n13224 ;
  assign n13324 = n13322 | n13323 ;
  assign n13325 = n13324 ^ x11 ^ 1'b0 ;
  assign n13326 = n13325 ^ n13313 ^ n13043 ;
  assign n13327 = ( ~n13043 & n13313 ) | ( ~n13043 & n13325 ) | ( n13313 & n13325 ) ;
  assign n13328 = n7188 & n10909 ;
  assign n13329 = ( n7190 & ~n10669 ) | ( n7190 & n13328 ) | ( ~n10669 & n13328 ) ;
  assign n13330 = n13328 | n13329 ;
  assign n13331 = ( n7192 & n10711 ) | ( n7192 & n13328 ) | ( n10711 & n13328 ) ;
  assign n13332 = n13330 | n13331 ;
  assign n13333 = n7196 & n13224 ;
  assign n13334 = n13332 | n13333 ;
  assign n13335 = n13334 ^ x23 ^ 1'b0 ;
  assign n13336 = ( n12947 & ~n13071 ) | ( n12947 & n13335 ) | ( ~n13071 & n13335 ) ;
  assign n13337 = n13335 ^ n13071 ^ n12947 ;
  assign n13338 = n7485 & n10711 ;
  assign n13339 = ( n7486 & n10909 ) | ( n7486 & n13338 ) | ( n10909 & n13338 ) ;
  assign n13340 = n13338 | n13339 ;
  assign n13341 = ( n7493 & ~n10669 ) | ( n7493 & n13338 ) | ( ~n10669 & n13338 ) ;
  assign n13342 = n13340 | n13341 ;
  assign n13343 = n7487 & n13224 ;
  assign n13344 = n13342 | n13343 ;
  assign n13345 = n13344 ^ x17 ^ 1'b0 ;
  assign n13346 = n13345 ^ n13249 ^ n13096 ;
  assign n13347 = ( n13096 & n13249 ) | ( n13096 & n13345 ) | ( n13249 & n13345 ) ;
  assign n13348 = n7037 & n10909 ;
  assign n13349 = n13167 ^ x29 ^ 1'b0 ;
  assign n13350 = ( n7036 & n10711 ) | ( n7036 & n13348 ) | ( n10711 & n13348 ) ;
  assign n13351 = n13348 | n13350 ;
  assign n13352 = ( n7052 & ~n10669 ) | ( n7052 & n13348 ) | ( ~n10669 & n13348 ) ;
  assign n13353 = n13351 | n13352 ;
  assign n13354 = n7035 & n13224 ;
  assign n13355 = n13353 | n13354 ;
  assign n13356 = n13355 ^ x26 ^ 1'b0 ;
  assign n13357 = n13356 ^ n13349 ^ n12736 ;
  assign n13358 = ( ~n12736 & n13349 ) | ( ~n12736 & n13356 ) | ( n13349 & n13356 ) ;
  assign n13359 = n7669 & n10711 ;
  assign n13360 = ( n7674 & ~n10669 ) | ( n7674 & n13359 ) | ( ~n10669 & n13359 ) ;
  assign n13361 = n13359 | n13360 ;
  assign n13362 = ( n7667 & n10909 ) | ( n7667 & n13359 ) | ( n10909 & n13359 ) ;
  assign n13363 = n13361 | n13362 ;
  assign n13364 = ( n7666 & n13224 ) | ( n7666 & n13363 ) | ( n13224 & n13363 ) ;
  assign n13365 = n13363 | n13364 ;
  assign n13366 = n13365 ^ x14 ^ 1'b0 ;
  assign n13367 = ( ~n13084 & n13258 ) | ( ~n13084 & n13366 ) | ( n13258 & n13366 ) ;
  assign n13368 = n13366 ^ n13258 ^ n13084 ;
  assign n13369 = n7339 & n10711 ;
  assign n13370 = ( n7337 & n10909 ) | ( n7337 & n13369 ) | ( n10909 & n13369 ) ;
  assign n13371 = n13369 | n13370 ;
  assign n13372 = ( n7338 & ~n10669 ) | ( n7338 & n13369 ) | ( ~n10669 & n13369 ) ;
  assign n13373 = n13371 | n13372 ;
  assign n13374 = ( n7340 & n13224 ) | ( n7340 & n13373 ) | ( n13224 & n13373 ) ;
  assign n13375 = n13373 | n13374 ;
  assign n13376 = n13375 ^ x20 ^ 1'b0 ;
  assign n13377 = ( n12803 & n13238 ) | ( n12803 & n13376 ) | ( n13238 & n13376 ) ;
  assign n13378 = n13376 ^ n13238 ^ n12803 ;
  assign n13379 = n8029 & n10711 ;
  assign n13380 = ( n8037 & ~n10669 ) | ( n8037 & n13379 ) | ( ~n10669 & n13379 ) ;
  assign n13381 = n13379 | n13380 ;
  assign n13382 = ( n8033 & n10909 ) | ( n8033 & n13379 ) | ( n10909 & n13379 ) ;
  assign n13383 = n13381 | n13382 ;
  assign n13384 = ( n8034 & n13224 ) | ( n8034 & n13383 ) | ( n13224 & n13383 ) ;
  assign n13385 = n13383 | n13384 ;
  assign n13386 = n13385 ^ x5 ^ 1'b0 ;
  assign n13387 = n13386 ^ n13214 ^ n12994 ;
  assign n13388 = ( n12994 & n13214 ) | ( n12994 & n13386 ) | ( n13214 & n13386 ) ;
  assign n13389 = n7932 & n10711 ;
  assign n13390 = ( n7943 & ~n10669 ) | ( n7943 & n13389 ) | ( ~n10669 & n13389 ) ;
  assign n13391 = n13389 | n13390 ;
  assign n13392 = ( n7929 & n10909 ) | ( n7929 & n13389 ) | ( n10909 & n13389 ) ;
  assign n13393 = n13391 | n13392 ;
  assign n13394 = ( n7930 & n13224 ) | ( n7930 & n13393 ) | ( n13224 & n13393 ) ;
  assign n13395 = n13393 | n13394 ;
  assign n13396 = n13395 ^ x8 ^ 1'b0 ;
  assign n13397 = n13396 ^ n13188 ^ n13007 ;
  assign n13398 = ( n13007 & n13188 ) | ( n13007 & n13396 ) | ( n13188 & n13396 ) ;
  assign n13399 = n13297 ^ n13174 ^ n6717 ;
  assign n13400 = ( n6717 & n13174 ) | ( n6717 & ~n13297 ) | ( n13174 & ~n13297 ) ;
  assign n13401 = n7485 & n10909 ;
  assign n13402 = ( n7486 & ~n10930 ) | ( n7486 & n13401 ) | ( ~n10930 & n13401 ) ;
  assign n13403 = n13401 | n13402 ;
  assign n13404 = ( n7493 & n10711 ) | ( n7493 & n13401 ) | ( n10711 & n13401 ) ;
  assign n13405 = n13403 | n13404 ;
  assign n13406 = n7487 & ~n13265 ;
  assign n13407 = n13405 | n13406 ;
  assign n13408 = n13407 ^ x17 ^ 1'b0 ;
  assign n13409 = n13408 ^ n13347 ^ n13147 ;
  assign n13410 = ( n13147 & n13347 ) | ( n13147 & n13408 ) | ( n13347 & n13408 ) ;
  assign n13411 = n8029 & n10909 ;
  assign n13412 = ( n8037 & n10711 ) | ( n8037 & n13411 ) | ( n10711 & n13411 ) ;
  assign n13413 = n13411 | n13412 ;
  assign n13414 = ( n8033 & ~n10930 ) | ( n8033 & n13411 ) | ( ~n10930 & n13411 ) ;
  assign n13415 = n13413 | n13414 ;
  assign n13416 = n8034 & ~n13265 ;
  assign n13417 = n13415 | n13416 ;
  assign n13418 = n13417 ^ x5 ^ 1'b0 ;
  assign n13419 = n13418 ^ n13388 ^ n13033 ;
  assign n13420 = ( n13033 & n13388 ) | ( n13033 & n13418 ) | ( n13388 & n13418 ) ;
  assign n13421 = n6791 & n10711 ;
  assign n13422 = ( n6788 & n10909 ) | ( n6788 & n13421 ) | ( n10909 & n13421 ) ;
  assign n13423 = n13421 | n13422 ;
  assign n13424 = ( n6790 & ~n10669 ) | ( n6790 & n13421 ) | ( ~n10669 & n13421 ) ;
  assign n13425 = n13423 | n13424 ;
  assign n13426 = n6901 & n10711 ;
  assign n13427 = ( n6906 & ~n10669 ) | ( n6906 & n13426 ) | ( ~n10669 & n13426 ) ;
  assign n13428 = n13426 | n13427 ;
  assign n13429 = ( n6907 & n10909 ) | ( n6907 & n13426 ) | ( n10909 & n13426 ) ;
  assign n13430 = n13428 | n13429 ;
  assign n13431 = ( n6918 & n13224 ) | ( n6918 & n13430 ) | ( n13224 & n13430 ) ;
  assign n13432 = n6789 & ~n13224 ;
  assign n13433 = ( n6789 & n13425 ) | ( n6789 & ~n13432 ) | ( n13425 & ~n13432 ) ;
  assign n13434 = n7932 & n10909 ;
  assign n13435 = n13430 | n13431 ;
  assign n13436 = ( n7943 & n10711 ) | ( n7943 & n13434 ) | ( n10711 & n13434 ) ;
  assign n13437 = n13434 | n13436 ;
  assign n13438 = ( n7929 & ~n10930 ) | ( n7929 & n13434 ) | ( ~n10930 & n13434 ) ;
  assign n13439 = n13437 | n13438 ;
  assign n13440 = n7930 & ~n13265 ;
  assign n13441 = n13439 | n13440 ;
  assign n13442 = n13441 ^ x8 ^ 1'b0 ;
  assign n13443 = ( n13023 & n13398 ) | ( n13023 & n13442 ) | ( n13398 & n13442 ) ;
  assign n13444 = n13442 ^ n13398 ^ n13023 ;
  assign n13445 = n7829 & n10909 ;
  assign n13446 = ( n7833 & n10711 ) | ( n7833 & n13445 ) | ( n10711 & n13445 ) ;
  assign n13447 = n13445 | n13446 ;
  assign n13448 = ( n7834 & ~n10930 ) | ( n7834 & n13445 ) | ( ~n10930 & n13445 ) ;
  assign n13449 = n13447 | n13448 ;
  assign n13450 = n7838 & ~n13265 ;
  assign n13451 = n13449 | n13450 ;
  assign n13452 = n13451 ^ x11 ^ 1'b0 ;
  assign n13453 = ( ~n13117 & n13327 ) | ( ~n13117 & n13452 ) | ( n13327 & n13452 ) ;
  assign n13454 = n13452 ^ n13327 ^ n13117 ;
  assign n13455 = n6901 & ~n10930 ;
  assign n13456 = ( n6906 & n10909 ) | ( n6906 & n13455 ) | ( n10909 & n13455 ) ;
  assign n13457 = n13455 | n13456 ;
  assign n13458 = ( n6907 & n10926 ) | ( n6907 & n13455 ) | ( n10926 & n13455 ) ;
  assign n13459 = n13457 | n13458 ;
  assign n13460 = n6918 & ~n13306 ;
  assign n13461 = n13459 & ~n13460 ;
  assign n13462 = n13461 ^ n13460 ^ x29 ;
  assign n13463 = n13433 ^ n6717 ^ n6638 ;
  assign n13464 = ( n6638 & ~n6717 ) | ( n6638 & n13433 ) | ( ~n6717 & n13433 ) ;
  assign n13465 = n13435 ^ x29 ^ 1'b0 ;
  assign n13466 = ( n13176 & n13399 ) | ( n13176 & n13462 ) | ( n13399 & n13462 ) ;
  assign n13467 = n13462 ^ n13399 ^ n13176 ;
  assign n13468 = ( n13155 & ~n13164 ) | ( n13155 & n13465 ) | ( ~n13164 & n13465 ) ;
  assign n13469 = n13465 ^ n13164 ^ n13155 ;
  assign n13470 = n13466 ^ n13463 ^ n13400 ;
  assign n13471 = ( n13400 & n13463 ) | ( n13400 & ~n13466 ) | ( n13463 & ~n13466 ) ;
  assign n13472 = n6901 & n10909 ;
  assign n13473 = ( n6906 & n10711 ) | ( n6906 & n13472 ) | ( n10711 & n13472 ) ;
  assign n13474 = ( n6907 & ~n10930 ) | ( n6907 & n13472 ) | ( ~n10930 & n13472 ) ;
  assign n13475 = n13472 | n13473 ;
  assign n13476 = n6918 & ~n13265 ;
  assign n13477 = n13474 | n13475 ;
  assign n13478 = n13476 | n13477 ;
  assign n13479 = n13478 ^ x29 ^ 1'b0 ;
  assign n13480 = n7035 & ~n13265 ;
  assign n13481 = n13479 ^ n13468 ^ n13175 ;
  assign n13482 = n7037 & ~n10930 ;
  assign n13483 = ( ~n13175 & n13468 ) | ( ~n13175 & n13479 ) | ( n13468 & n13479 ) ;
  assign n13484 = ( n7036 & n10909 ) | ( n7036 & n13482 ) | ( n10909 & n13482 ) ;
  assign n13485 = n13482 | n13484 ;
  assign n13486 = ( n7052 & n10711 ) | ( n7052 & n13482 ) | ( n10711 & n13482 ) ;
  assign n13487 = n13485 | n13486 ;
  assign n13488 = n13480 | n13487 ;
  assign n13489 = n13488 ^ x26 ^ 1'b0 ;
  assign n13490 = ( ~n13138 & n13358 ) | ( ~n13138 & n13489 ) | ( n13358 & n13489 ) ;
  assign n13491 = n7339 & n10909 ;
  assign n13492 = ( n7337 & ~n10930 ) | ( n7337 & n13491 ) | ( ~n10930 & n13491 ) ;
  assign n13493 = n13491 | n13492 ;
  assign n13494 = ( n7338 & n10711 ) | ( n7338 & n13491 ) | ( n10711 & n13491 ) ;
  assign n13495 = n13493 | n13494 ;
  assign n13496 = n7340 & ~n13265 ;
  assign n13497 = n13495 | n13496 ;
  assign n13498 = n13497 ^ x20 ^ 1'b0 ;
  assign n13499 = n7340 & ~n13306 ;
  assign n13500 = n13489 ^ n13358 ^ n13138 ;
  assign n13501 = n7339 & ~n10930 ;
  assign n13502 = ( n12805 & ~n13058 ) | ( n12805 & n13498 ) | ( ~n13058 & n13498 ) ;
  assign n13503 = n13498 ^ n13058 ^ n12805 ;
  assign n13504 = ( n7337 & n10926 ) | ( n7337 & n13501 ) | ( n10926 & n13501 ) ;
  assign n13505 = ( n7338 & n10909 ) | ( n7338 & n13501 ) | ( n10909 & n13501 ) ;
  assign n13506 = n13501 | n13504 ;
  assign n13507 = n7669 & n10909 ;
  assign n13508 = n13505 | n13506 ;
  assign n13509 = ( n7674 & n10711 ) | ( n7674 & n13507 ) | ( n10711 & n13507 ) ;
  assign n13510 = n13507 | n13509 ;
  assign n13511 = ( n7667 & ~n10930 ) | ( n7667 & n13507 ) | ( ~n10930 & n13507 ) ;
  assign n13512 = n13499 | n13508 ;
  assign n13513 = n7188 & ~n10930 ;
  assign n13514 = n13510 | n13511 ;
  assign n13515 = n13512 ^ x20 ^ 1'b0 ;
  assign n13516 = ( n7190 & n10711 ) | ( n7190 & n13513 ) | ( n10711 & n13513 ) ;
  assign n13517 = n13513 | n13516 ;
  assign n13518 = ( n7192 & n10909 ) | ( n7192 & n13513 ) | ( n10909 & n13513 ) ;
  assign n13519 = n13517 | n13518 ;
  assign n13520 = n7666 & ~n13265 ;
  assign n13521 = n13514 & ~n13520 ;
  assign n13522 = n13521 ^ n13520 ^ x14 ;
  assign n13523 = n7665 ^ x14 ^ 1'b0 ;
  assign n13524 = n13523 ^ n6717 ^ n6641 ;
  assign n13525 = ( n6641 & ~n6717 ) | ( n6641 & n13523 ) | ( ~n6717 & n13523 ) ;
  assign n13526 = n6789 & ~n13265 ;
  assign n13527 = n7196 & ~n13265 ;
  assign n13528 = n13519 | n13527 ;
  assign n13529 = ( ~n13107 & n13367 ) | ( ~n13107 & n13522 ) | ( n13367 & n13522 ) ;
  assign n13530 = n13522 ^ n13367 ^ n13107 ;
  assign n13531 = ( n13059 & n13295 ) | ( n13059 & n13515 ) | ( n13295 & n13515 ) ;
  assign n13532 = n13515 ^ n13295 ^ n13059 ;
  assign n13533 = n6791 & n10909 ;
  assign n13534 = n13528 ^ x23 ^ 1'b0 ;
  assign n13535 = ( n6788 & ~n10930 ) | ( n6788 & n13533 ) | ( ~n10930 & n13533 ) ;
  assign n13536 = n13533 | n13535 ;
  assign n13537 = ( n6790 & n10711 ) | ( n6790 & n13533 ) | ( n10711 & n13533 ) ;
  assign n13538 = n13536 | n13537 ;
  assign n13539 = n13534 ^ n13336 ^ n13085 ;
  assign n13540 = ( ~n13085 & n13336 ) | ( ~n13085 & n13534 ) | ( n13336 & n13534 ) ;
  assign n13541 = n13526 | n13538 ;
  assign n13542 = ( n13464 & n13524 ) | ( n13464 & n13541 ) | ( n13524 & n13541 ) ;
  assign n13543 = n13541 ^ n13524 ^ n13464 ;
  assign n13544 = n7037 & n10926 ;
  assign n13545 = ( n7036 & ~n10930 ) | ( n7036 & n13544 ) | ( ~n10930 & n13544 ) ;
  assign n13546 = n13544 | n13545 ;
  assign n13547 = ( n7052 & n10909 ) | ( n7052 & n13544 ) | ( n10909 & n13544 ) ;
  assign n13548 = n13546 | n13547 ;
  assign n13549 = n7035 & ~n13306 ;
  assign n13550 = n13548 | n13549 ;
  assign n13551 = n13550 ^ x26 ^ 1'b0 ;
  assign n13552 = ( n13137 & ~n13283 ) | ( n13137 & n13551 ) | ( ~n13283 & n13551 ) ;
  assign n13553 = n13551 ^ n13283 ^ n13137 ;
  assign n13554 = n7485 & ~n10930 ;
  assign n13555 = ( n7486 & n10926 ) | ( n7486 & n13554 ) | ( n10926 & n13554 ) ;
  assign n13556 = n13554 | n13555 ;
  assign n13557 = ( n7493 & n10909 ) | ( n7493 & n13554 ) | ( n10909 & n13554 ) ;
  assign n13558 = n13556 | n13557 ;
  assign n13559 = n7487 & ~n13306 ;
  assign n13560 = n13558 | n13559 ;
  assign n13561 = n13560 ^ x17 ^ 1'b0 ;
  assign n13562 = n13561 ^ n13410 ^ n13239 ;
  assign n13563 = ( n13239 & n13410 ) | ( n13239 & n13561 ) | ( n13410 & n13561 ) ;
  assign n13564 = n7188 & n10926 ;
  assign n13565 = ( n7190 & n10909 ) | ( n7190 & n13564 ) | ( n10909 & n13564 ) ;
  assign n13566 = n13564 | n13565 ;
  assign n13567 = ( n7192 & ~n10930 ) | ( n7192 & n13564 ) | ( ~n10930 & n13564 ) ;
  assign n13568 = n13566 | n13567 ;
  assign n13569 = n7196 & ~n13306 ;
  assign n13570 = n13568 | n13569 ;
  assign n13571 = n13570 ^ x23 ^ 1'b0 ;
  assign n13572 = n13571 ^ n13216 ^ n13086 ;
  assign n13573 = ( n13086 & n13216 ) | ( n13086 & n13571 ) | ( n13216 & n13571 ) ;
  assign n13574 = n8029 & ~n10930 ;
  assign n13575 = ( n8037 & n10909 ) | ( n8037 & n13574 ) | ( n10909 & n13574 ) ;
  assign n13576 = n13574 | n13575 ;
  assign n13577 = ( n8033 & n10926 ) | ( n8033 & n13574 ) | ( n10926 & n13574 ) ;
  assign n13578 = n13576 | n13577 ;
  assign n13579 = n8034 & ~n13306 ;
  assign n13580 = n13578 | n13579 ;
  assign n13581 = n13580 ^ x5 ^ 1'b0 ;
  assign n13582 = ( n13187 & n13420 ) | ( n13187 & n13581 ) | ( n13420 & n13581 ) ;
  assign n13583 = n13581 ^ n13420 ^ n13187 ;
  assign n13584 = n7932 & ~n10930 ;
  assign n13585 = ( n7943 & n10909 ) | ( n7943 & n13584 ) | ( n10909 & n13584 ) ;
  assign n13586 = n13584 | n13585 ;
  assign n13587 = ( n7929 & n10926 ) | ( n7929 & n13584 ) | ( n10926 & n13584 ) ;
  assign n13588 = n13586 | n13587 ;
  assign n13589 = n7930 & ~n13306 ;
  assign n13590 = n13588 | n13589 ;
  assign n13591 = n13590 ^ x8 ^ 1'b0 ;
  assign n13592 = ( n13312 & n13443 ) | ( n13312 & n13591 ) | ( n13443 & n13591 ) ;
  assign n13593 = n13591 ^ n13443 ^ n13312 ;
  assign n13594 = n7669 & ~n10930 ;
  assign n13595 = ( n7674 & n10909 ) | ( n7674 & n13594 ) | ( n10909 & n13594 ) ;
  assign n13596 = n13594 | n13595 ;
  assign n13597 = ( n7667 & n10926 ) | ( n7667 & n13594 ) | ( n10926 & n13594 ) ;
  assign n13598 = n13596 | n13597 ;
  assign n13599 = n7666 & ~n13306 ;
  assign n13600 = n13598 & ~n13599 ;
  assign n13601 = n13600 ^ n13599 ^ x14 ;
  assign n13602 = n13601 ^ n13529 ^ n13248 ;
  assign n13603 = ( n13248 & n13529 ) | ( n13248 & n13601 ) | ( n13529 & n13601 ) ;
  assign n13604 = n6789 & ~n13306 ;
  assign n13605 = ( n6791 & ~n10930 ) | ( n6791 & n13604 ) | ( ~n10930 & n13604 ) ;
  assign n13606 = n13604 | n13605 ;
  assign n13607 = ( n6790 & n10909 ) | ( n6790 & n13604 ) | ( n10909 & n13604 ) ;
  assign n13608 = n13606 | n13607 ;
  assign n13609 = n7829 & ~n10930 ;
  assign n13610 = n7838 & ~n13306 ;
  assign n13611 = ( n7833 & n10909 ) | ( n7833 & n13609 ) | ( n10909 & n13609 ) ;
  assign n13612 = n13609 | n13611 ;
  assign n13613 = ( n10926 & ~n10930 ) | ( n10926 & n13298 ) | ( ~n10930 & n13298 ) ;
  assign n13614 = ( n7834 & n10926 ) | ( n7834 & n13609 ) | ( n10926 & n13609 ) ;
  assign n13615 = n13612 | n13614 ;
  assign n13616 = n13613 ^ n10938 ^ n10926 ;
  assign n13617 = n13610 | n13615 ;
  assign n13618 = n13617 ^ x11 ^ 1'b0 ;
  assign n13619 = ( n13260 & n13453 ) | ( n13260 & n13618 ) | ( n13453 & n13618 ) ;
  assign n13620 = n13618 ^ n13453 ^ n13260 ;
  assign n13621 = n8086 & ~n10930 ;
  assign n13622 = ( n8088 & n10926 ) | ( n8088 & n13621 ) | ( n10926 & n13621 ) ;
  assign n13623 = n13621 | n13622 ;
  assign n13624 = ( n8090 & ~n10938 ) | ( n8090 & n13621 ) | ( ~n10938 & n13621 ) ;
  assign n13625 = n13623 | n13624 ;
  assign n13626 = n8089 & ~n13616 ;
  assign n13627 = n13625 | n13626 ;
  assign n13628 = n13627 ^ x2 ^ 1'b0 ;
  assign n13629 = ( n13317 & n13387 ) | ( n13317 & n13628 ) | ( n13387 & n13628 ) ;
  assign n13630 = n7669 & n10926 ;
  assign n13631 = ( n7667 & ~n10938 ) | ( n7667 & n13630 ) | ( ~n10938 & n13630 ) ;
  assign n13632 = ( n7674 & ~n10930 ) | ( n7674 & n13630 ) | ( ~n10930 & n13630 ) ;
  assign n13633 = n13630 | n13632 ;
  assign n13634 = n13631 | n13633 ;
  assign n13635 = n7339 & n10926 ;
  assign n13636 = ( n7337 & ~n10938 ) | ( n7337 & n13635 ) | ( ~n10938 & n13635 ) ;
  assign n13637 = n13635 | n13636 ;
  assign n13638 = ( n7338 & ~n10930 ) | ( n7338 & n13635 ) | ( ~n10930 & n13635 ) ;
  assign n13639 = n13637 | n13638 ;
  assign n13640 = n7340 & ~n13616 ;
  assign n13641 = n13639 | n13640 ;
  assign n13642 = n13641 ^ x20 ^ 1'b0 ;
  assign n13643 = ( n13294 & ~n13337 ) | ( n13294 & n13642 ) | ( ~n13337 & n13642 ) ;
  assign n13644 = n7493 ^ n7492 ^ x17 ;
  assign n13645 = n13642 ^ n13337 ^ n13294 ;
  assign n13646 = n7037 & ~n10938 ;
  assign n13647 = ( n7036 & n10926 ) | ( n7036 & n13646 ) | ( n10926 & n13646 ) ;
  assign n13648 = n13646 | n13647 ;
  assign n13649 = ( n7052 & ~n10930 ) | ( n7052 & n13646 ) | ( ~n10930 & n13646 ) ;
  assign n13650 = n13648 | n13649 ;
  assign n13651 = n7666 & ~n13616 ;
  assign n13652 = n13634 & ~n13651 ;
  assign n13653 = n13652 ^ n13651 ^ x14 ;
  assign n13654 = n7035 & ~n13616 ;
  assign n13655 = n13650 | n13654 ;
  assign n13656 = ( n13346 & n13603 ) | ( n13346 & n13653 ) | ( n13603 & n13653 ) ;
  assign n13657 = n13653 ^ n13603 ^ n13346 ;
  assign n13658 = n13655 ^ x26 ^ 1'b0 ;
  assign n13659 = ( n13284 & ~n13469 ) | ( n13284 & n13658 ) | ( ~n13469 & n13658 ) ;
  assign n13660 = n13658 ^ n13469 ^ n13284 ;
  assign n13661 = n7669 & ~n10938 ;
  assign n13662 = ( n7674 & n10926 ) | ( n7674 & n13661 ) | ( n10926 & n13661 ) ;
  assign n13663 = n13661 | n13662 ;
  assign n13664 = ( n7667 & n10964 ) | ( n7667 & n13661 ) | ( n10964 & n13661 ) ;
  assign n13665 = n13663 | n13664 ;
  assign n13666 = ( n10926 & ~n10938 ) | ( n10926 & n13613 ) | ( ~n10938 & n13613 ) ;
  assign n13667 = n8029 & n10926 ;
  assign n13668 = ( n8037 & ~n10930 ) | ( n8037 & n13667 ) | ( ~n10930 & n13667 ) ;
  assign n13669 = n13667 | n13668 ;
  assign n13670 = ( n8033 & ~n10938 ) | ( n8033 & n13667 ) | ( ~n10938 & n13667 ) ;
  assign n13671 = n13669 | n13670 ;
  assign n13672 = n8034 & ~n13616 ;
  assign n13673 = n13671 | n13672 ;
  assign n13674 = n13673 ^ x5 ^ 1'b0 ;
  assign n13675 = n13674 ^ n13582 ^ n13397 ;
  assign n13676 = ( n13397 & n13582 ) | ( n13397 & n13674 ) | ( n13582 & n13674 ) ;
  assign n13677 = n13666 ^ n10964 ^ n10938 ;
  assign n13678 = n7666 & ~n13677 ;
  assign n13679 = n13665 & ~n13678 ;
  assign n13680 = n13679 ^ n13678 ^ x14 ;
  assign n13681 = n13680 ^ n13656 ^ n13409 ;
  assign n13682 = ( n13409 & n13656 ) | ( n13409 & n13680 ) | ( n13656 & n13680 ) ;
  assign n13683 = n6901 & ~n10938 ;
  assign n13684 = ( n6906 & n10926 ) | ( n6906 & n13683 ) | ( n10926 & n13683 ) ;
  assign n13685 = n13683 | n13684 ;
  assign n13686 = ( n6907 & n10964 ) | ( n6907 & n13683 ) | ( n10964 & n13683 ) ;
  assign n13687 = n13685 | n13686 ;
  assign n13688 = n6918 & ~n13677 ;
  assign n13689 = n13687 | n13688 ;
  assign n13690 = n13689 ^ x29 ^ 1'b0 ;
  assign n13691 = n13690 ^ n13543 ^ n13471 ;
  assign n13692 = ( ~n13471 & n13543 ) | ( ~n13471 & n13690 ) | ( n13543 & n13690 ) ;
  assign n13693 = n8086 & n10926 ;
  assign n13694 = ( n8088 & ~n10938 ) | ( n8088 & n13693 ) | ( ~n10938 & n13693 ) ;
  assign n13695 = n13693 | n13694 ;
  assign n13696 = ( n8090 & n10964 ) | ( n8090 & n13693 ) | ( n10964 & n13693 ) ;
  assign n13697 = n13695 | n13696 ;
  assign n13698 = n8089 & ~n13677 ;
  assign n13699 = n13697 & ~n13698 ;
  assign n13700 = n13699 ^ n13698 ^ x2 ;
  assign n13701 = n7035 & ~n13677 ;
  assign n13702 = ( n13419 & n13629 ) | ( n13419 & n13700 ) | ( n13629 & n13700 ) ;
  assign n13703 = n7037 & n10964 ;
  assign n13704 = ( n7036 & ~n10938 ) | ( n7036 & n13703 ) | ( ~n10938 & n13703 ) ;
  assign n13705 = n13703 | n13704 ;
  assign n13706 = ( n7052 & n10926 ) | ( n7052 & n13703 ) | ( n10926 & n13703 ) ;
  assign n13707 = n13705 | n13706 ;
  assign n13708 = n13701 | n13707 ;
  assign n13709 = n13708 ^ x26 ^ 1'b0 ;
  assign n13710 = n13709 ^ n13659 ^ n13481 ;
  assign n13711 = ( ~n13481 & n13659 ) | ( ~n13481 & n13709 ) | ( n13659 & n13709 ) ;
  assign n13712 = n6791 & ~n10938 ;
  assign n13713 = ( n6788 & n10964 ) | ( n6788 & n13712 ) | ( n10964 & n13712 ) ;
  assign n13714 = n13712 | n13713 ;
  assign n13715 = ( n6790 & n10926 ) | ( n6790 & n13712 ) | ( n10926 & n13712 ) ;
  assign n13716 = n13714 | n13715 ;
  assign n13717 = n6788 & ~n10926 ;
  assign n13718 = ( n6788 & n13608 ) | ( n6788 & ~n13717 ) | ( n13608 & ~n13717 ) ;
  assign n13719 = n13718 ^ n13525 ^ n6660 ;
  assign n13720 = ( n6660 & n13525 ) | ( n6660 & ~n13718 ) | ( n13525 & ~n13718 ) ;
  assign n13721 = ( n6660 & n6713 ) | ( n6660 & ~n13720 ) | ( n6713 & ~n13720 ) ;
  assign n13722 = n13720 ^ n6713 ^ n6660 ;
  assign n13723 = n13644 ^ n6778 ^ n6713 ;
  assign n13724 = ( n6713 & ~n6778 ) | ( n6713 & n13644 ) | ( ~n6778 & n13644 ) ;
  assign n13725 = n6789 & ~n13677 ;
  assign n13726 = n13716 | n13725 ;
  assign n13727 = n13726 ^ n13723 ^ n13721 ;
  assign n13728 = ( n13721 & n13723 ) | ( n13721 & n13726 ) | ( n13723 & n13726 ) ;
  assign n13729 = n7485 & ~n10938 ;
  assign n13730 = ( n7486 & n10964 ) | ( n7486 & n13729 ) | ( n10964 & n13729 ) ;
  assign n13731 = n13729 | n13730 ;
  assign n13732 = ( n7493 & n10926 ) | ( n7493 & n13729 ) | ( n10926 & n13729 ) ;
  assign n13733 = n13731 | n13732 ;
  assign n13734 = n7487 & ~n13677 ;
  assign n13735 = n13733 | n13734 ;
  assign n13736 = n13735 ^ x17 ^ 1'b0 ;
  assign n13737 = ( n13377 & ~n13503 ) | ( n13377 & n13736 ) | ( ~n13503 & n13736 ) ;
  assign n13738 = n13736 ^ n13503 ^ n13377 ;
  assign n13739 = n7188 & ~n10938 ;
  assign n13740 = ( n7190 & ~n10930 ) | ( n7190 & n13739 ) | ( ~n10930 & n13739 ) ;
  assign n13741 = n13739 | n13740 ;
  assign n13742 = ( n7192 & n10926 ) | ( n7192 & n13739 ) | ( n10926 & n13739 ) ;
  assign n13743 = n13741 | n13742 ;
  assign n13744 = n7196 & ~n13616 ;
  assign n13745 = n13743 | n13744 ;
  assign n13746 = n13745 ^ x23 ^ 1'b0 ;
  assign n13747 = ( n13218 & ~n13357 ) | ( n13218 & n13746 ) | ( ~n13357 & n13746 ) ;
  assign n13748 = n13746 ^ n13357 ^ n13218 ;
  assign n13749 = n7188 & n10964 ;
  assign n13750 = ( n7190 & n10926 ) | ( n7190 & n13749 ) | ( n10926 & n13749 ) ;
  assign n13751 = n13749 | n13750 ;
  assign n13752 = ( n7192 & ~n10938 ) | ( n7192 & n13749 ) | ( ~n10938 & n13749 ) ;
  assign n13753 = n13751 | n13752 ;
  assign n13754 = n7196 & ~n13677 ;
  assign n13755 = n13753 | n13754 ;
  assign n13756 = n13755 ^ x23 ^ 1'b0 ;
  assign n13757 = n13756 ^ n13747 ^ n13500 ;
  assign n13758 = ( ~n13500 & n13747 ) | ( ~n13500 & n13756 ) | ( n13747 & n13756 ) ;
  assign n13759 = n7485 & n10926 ;
  assign n13760 = ( n7486 & ~n10938 ) | ( n7486 & n13759 ) | ( ~n10938 & n13759 ) ;
  assign n13761 = n13759 | n13760 ;
  assign n13762 = ( n7493 & ~n10930 ) | ( n7493 & n13759 ) | ( ~n10930 & n13759 ) ;
  assign n13763 = n13761 | n13762 ;
  assign n13764 = n7487 & ~n13616 ;
  assign n13765 = n13763 | n13764 ;
  assign n13766 = n13765 ^ x17 ^ 1'b0 ;
  assign n13767 = n13766 ^ n13563 ^ n13378 ;
  assign n13768 = ( n13378 & n13563 ) | ( n13378 & n13766 ) | ( n13563 & n13766 ) ;
  assign n13769 = n7829 & n10926 ;
  assign n13770 = ( n7833 & ~n10930 ) | ( n7833 & n13769 ) | ( ~n10930 & n13769 ) ;
  assign n13771 = n13769 | n13770 ;
  assign n13772 = ( n7834 & ~n10938 ) | ( n7834 & n13769 ) | ( ~n10938 & n13769 ) ;
  assign n13773 = n13771 | n13772 ;
  assign n13774 = n7838 & ~n13616 ;
  assign n13775 = n13773 | n13774 ;
  assign n13776 = n13775 ^ x11 ^ 1'b0 ;
  assign n13777 = n13776 ^ n13619 ^ n13368 ;
  assign n13778 = ( ~n13368 & n13619 ) | ( ~n13368 & n13776 ) | ( n13619 & n13776 ) ;
  assign n13779 = n7339 & ~n10938 ;
  assign n13780 = ( n7337 & n10964 ) | ( n7337 & n13779 ) | ( n10964 & n13779 ) ;
  assign n13781 = n13779 | n13780 ;
  assign n13782 = ( n7338 & n10926 ) | ( n7338 & n13779 ) | ( n10926 & n13779 ) ;
  assign n13783 = n13781 | n13782 ;
  assign n13784 = n7340 & ~n13677 ;
  assign n13785 = n13783 | n13784 ;
  assign n13786 = n7930 & ~n13616 ;
  assign n13787 = n13785 ^ x20 ^ 1'b0 ;
  assign n13788 = ( ~n13539 & n13643 ) | ( ~n13539 & n13787 ) | ( n13643 & n13787 ) ;
  assign n13789 = n13787 ^ n13643 ^ n13539 ;
  assign n13790 = n7932 & n10926 ;
  assign n13791 = ( n7943 & ~n10930 ) | ( n7943 & n13790 ) | ( ~n10930 & n13790 ) ;
  assign n13792 = n13790 | n13791 ;
  assign n13793 = ( n7929 & ~n10938 ) | ( n7929 & n13790 ) | ( ~n10938 & n13790 ) ;
  assign n13794 = n13792 | n13793 ;
  assign n13795 = ~n13786 & n13794 ;
  assign n13796 = n8029 & ~n10938 ;
  assign n13797 = n13795 ^ n13786 ^ x8 ;
  assign n13798 = ( n8037 & n10926 ) | ( n8037 & n13796 ) | ( n10926 & n13796 ) ;
  assign n13799 = n13796 | n13798 ;
  assign n13800 = ( n8033 & n10964 ) | ( n8033 & n13796 ) | ( n10964 & n13796 ) ;
  assign n13801 = n13799 | n13800 ;
  assign n13802 = n13797 ^ n13592 ^ n13326 ;
  assign n13803 = ( ~n13326 & n13592 ) | ( ~n13326 & n13797 ) | ( n13592 & n13797 ) ;
  assign n13804 = n7932 & ~n10938 ;
  assign n13805 = ( n7943 & n10926 ) | ( n7943 & n13804 ) | ( n10926 & n13804 ) ;
  assign n13806 = n13804 | n13805 ;
  assign n13807 = ( n7929 & n10964 ) | ( n7929 & n13804 ) | ( n10964 & n13804 ) ;
  assign n13808 = n13806 | n13807 ;
  assign n13809 = n8034 & ~n13677 ;
  assign n13810 = n13801 & ~n13809 ;
  assign n13811 = n13810 ^ n13809 ^ x5 ;
  assign n13812 = n7838 & ~n13677 ;
  assign n13813 = n7930 & ~n13677 ;
  assign n13814 = n13808 & ~n13813 ;
  assign n13815 = n13814 ^ n13813 ^ x8 ;
  assign n13816 = n13811 ^ n13676 ^ n13444 ;
  assign n13817 = ( n13444 & n13676 ) | ( n13444 & n13811 ) | ( n13676 & n13811 ) ;
  assign n13818 = ( ~n13454 & n13803 ) | ( ~n13454 & n13815 ) | ( n13803 & n13815 ) ;
  assign n13819 = n13815 ^ n13803 ^ n13454 ;
  assign n13820 = n6791 & n10926 ;
  assign n13821 = n7829 & ~n10938 ;
  assign n13822 = ( n7833 & n10926 ) | ( n7833 & n13821 ) | ( n10926 & n13821 ) ;
  assign n13823 = n13821 | n13822 ;
  assign n13824 = ( n7834 & n10964 ) | ( n7834 & n13821 ) | ( n10964 & n13821 ) ;
  assign n13825 = n13823 | n13824 ;
  assign n13826 = n6918 & ~n13616 ;
  assign n13827 = n6789 & ~n13616 ;
  assign n13828 = n13812 | n13825 ;
  assign n13829 = ( n6788 & ~n10938 ) | ( n6788 & n13820 ) | ( ~n10938 & n13820 ) ;
  assign n13830 = n13820 | n13829 ;
  assign n13831 = ( n6790 & ~n10930 ) | ( n6790 & n13820 ) | ( ~n10930 & n13820 ) ;
  assign n13832 = n13828 ^ x11 ^ 1'b0 ;
  assign n13833 = n13830 | n13831 ;
  assign n13834 = n6901 & n10926 ;
  assign n13835 = ( n6907 & ~n10938 ) | ( n6907 & n13834 ) | ( ~n10938 & n13834 ) ;
  assign n13836 = ( n6906 & ~n10930 ) | ( n6906 & n13834 ) | ( ~n10930 & n13834 ) ;
  assign n13837 = n13834 | n13836 ;
  assign n13838 = n13832 ^ n13778 ^ n13530 ;
  assign n13839 = ( ~n13530 & n13778 ) | ( ~n13530 & n13832 ) | ( n13778 & n13832 ) ;
  assign n13840 = n13827 | n13833 ;
  assign n13841 = n13835 | n13837 ;
  assign n13842 = n13826 | n13841 ;
  assign n13843 = n8086 & ~n10938 ;
  assign n13844 = ( n8090 & n10944 ) | ( n8090 & n13843 ) | ( n10944 & n13843 ) ;
  assign n13845 = ( n8088 & n10964 ) | ( n8088 & n13843 ) | ( n10964 & n13843 ) ;
  assign n13846 = n13843 | n13845 ;
  assign n13847 = n13844 | n13846 ;
  assign n13848 = ( ~n10938 & n10964 ) | ( ~n10938 & n13666 ) | ( n10964 & n13666 ) ;
  assign n13849 = n13848 ^ n10964 ^ n10944 ;
  assign n13850 = ( n8089 & n13847 ) | ( n8089 & n13849 ) | ( n13847 & n13849 ) ;
  assign n13851 = n13847 | n13850 ;
  assign n13852 = n7339 & n10964 ;
  assign n13853 = n13851 ^ x2 ^ 1'b0 ;
  assign n13854 = ( n13583 & n13702 ) | ( n13583 & n13853 ) | ( n13702 & n13853 ) ;
  assign n13855 = ( n7337 & n10944 ) | ( n7337 & n13852 ) | ( n10944 & n13852 ) ;
  assign n13856 = n13852 | n13855 ;
  assign n13857 = n7340 & n13849 ;
  assign n13858 = ( n7338 & ~n10938 ) | ( n7338 & n13852 ) | ( ~n10938 & n13852 ) ;
  assign n13859 = n13856 | n13858 ;
  assign n13860 = n13857 | n13859 ;
  assign n13861 = n13860 ^ x20 ^ 1'b0 ;
  assign n13862 = n13861 ^ n13572 ^ n13540 ;
  assign n13863 = n7188 & n10944 ;
  assign n13864 = ( n13540 & n13572 ) | ( n13540 & n13861 ) | ( n13572 & n13861 ) ;
  assign n13865 = ( n7190 & ~n10938 ) | ( n7190 & n13863 ) | ( ~n10938 & n13863 ) ;
  assign n13866 = n13863 | n13865 ;
  assign n13867 = n7487 & n13849 ;
  assign n13868 = ( n7192 & n10964 ) | ( n7192 & n13863 ) | ( n10964 & n13863 ) ;
  assign n13869 = n13866 | n13868 ;
  assign n13870 = n7196 & n13849 ;
  assign n13871 = n13869 | n13870 ;
  assign n13872 = n13871 ^ x23 ^ 1'b0 ;
  assign n13873 = n13872 ^ n13553 ^ n13490 ;
  assign n13874 = ( n13490 & ~n13553 ) | ( n13490 & n13872 ) | ( ~n13553 & n13872 ) ;
  assign n13875 = n7485 & n10964 ;
  assign n13876 = ( n7486 & n10944 ) | ( n7486 & n13875 ) | ( n10944 & n13875 ) ;
  assign n13877 = n13875 | n13876 ;
  assign n13878 = ( n7493 & ~n10938 ) | ( n7493 & n13875 ) | ( ~n10938 & n13875 ) ;
  assign n13879 = n13877 | n13878 ;
  assign n13880 = n13867 | n13879 ;
  assign n13881 = n7829 & n10964 ;
  assign n13882 = ( n7833 & ~n10938 ) | ( n7833 & n13881 ) | ( ~n10938 & n13881 ) ;
  assign n13883 = n13881 | n13882 ;
  assign n13884 = ( n7834 & n10944 ) | ( n7834 & n13881 ) | ( n10944 & n13881 ) ;
  assign n13885 = n13880 ^ x17 ^ 1'b0 ;
  assign n13886 = n13883 | n13884 ;
  assign n13887 = ( n13502 & n13532 ) | ( n13502 & n13885 ) | ( n13532 & n13885 ) ;
  assign n13888 = n13885 ^ n13532 ^ n13502 ;
  assign n13889 = n7838 & n13849 ;
  assign n13890 = n13886 | n13889 ;
  assign n13891 = n13890 ^ x11 ^ 1'b0 ;
  assign n13892 = ( n13602 & n13839 ) | ( n13602 & n13891 ) | ( n13839 & n13891 ) ;
  assign n13893 = n13891 ^ n13839 ^ n13602 ;
  assign n13894 = n8029 & n10964 ;
  assign n13895 = ( n8037 & ~n10938 ) | ( n8037 & n13894 ) | ( ~n10938 & n13894 ) ;
  assign n13896 = n13894 | n13895 ;
  assign n13897 = ( n8033 & n10944 ) | ( n8033 & n13894 ) | ( n10944 & n13894 ) ;
  assign n13898 = n13896 | n13897 ;
  assign n13899 = ( n8034 & n13849 ) | ( n8034 & n13898 ) | ( n13849 & n13898 ) ;
  assign n13900 = n13898 | n13899 ;
  assign n13901 = n13900 ^ x5 ^ 1'b0 ;
  assign n13902 = ( n13593 & n13817 ) | ( n13593 & n13901 ) | ( n13817 & n13901 ) ;
  assign n13903 = n13901 ^ n13817 ^ n13593 ;
  assign n13904 = n7037 & n10944 ;
  assign n13905 = ( n7036 & n10964 ) | ( n7036 & n13904 ) | ( n10964 & n13904 ) ;
  assign n13906 = n13904 | n13905 ;
  assign n13907 = ( n7052 & ~n10938 ) | ( n7052 & n13904 ) | ( ~n10938 & n13904 ) ;
  assign n13908 = n13906 | n13907 ;
  assign n13909 = n7035 & n13849 ;
  assign n13910 = n13908 | n13909 ;
  assign n13911 = n13910 ^ x26 ^ 1'b0 ;
  assign n13912 = n13911 ^ n13483 ^ n13467 ;
  assign n13913 = ( n13467 & n13483 ) | ( n13467 & n13911 ) | ( n13483 & n13911 ) ;
  assign n13914 = n7932 & n10964 ;
  assign n13915 = ( n7943 & ~n10938 ) | ( n7943 & n13914 ) | ( ~n10938 & n13914 ) ;
  assign n13916 = n13914 | n13915 ;
  assign n13917 = ( n7929 & n10944 ) | ( n7929 & n13914 ) | ( n10944 & n13914 ) ;
  assign n13918 = n13916 | n13917 ;
  assign n13919 = ( n7930 & n13849 ) | ( n7930 & n13918 ) | ( n13849 & n13918 ) ;
  assign n13920 = n13918 | n13919 ;
  assign n13921 = n13920 ^ x8 ^ 1'b0 ;
  assign n13922 = n13921 ^ n13818 ^ n13620 ;
  assign n13923 = ( n13620 & n13818 ) | ( n13620 & n13921 ) | ( n13818 & n13921 ) ;
  assign n13924 = n6901 & n10964 ;
  assign n13925 = ( n6906 & ~n10938 ) | ( n6906 & n13924 ) | ( ~n10938 & n13924 ) ;
  assign n13926 = n13924 | n13925 ;
  assign n13927 = ( n6907 & n10944 ) | ( n6907 & n13924 ) | ( n10944 & n13924 ) ;
  assign n13928 = n13926 | n13927 ;
  assign n13929 = ( n6918 & n13849 ) | ( n6918 & n13928 ) | ( n13849 & n13928 ) ;
  assign n13930 = n13928 | n13929 ;
  assign n13931 = n13930 ^ x29 ^ 1'b0 ;
  assign n13932 = n13931 ^ n13719 ^ n13542 ;
  assign n13933 = ( n13542 & n13719 ) | ( n13542 & n13931 ) | ( n13719 & n13931 ) ;
  assign n13934 = n7669 & n10964 ;
  assign n13935 = ( n7674 & ~n10938 ) | ( n7674 & n13934 ) | ( ~n10938 & n13934 ) ;
  assign n13936 = n13934 | n13935 ;
  assign n13937 = ( n7667 & n10944 ) | ( n7667 & n13934 ) | ( n10944 & n13934 ) ;
  assign n13938 = n13936 | n13937 ;
  assign n13939 = ( n7666 & n13849 ) | ( n7666 & n13938 ) | ( n13849 & n13938 ) ;
  assign n13940 = n6789 & n13849 ;
  assign n13941 = n13938 | n13939 ;
  assign n13942 = ( n6791 & n10964 ) | ( n6791 & n13940 ) | ( n10964 & n13940 ) ;
  assign n13943 = n13940 | n13942 ;
  assign n13944 = ( n6790 & ~n10938 ) | ( n6790 & n13940 ) | ( ~n10938 & n13940 ) ;
  assign n13945 = n13943 | n13944 ;
  assign n13946 = n13941 ^ x14 ^ 1'b0 ;
  assign n13947 = n13946 ^ n13682 ^ n13562 ;
  assign n13948 = ( n13562 & n13682 ) | ( n13562 & n13946 ) | ( n13682 & n13946 ) ;
  assign n13949 = n8086 & n10964 ;
  assign n13950 = ( n8088 & n10944 ) | ( n8088 & n13949 ) | ( n10944 & n13949 ) ;
  assign n13951 = ( n8090 & n10952 ) | ( n8090 & n13949 ) | ( n10952 & n13949 ) ;
  assign n13952 = n13949 | n13950 ;
  assign n13953 = ( n10944 & n10964 ) | ( n10944 & n13848 ) | ( n10964 & n13848 ) ;
  assign n13954 = n13953 ^ n10952 ^ n10944 ;
  assign n13955 = n13951 | n13952 ;
  assign n13956 = ( n8089 & n13954 ) | ( n8089 & n13955 ) | ( n13954 & n13955 ) ;
  assign n13957 = n13955 | n13956 ;
  assign n13958 = n13957 ^ x2 ^ 1'b0 ;
  assign n13959 = n6901 & n10944 ;
  assign n13960 = ( n13675 & n13854 ) | ( n13675 & n13958 ) | ( n13854 & n13958 ) ;
  assign n13961 = n7669 & n10944 ;
  assign n13962 = ( n7674 & n10964 ) | ( n7674 & n13961 ) | ( n10964 & n13961 ) ;
  assign n13963 = n13961 | n13962 ;
  assign n13964 = ( n7667 & n10952 ) | ( n7667 & n13961 ) | ( n10952 & n13961 ) ;
  assign n13965 = n13963 | n13964 ;
  assign n13966 = ( n7666 & n13954 ) | ( n7666 & n13965 ) | ( n13954 & n13965 ) ;
  assign n13967 = n13965 | n13966 ;
  assign n13968 = ( n6906 & n10964 ) | ( n6906 & n13959 ) | ( n10964 & n13959 ) ;
  assign n13969 = n13967 ^ x14 ^ 1'b0 ;
  assign n13970 = n13959 | n13968 ;
  assign n13971 = ( n6907 & n10952 ) | ( n6907 & n13959 ) | ( n10952 & n13959 ) ;
  assign n13972 = n13970 | n13971 ;
  assign n13973 = n13969 ^ n13948 ^ n13767 ;
  assign n13974 = ( n13767 & n13948 ) | ( n13767 & n13969 ) | ( n13948 & n13969 ) ;
  assign n13975 = n8029 & n10944 ;
  assign n13976 = ( n8037 & n10964 ) | ( n8037 & n13975 ) | ( n10964 & n13975 ) ;
  assign n13977 = n13975 | n13976 ;
  assign n13978 = ( n8033 & n10952 ) | ( n8033 & n13975 ) | ( n10952 & n13975 ) ;
  assign n13979 = n13977 | n13978 ;
  assign n13980 = n8034 & n13954 ;
  assign n13981 = n13979 | n13980 ;
  assign n13982 = ( n6918 & n13954 ) | ( n6918 & n13972 ) | ( n13954 & n13972 ) ;
  assign n13983 = n13972 | n13982 ;
  assign n13984 = n13981 ^ x5 ^ 1'b0 ;
  assign n13985 = n13983 ^ x29 ^ 1'b0 ;
  assign n13986 = ( ~n13722 & n13840 ) | ( ~n13722 & n13985 ) | ( n13840 & n13985 ) ;
  assign n13987 = n13985 ^ n13840 ^ n13722 ;
  assign n13988 = n7829 & n10944 ;
  assign n13989 = n13984 ^ n13902 ^ n13802 ;
  assign n13990 = ( ~n13802 & n13902 ) | ( ~n13802 & n13984 ) | ( n13902 & n13984 ) ;
  assign n13991 = ( n7833 & n10964 ) | ( n7833 & n13988 ) | ( n10964 & n13988 ) ;
  assign n13992 = n13988 | n13991 ;
  assign n13993 = ( n7834 & n10952 ) | ( n7834 & n13988 ) | ( n10952 & n13988 ) ;
  assign n13994 = n7838 & n13954 ;
  assign n13995 = n13992 | n13993 ;
  assign n13996 = n13994 | n13995 ;
  assign n13997 = n13996 ^ x11 ^ 1'b0 ;
  assign n13998 = n13997 ^ n13892 ^ n13657 ;
  assign n13999 = ( n13657 & n13892 ) | ( n13657 & n13997 ) | ( n13892 & n13997 ) ;
  assign n14000 = n7037 & n10952 ;
  assign n14001 = ( n7036 & n10944 ) | ( n7036 & n14000 ) | ( n10944 & n14000 ) ;
  assign n14002 = n14000 | n14001 ;
  assign n14003 = n13842 ^ x29 ^ 1'b0 ;
  assign n14004 = ( n7052 & n10964 ) | ( n7052 & n14000 ) | ( n10964 & n14000 ) ;
  assign n14005 = n14002 | n14004 ;
  assign n14006 = n7035 & n13954 ;
  assign n14007 = n14005 | n14006 ;
  assign n14008 = n14007 ^ x26 ^ 1'b0 ;
  assign n14009 = n14008 ^ n14003 ^ n13470 ;
  assign n14010 = ( n13470 & n14003 ) | ( n13470 & n14008 ) | ( n14003 & n14008 ) ;
  assign n14011 = n7485 & n10944 ;
  assign n14012 = ( n7486 & n10952 ) | ( n7486 & n14011 ) | ( n10952 & n14011 ) ;
  assign n14013 = n14011 | n14012 ;
  assign n14014 = ( n7493 & n10964 ) | ( n7493 & n14011 ) | ( n10964 & n14011 ) ;
  assign n14015 = n14013 | n14014 ;
  assign n14016 = n7487 & n13954 ;
  assign n14017 = n14015 | n14016 ;
  assign n14018 = n14017 ^ x17 ^ 1'b0 ;
  assign n14019 = ( n13531 & ~n13645 ) | ( n13531 & n14018 ) | ( ~n13645 & n14018 ) ;
  assign n14020 = n14018 ^ n13645 ^ n13531 ;
  assign n14021 = n7188 & n10952 ;
  assign n14022 = ( n7190 & n10964 ) | ( n7190 & n14021 ) | ( n10964 & n14021 ) ;
  assign n14023 = n14021 | n14022 ;
  assign n14024 = ( n7192 & n10944 ) | ( n7192 & n14021 ) | ( n10944 & n14021 ) ;
  assign n14025 = n14023 | n14024 ;
  assign n14026 = n7196 & n13954 ;
  assign n14027 = n14025 | n14026 ;
  assign n14028 = n14027 ^ x23 ^ 1'b0 ;
  assign n14029 = ( n13552 & ~n13660 ) | ( n13552 & n14028 ) | ( ~n13660 & n14028 ) ;
  assign n14030 = n14028 ^ n13660 ^ n13552 ;
  assign n14031 = n7339 & n10944 ;
  assign n14032 = ( n7337 & n10952 ) | ( n7337 & n14031 ) | ( n10952 & n14031 ) ;
  assign n14033 = n14031 | n14032 ;
  assign n14034 = ( n7338 & n10964 ) | ( n7338 & n14031 ) | ( n10964 & n14031 ) ;
  assign n14035 = n14033 | n14034 ;
  assign n14036 = n7340 & n13954 ;
  assign n14037 = n14035 | n14036 ;
  assign n14038 = n14037 ^ x20 ^ 1'b0 ;
  assign n14039 = n14038 ^ n13748 ^ n13573 ;
  assign n14040 = ( n13573 & ~n13748 ) | ( n13573 & n14038 ) | ( ~n13748 & n14038 ) ;
  assign n14041 = n6791 & n10944 ;
  assign n14042 = ( n6788 & n10952 ) | ( n6788 & n14041 ) | ( n10952 & n14041 ) ;
  assign n14043 = n14041 | n14042 ;
  assign n14044 = ( n6790 & n10964 ) | ( n6790 & n14041 ) | ( n10964 & n14041 ) ;
  assign n14045 = n14043 | n14044 ;
  assign n14046 = n7932 & n10944 ;
  assign n14047 = ( n7943 & n10964 ) | ( n7943 & n14046 ) | ( n10964 & n14046 ) ;
  assign n14048 = n14046 | n14047 ;
  assign n14049 = ( n7929 & n10952 ) | ( n7929 & n14046 ) | ( n10952 & n14046 ) ;
  assign n14050 = n14048 | n14049 ;
  assign n14051 = ( n7930 & n13954 ) | ( n7930 & n14050 ) | ( n13954 & n14050 ) ;
  assign n14052 = n14050 | n14051 ;
  assign n14053 = n14052 ^ x8 ^ 1'b0 ;
  assign n14054 = n14053 ^ n13923 ^ n13777 ;
  assign n14055 = ( ~n13777 & n13923 ) | ( ~n13777 & n14053 ) | ( n13923 & n14053 ) ;
  assign n14056 = n6789 & ~n13954 ;
  assign n14057 = ( n6789 & n14045 ) | ( n6789 & ~n14056 ) | ( n14045 & ~n14056 ) ;
  assign n14058 = ( n10944 & n10952 ) | ( n10944 & n13953 ) | ( n10952 & n13953 ) ;
  assign n14059 = n14058 ^ n10965 ^ n10952 ;
  assign n14060 = n8086 & n10944 ;
  assign n14061 = ( n8088 & n10952 ) | ( n8088 & n14060 ) | ( n10952 & n14060 ) ;
  assign n14062 = n14060 | n14061 ;
  assign n14063 = ( n8090 & n10965 ) | ( n8090 & n14060 ) | ( n10965 & n14060 ) ;
  assign n14064 = n14062 | n14063 ;
  assign n14065 = n8089 & n14059 ;
  assign n14066 = n14064 | n14065 ;
  assign n14067 = n8086 & n10952 ;
  assign n14068 = n14066 ^ x2 ^ 1'b0 ;
  assign n14069 = ( n13816 & n13960 ) | ( n13816 & n14068 ) | ( n13960 & n14068 ) ;
  assign n14070 = ( n8088 & n10965 ) | ( n8088 & n14067 ) | ( n10965 & n14067 ) ;
  assign n14071 = n14067 | n14070 ;
  assign n14072 = n6788 & ~n10944 ;
  assign n14073 = ( n6788 & n13945 ) | ( n6788 & ~n14072 ) | ( n13945 & ~n14072 ) ;
  assign n14074 = ( n6342 & ~n13724 ) | ( n6342 & n14073 ) | ( ~n13724 & n14073 ) ;
  assign n14075 = ( n8090 & n10957 ) | ( n8090 & n14067 ) | ( n10957 & n14067 ) ;
  assign n14076 = n14071 | n14075 ;
  assign n14077 = n14073 ^ n13724 ^ n6342 ;
  assign n14078 = ( n10952 & n10965 ) | ( n10952 & n14058 ) | ( n10965 & n14058 ) ;
  assign n14079 = n14078 ^ n10965 ^ n10957 ;
  assign n14080 = n8089 & n14079 ;
  assign n14081 = n14076 | n14080 ;
  assign n14082 = n14081 ^ x2 ^ 1'b0 ;
  assign n14083 = ( n13903 & n14069 ) | ( n13903 & n14082 ) | ( n14069 & n14082 ) ;
  assign n14084 = n6901 & n10965 ;
  assign n14085 = ( n6906 & n10952 ) | ( n6906 & n14084 ) | ( n10952 & n14084 ) ;
  assign n14086 = n14084 | n14085 ;
  assign n14087 = n7829 & n10952 ;
  assign n14088 = ( n6907 & n10957 ) | ( n6907 & n14084 ) | ( n10957 & n14084 ) ;
  assign n14089 = n14086 | n14088 ;
  assign n14090 = ( n6918 & n14079 ) | ( n6918 & n14089 ) | ( n14079 & n14089 ) ;
  assign n14091 = n14089 | n14090 ;
  assign n14092 = n14091 ^ x29 ^ 1'b0 ;
  assign n14093 = ( n7833 & n10944 ) | ( n7833 & n14087 ) | ( n10944 & n14087 ) ;
  assign n14094 = n14087 | n14093 ;
  assign n14095 = ( n7834 & n10965 ) | ( n7834 & n14087 ) | ( n10965 & n14087 ) ;
  assign n14096 = n14094 | n14095 ;
  assign n14097 = n7838 & n14059 ;
  assign n14098 = n14096 | n14097 ;
  assign n14099 = ( n6342 & ~n6779 ) | ( n6342 & n14057 ) | ( ~n6779 & n14057 ) ;
  assign n14100 = n14098 ^ x11 ^ 1'b0 ;
  assign n14101 = n14057 ^ n6779 ^ n6342 ;
  assign n14102 = n14100 ^ n13999 ^ n13681 ;
  assign n14103 = ( n13681 & n13999 ) | ( n13681 & n14100 ) | ( n13999 & n14100 ) ;
  assign n14104 = n14092 ^ n14077 ^ n13728 ;
  assign n14105 = n7196 & n14059 ;
  assign n14106 = ( n13728 & ~n14077 ) | ( n13728 & n14092 ) | ( ~n14077 & n14092 ) ;
  assign n14107 = n7188 & n10965 ;
  assign n14108 = n14106 ^ n14101 ^ n14074 ;
  assign n14109 = ( n14074 & ~n14101 ) | ( n14074 & n14106 ) | ( ~n14101 & n14106 ) ;
  assign n14110 = ( n7190 & n10944 ) | ( n7190 & n14107 ) | ( n10944 & n14107 ) ;
  assign n14111 = ( n7192 & n10952 ) | ( n7192 & n14107 ) | ( n10952 & n14107 ) ;
  assign n14112 = n14107 | n14110 ;
  assign n14113 = n14111 | n14112 ;
  assign n14114 = n14105 | n14113 ;
  assign n14115 = n14114 ^ x23 ^ 1'b0 ;
  assign n14116 = ( ~n13710 & n14029 ) | ( ~n13710 & n14115 ) | ( n14029 & n14115 ) ;
  assign n14117 = n14115 ^ n14029 ^ n13710 ;
  assign n14118 = n7339 & n10952 ;
  assign n14119 = ( n7337 & n10965 ) | ( n7337 & n14118 ) | ( n10965 & n14118 ) ;
  assign n14120 = n14118 | n14119 ;
  assign n14121 = ( n7338 & n10944 ) | ( n7338 & n14118 ) | ( n10944 & n14118 ) ;
  assign n14122 = n14120 | n14121 ;
  assign n14123 = n7340 & n14059 ;
  assign n14124 = n14122 | n14123 ;
  assign n14125 = n14124 ^ x20 ^ 1'b0 ;
  assign n14126 = ( ~n13757 & n14040 ) | ( ~n13757 & n14125 ) | ( n14040 & n14125 ) ;
  assign n14127 = n14125 ^ n14040 ^ n13757 ;
  assign n14128 = n8029 & n10952 ;
  assign n14129 = ( n8037 & n10944 ) | ( n8037 & n14128 ) | ( n10944 & n14128 ) ;
  assign n14130 = n14128 | n14129 ;
  assign n14131 = ( n8033 & n10965 ) | ( n8033 & n14128 ) | ( n10965 & n14128 ) ;
  assign n14132 = n14130 | n14131 ;
  assign n14133 = n8034 & n14059 ;
  assign n14134 = n14132 | n14133 ;
  assign n14135 = n14134 ^ x5 ^ 1'b0 ;
  assign n14136 = ( ~n13819 & n13990 ) | ( ~n13819 & n14135 ) | ( n13990 & n14135 ) ;
  assign n14137 = n14135 ^ n13990 ^ n13819 ;
  assign n14138 = n8029 & n10965 ;
  assign n14139 = ( n8037 & n10952 ) | ( n8037 & n14138 ) | ( n10952 & n14138 ) ;
  assign n14140 = n14138 | n14139 ;
  assign n14141 = ( n8033 & n10957 ) | ( n8033 & n14138 ) | ( n10957 & n14138 ) ;
  assign n14142 = n14140 | n14141 ;
  assign n14143 = n8034 & n14079 ;
  assign n14144 = n14142 | n14143 ;
  assign n14145 = n14144 ^ x5 ^ 1'b0 ;
  assign n14146 = ( n13922 & n14136 ) | ( n13922 & n14145 ) | ( n14136 & n14145 ) ;
  assign n14147 = n14145 ^ n14136 ^ n13922 ;
  assign n14148 = n6901 & n10952 ;
  assign n14149 = ( n6906 & n10944 ) | ( n6906 & n14148 ) | ( n10944 & n14148 ) ;
  assign n14150 = n14148 | n14149 ;
  assign n14151 = ( n6907 & n10965 ) | ( n6907 & n14148 ) | ( n10965 & n14148 ) ;
  assign n14152 = n14150 | n14151 ;
  assign n14153 = n6918 & n14059 ;
  assign n14154 = n14152 | n14153 ;
  assign n14155 = n14154 ^ x29 ^ 1'b0 ;
  assign n14156 = ( n13727 & n13986 ) | ( n13727 & n14155 ) | ( n13986 & n14155 ) ;
  assign n14157 = n14155 ^ n13986 ^ n13727 ;
  assign n14158 = n7037 & n10957 ;
  assign n14159 = ( n7036 & n10965 ) | ( n7036 & n14158 ) | ( n10965 & n14158 ) ;
  assign n14160 = n14158 | n14159 ;
  assign n14161 = ( n7052 & n10952 ) | ( n7052 & n14158 ) | ( n10952 & n14158 ) ;
  assign n14162 = n14160 | n14161 ;
  assign n14163 = n7035 & n14079 ;
  assign n14164 = n14162 | n14163 ;
  assign n14165 = n14164 ^ x26 ^ 1'b0 ;
  assign n14166 = n14165 ^ n13932 ^ n13692 ;
  assign n14167 = ( n13692 & n13932 ) | ( n13692 & n14165 ) | ( n13932 & n14165 ) ;
  assign n14168 = n7829 & n10965 ;
  assign n14169 = ( n7833 & n10952 ) | ( n7833 & n14168 ) | ( n10952 & n14168 ) ;
  assign n14170 = n14168 | n14169 ;
  assign n14171 = ( n7834 & n10957 ) | ( n7834 & n14168 ) | ( n10957 & n14168 ) ;
  assign n14172 = n14170 | n14171 ;
  assign n14173 = n7838 & n14079 ;
  assign n14174 = n14172 | n14173 ;
  assign n14175 = n14174 ^ x11 ^ 1'b0 ;
  assign n14176 = n14175 ^ n14103 ^ n13947 ;
  assign n14177 = ( n13947 & n14103 ) | ( n13947 & n14175 ) | ( n14103 & n14175 ) ;
  assign n14178 = n7669 & n10952 ;
  assign n14179 = ( n7674 & n10944 ) | ( n7674 & n14178 ) | ( n10944 & n14178 ) ;
  assign n14180 = n14178 | n14179 ;
  assign n14181 = ( n7667 & n10965 ) | ( n7667 & n14178 ) | ( n10965 & n14178 ) ;
  assign n14182 = n14180 | n14181 ;
  assign n14183 = n7666 & n14059 ;
  assign n14184 = n14182 | n14183 ;
  assign n14185 = n14184 ^ x14 ^ 1'b0 ;
  assign n14186 = n14185 ^ n13768 ^ n13738 ;
  assign n14187 = ( ~n13738 & n13768 ) | ( ~n13738 & n14185 ) | ( n13768 & n14185 ) ;
  assign n14188 = n7037 & n10965 ;
  assign n14189 = ( n7036 & n10952 ) | ( n7036 & n14188 ) | ( n10952 & n14188 ) ;
  assign n14190 = n14188 | n14189 ;
  assign n14191 = ( n7052 & n10944 ) | ( n7052 & n14188 ) | ( n10944 & n14188 ) ;
  assign n14192 = n14190 | n14191 ;
  assign n14193 = n7035 & n14059 ;
  assign n14194 = n14192 | n14193 ;
  assign n14195 = n14194 ^ x26 ^ 1'b0 ;
  assign n14196 = n14195 ^ n14010 ^ n13691 ;
  assign n14197 = ( ~n13691 & n14010 ) | ( ~n13691 & n14195 ) | ( n14010 & n14195 ) ;
  assign n14198 = n7485 & n10952 ;
  assign n14199 = ( n7486 & n10965 ) | ( n7486 & n14198 ) | ( n10965 & n14198 ) ;
  assign n14200 = n14198 | n14199 ;
  assign n14201 = ( n7493 & n10944 ) | ( n7493 & n14198 ) | ( n10944 & n14198 ) ;
  assign n14202 = n14200 | n14201 ;
  assign n14203 = n7487 & n14059 ;
  assign n14204 = n14202 | n14203 ;
  assign n14205 = n14204 ^ x17 ^ 1'b0 ;
  assign n14206 = ( ~n13789 & n14019 ) | ( ~n13789 & n14205 ) | ( n14019 & n14205 ) ;
  assign n14207 = n14205 ^ n14019 ^ n13789 ;
  assign n14208 = n7932 & n10952 ;
  assign n14209 = ( n7943 & n10944 ) | ( n7943 & n14208 ) | ( n10944 & n14208 ) ;
  assign n14210 = n14208 | n14209 ;
  assign n14211 = ( n7929 & n10965 ) | ( n7929 & n14208 ) | ( n10965 & n14208 ) ;
  assign n14212 = n14210 | n14211 ;
  assign n14213 = n6789 & ~n14059 ;
  assign n14214 = ( n7930 & n14059 ) | ( n7930 & n14212 ) | ( n14059 & n14212 ) ;
  assign n14215 = n14212 | n14214 ;
  assign n14216 = n14215 ^ x8 ^ 1'b0 ;
  assign n14217 = ( ~n13838 & n14055 ) | ( ~n13838 & n14216 ) | ( n14055 & n14216 ) ;
  assign n14218 = n14216 ^ n14055 ^ n13838 ;
  assign n14219 = n6791 & n10952 ;
  assign n14220 = ( n6790 & n10944 ) | ( n6790 & n14219 ) | ( n10944 & n14219 ) ;
  assign n14221 = ( n6788 & n10965 ) | ( n6788 & n14219 ) | ( n10965 & n14219 ) ;
  assign n14222 = n14219 | n14221 ;
  assign n14223 = n14220 | n14222 ;
  assign n14224 = ( n6789 & ~n14213 ) | ( n6789 & n14223 ) | ( ~n14213 & n14223 ) ;
  assign n14225 = n7188 & n10957 ;
  assign n14226 = ( n7190 & n10952 ) | ( n7190 & n14225 ) | ( n10952 & n14225 ) ;
  assign n14227 = n14225 | n14226 ;
  assign n14228 = ( n7192 & n10965 ) | ( n7192 & n14225 ) | ( n10965 & n14225 ) ;
  assign n14229 = n14227 | n14228 ;
  assign n14230 = n7196 & n14079 ;
  assign n14231 = n14229 | n14230 ;
  assign n14232 = n14231 ^ x23 ^ 1'b0 ;
  assign n14233 = ( n13711 & n13912 ) | ( n13711 & n14232 ) | ( n13912 & n14232 ) ;
  assign n14234 = n14232 ^ n13912 ^ n13711 ;
  assign n14235 = n7339 & n10965 ;
  assign n14236 = ( n7337 & n10957 ) | ( n7337 & n14235 ) | ( n10957 & n14235 ) ;
  assign n14237 = n14235 | n14236 ;
  assign n14238 = ( n7338 & n10952 ) | ( n7338 & n14235 ) | ( n10952 & n14235 ) ;
  assign n14239 = n14237 | n14238 ;
  assign n14240 = n7340 & n14079 ;
  assign n14241 = n14239 | n14240 ;
  assign n14242 = n14241 ^ x20 ^ 1'b0 ;
  assign n14243 = n14242 ^ n13873 ^ n13758 ;
  assign n14244 = ( n13758 & ~n13873 ) | ( n13758 & n14242 ) | ( ~n13873 & n14242 ) ;
  assign n14245 = n7485 & n10965 ;
  assign n14246 = ( n7486 & n10957 ) | ( n7486 & n14245 ) | ( n10957 & n14245 ) ;
  assign n14247 = n14245 | n14246 ;
  assign n14248 = ( n7493 & n10952 ) | ( n7493 & n14245 ) | ( n10952 & n14245 ) ;
  assign n14249 = n14247 | n14248 ;
  assign n14250 = n7487 & n14079 ;
  assign n14251 = n14249 | n14250 ;
  assign n14252 = n14251 ^ x17 ^ 1'b0 ;
  assign n14253 = n14252 ^ n13862 ^ n13788 ;
  assign n14254 = ( n13788 & n13862 ) | ( n13788 & n14252 ) | ( n13862 & n14252 ) ;
  assign n14255 = n7669 & n10965 ;
  assign n14256 = ( n7674 & n10952 ) | ( n7674 & n14255 ) | ( n10952 & n14255 ) ;
  assign n14257 = n14255 | n14256 ;
  assign n14258 = ( n7667 & n10957 ) | ( n7667 & n14255 ) | ( n10957 & n14255 ) ;
  assign n14259 = n14257 | n14258 ;
  assign n14260 = n7666 & n14079 ;
  assign n14261 = n14259 | n14260 ;
  assign n14262 = n14261 ^ x14 ^ 1'b0 ;
  assign n14263 = n14262 ^ n13888 ^ n13737 ;
  assign n14264 = ( n13737 & n13888 ) | ( n13737 & n14262 ) | ( n13888 & n14262 ) ;
  assign n14265 = n7932 & n10965 ;
  assign n14266 = ( n7943 & n10952 ) | ( n7943 & n14265 ) | ( n10952 & n14265 ) ;
  assign n14267 = n14265 | n14266 ;
  assign n14268 = ( n7929 & n10957 ) | ( n7929 & n14265 ) | ( n10957 & n14265 ) ;
  assign n14269 = n14267 | n14268 ;
  assign n14270 = ( n7930 & n14079 ) | ( n7930 & n14269 ) | ( n14079 & n14269 ) ;
  assign n14271 = n6789 & n14079 ;
  assign n14272 = n14269 | n14270 ;
  assign n14273 = ( n6791 & n10965 ) | ( n6791 & n14271 ) | ( n10965 & n14271 ) ;
  assign n14274 = n14271 | n14273 ;
  assign n14275 = ( n6790 & n10952 ) | ( n6790 & n14271 ) | ( n10952 & n14271 ) ;
  assign n14276 = n14272 ^ x8 ^ 1'b0 ;
  assign n14277 = ( n13893 & n14217 ) | ( n13893 & n14276 ) | ( n14217 & n14276 ) ;
  assign n14278 = n14276 ^ n14217 ^ n13893 ;
  assign n14279 = n14274 | n14275 ;
  assign n14280 = ( n10957 & n10965 ) | ( n10957 & n14078 ) | ( n10965 & n14078 ) ;
  assign n14281 = n14280 ^ n10957 ^ n10954 ;
  assign n14282 = n7669 & n10957 ;
  assign n14283 = ( n7674 & n10965 ) | ( n7674 & n14282 ) | ( n10965 & n14282 ) ;
  assign n14284 = ( ~n10954 & n10957 ) | ( ~n10954 & n14280 ) | ( n10957 & n14280 ) ;
  assign n14285 = n14282 | n14283 ;
  assign n14286 = ( n7667 & ~n10954 ) | ( n7667 & n14282 ) | ( ~n10954 & n14282 ) ;
  assign n14287 = n14285 | n14286 ;
  assign n14288 = n8029 & n10957 ;
  assign n14289 = n7666 & ~n14281 ;
  assign n14290 = n14287 | n14289 ;
  assign n14291 = n14290 ^ x14 ^ 1'b0 ;
  assign n14292 = ( n13887 & ~n14020 ) | ( n13887 & n14291 ) | ( ~n14020 & n14291 ) ;
  assign n14293 = n14291 ^ n14020 ^ n13887 ;
  assign n14294 = ( n8037 & n10965 ) | ( n8037 & n14288 ) | ( n10965 & n14288 ) ;
  assign n14295 = n14288 | n14294 ;
  assign n14296 = ( n8033 & ~n10954 ) | ( n8033 & n14288 ) | ( ~n10954 & n14288 ) ;
  assign n14297 = n14295 | n14296 ;
  assign n14298 = n8034 & ~n14281 ;
  assign n14299 = n14297 | n14298 ;
  assign n14300 = n7932 & n10957 ;
  assign n14301 = ( n7943 & n10965 ) | ( n7943 & n14300 ) | ( n10965 & n14300 ) ;
  assign n14302 = n14299 ^ x5 ^ 1'b0 ;
  assign n14303 = n14300 | n14301 ;
  assign n14304 = ( n7929 & ~n10954 ) | ( n7929 & n14300 ) | ( ~n10954 & n14300 ) ;
  assign n14305 = n14303 | n14304 ;
  assign n14306 = n14302 ^ n14146 ^ n14054 ;
  assign n14307 = ( ~n14054 & n14146 ) | ( ~n14054 & n14302 ) | ( n14146 & n14302 ) ;
  assign n14308 = n7930 & ~n14281 ;
  assign n14309 = ( n8086 & n8090 ) | ( n8086 & n10969 ) | ( n8090 & n10969 ) ;
  assign n14310 = n14305 & ~n14308 ;
  assign n14311 = n8084 | n14309 ;
  assign n14312 = n14310 ^ n14308 ^ x8 ;
  assign n14313 = ( n10954 & n10959 ) | ( n10954 & ~n14284 ) | ( n10959 & ~n14284 ) ;
  assign n14314 = n14312 ^ n14277 ^ n13998 ;
  assign n14315 = ( n13998 & n14277 ) | ( n13998 & n14312 ) | ( n14277 & n14312 ) ;
  assign n14316 = n8086 & n10965 ;
  assign n14317 = ( n8088 & n10957 ) | ( n8088 & n14316 ) | ( n10957 & n14316 ) ;
  assign n14318 = n14316 | n14317 ;
  assign n14319 = ( n8090 & ~n10954 ) | ( n8090 & n14316 ) | ( ~n10954 & n14316 ) ;
  assign n14320 = n14318 | n14319 ;
  assign n14321 = n8089 & ~n14281 ;
  assign n14322 = n14320 & ~n14321 ;
  assign n14323 = n14322 ^ n14321 ^ x2 ;
  assign n14324 = n14323 ^ n14083 ^ n13989 ;
  assign n14325 = ( ~n13989 & n14083 ) | ( ~n13989 & n14323 ) | ( n14083 & n14323 ) ;
  assign n14326 = n7932 & ~n10954 ;
  assign n14327 = n14284 ^ n10959 ^ n10954 ;
  assign n14328 = ( n7943 & n10957 ) | ( n7943 & n14326 ) | ( n10957 & n14326 ) ;
  assign n14329 = n14326 | n14328 ;
  assign n14330 = ( n7929 & ~n10959 ) | ( n7929 & n14326 ) | ( ~n10959 & n14326 ) ;
  assign n14331 = n14329 | n14330 ;
  assign n14332 = n14311 ^ x2 ^ 1'b0 ;
  assign n14333 = ( n7930 & n14327 ) | ( n7930 & n14331 ) | ( n14327 & n14331 ) ;
  assign n14334 = n14331 | n14333 ;
  assign n14335 = n14334 ^ x8 ^ 1'b0 ;
  assign n14336 = ( n14102 & n14315 ) | ( n14102 & n14335 ) | ( n14315 & n14335 ) ;
  assign n14337 = n14335 ^ n14315 ^ n14102 ;
  assign n14338 = n7829 & n10957 ;
  assign n14339 = ( n7833 & n10965 ) | ( n7833 & n14338 ) | ( n10965 & n14338 ) ;
  assign n14340 = n14338 | n14339 ;
  assign n14341 = ( n7834 & ~n10954 ) | ( n7834 & n14338 ) | ( ~n10954 & n14338 ) ;
  assign n14342 = n14340 | n14341 ;
  assign n14343 = n7838 & ~n14281 ;
  assign n14344 = n14342 | n14343 ;
  assign n14345 = n14344 ^ x11 ^ 1'b0 ;
  assign n14346 = n14345 ^ n14177 ^ n13973 ;
  assign n14347 = ( n13973 & n14177 ) | ( n13973 & n14345 ) | ( n14177 & n14345 ) ;
  assign n14348 = n8029 & ~n10954 ;
  assign n14349 = n7932 & ~n10959 ;
  assign n14350 = ( n7943 & ~n10954 ) | ( n7943 & n14349 ) | ( ~n10954 & n14349 ) ;
  assign n14351 = n14349 | n14350 ;
  assign n14352 = ( n7929 & n10951 ) | ( n7929 & n14349 ) | ( n10951 & n14349 ) ;
  assign n14353 = n14351 | n14352 ;
  assign n14354 = ( n8037 & n10957 ) | ( n8037 & n14348 ) | ( n10957 & n14348 ) ;
  assign n14355 = n14348 | n14354 ;
  assign n14356 = ( n8033 & ~n10959 ) | ( n8033 & n14348 ) | ( ~n10959 & n14348 ) ;
  assign n14357 = n14355 | n14356 ;
  assign n14358 = n8034 & n14327 ;
  assign n14359 = n14357 | n14358 ;
  assign n14360 = n14359 ^ x5 ^ 1'b0 ;
  assign n14361 = n14360 ^ n14307 ^ n14218 ;
  assign n14362 = ( ~n14218 & n14307 ) | ( ~n14218 & n14360 ) | ( n14307 & n14360 ) ;
  assign n14363 = n14313 ^ n10959 ^ n10951 ;
  assign n14364 = ( n7930 & n14353 ) | ( n7930 & n14363 ) | ( n14353 & n14363 ) ;
  assign n14365 = n14353 | n14364 ;
  assign n14366 = n14365 ^ x8 ^ 1'b0 ;
  assign n14367 = n14366 ^ n14336 ^ n14176 ;
  assign n14368 = ( n14176 & n14336 ) | ( n14176 & n14366 ) | ( n14336 & n14366 ) ;
  assign n14369 = n8086 & n10957 ;
  assign n14370 = ( n8088 & ~n10954 ) | ( n8088 & n14369 ) | ( ~n10954 & n14369 ) ;
  assign n14371 = n14369 | n14370 ;
  assign n14372 = ( n8090 & ~n10959 ) | ( n8090 & n14369 ) | ( ~n10959 & n14369 ) ;
  assign n14373 = n14371 | n14372 ;
  assign n14374 = ( n8089 & n14327 ) | ( n8089 & n14373 ) | ( n14327 & n14373 ) ;
  assign n14375 = n14373 | n14374 ;
  assign n14376 = n14375 ^ x2 ^ 1'b0 ;
  assign n14377 = ( ~n14137 & n14325 ) | ( ~n14137 & n14376 ) | ( n14325 & n14376 ) ;
  assign n14378 = n14376 ^ n14325 ^ n14137 ;
  assign n14379 = n8029 & ~n10959 ;
  assign n14380 = ( n8037 & ~n10954 ) | ( n8037 & n14379 ) | ( ~n10954 & n14379 ) ;
  assign n14381 = n14379 | n14380 ;
  assign n14382 = ( n8033 & n10951 ) | ( n8033 & n14379 ) | ( n10951 & n14379 ) ;
  assign n14383 = n14381 | n14382 ;
  assign n14384 = n8034 & n14363 ;
  assign n14385 = n14383 | n14384 ;
  assign n14386 = n14385 ^ x5 ^ 1'b0 ;
  assign n14387 = ( n14278 & n14362 ) | ( n14278 & n14386 ) | ( n14362 & n14386 ) ;
  assign n14388 = n14386 ^ n14362 ^ n14278 ;
  assign n14389 = n7829 & ~n10959 ;
  assign n14390 = ( n7833 & ~n10954 ) | ( n7833 & n14389 ) | ( ~n10954 & n14389 ) ;
  assign n14391 = n14389 | n14390 ;
  assign n14392 = ( n7834 & n10951 ) | ( n7834 & n14389 ) | ( n10951 & n14389 ) ;
  assign n14393 = n14391 | n14392 ;
  assign n14394 = n7838 & n14363 ;
  assign n14395 = n14393 | n14394 ;
  assign n14396 = n14395 ^ x11 ^ 1'b0 ;
  assign n14397 = ( n14187 & n14263 ) | ( n14187 & n14396 ) | ( n14263 & n14396 ) ;
  assign n14398 = n14396 ^ n14263 ^ n14187 ;
  assign n14399 = n7829 & ~n10954 ;
  assign n14400 = ( n7833 & n10957 ) | ( n7833 & n14399 ) | ( n10957 & n14399 ) ;
  assign n14401 = n14399 | n14400 ;
  assign n14402 = ( ~n10951 & n10959 ) | ( ~n10951 & n14313 ) | ( n10959 & n14313 ) ;
  assign n14403 = ( n7834 & ~n10959 ) | ( n7834 & n14399 ) | ( ~n10959 & n14399 ) ;
  assign n14404 = n14401 | n14403 ;
  assign n14405 = n7838 & n14327 ;
  assign n14406 = n14404 | n14405 ;
  assign n14407 = n14406 ^ x11 ^ 1'b0 ;
  assign n14408 = ( n13974 & ~n14186 ) | ( n13974 & n14407 ) | ( ~n14186 & n14407 ) ;
  assign n14409 = n14407 ^ n14186 ^ n13974 ;
  assign n14410 = n8086 & ~n10954 ;
  assign n14411 = ( n8088 & ~n10959 ) | ( n8088 & n14410 ) | ( ~n10959 & n14410 ) ;
  assign n14412 = n14410 | n14411 ;
  assign n14413 = ( n8090 & n10951 ) | ( n8090 & n14410 ) | ( n10951 & n14410 ) ;
  assign n14414 = n14412 | n14413 ;
  assign n14415 = ( n8089 & n14363 ) | ( n8089 & n14414 ) | ( n14363 & n14414 ) ;
  assign n14416 = n14414 | n14415 ;
  assign n14417 = n14416 ^ x2 ^ 1'b0 ;
  assign n14418 = n14417 ^ n14377 ^ n14147 ;
  assign n14419 = ( n14147 & n14377 ) | ( n14147 & n14417 ) | ( n14377 & n14417 ) ;
  assign n14420 = n7932 & n10951 ;
  assign n14421 = ( n7929 & ~n10956 ) | ( n7929 & n14420 ) | ( ~n10956 & n14420 ) ;
  assign n14422 = ( n7943 & ~n10959 ) | ( n7943 & n14420 ) | ( ~n10959 & n14420 ) ;
  assign n14423 = n14420 | n14422 ;
  assign n14424 = n14421 | n14423 ;
  assign n14425 = n14402 ^ n10956 ^ n10951 ;
  assign n14426 = ( n7930 & n14424 ) | ( n7930 & n14425 ) | ( n14424 & n14425 ) ;
  assign n14427 = n14424 | n14426 ;
  assign n14428 = n14427 ^ x8 ^ 1'b0 ;
  assign n14429 = n14428 ^ n14368 ^ n14346 ;
  assign n14430 = n7932 & ~n10956 ;
  assign n14431 = ( n14346 & n14368 ) | ( n14346 & n14428 ) | ( n14368 & n14428 ) ;
  assign n14432 = ( n7943 & n10951 ) | ( n7943 & n14430 ) | ( n10951 & n14430 ) ;
  assign n14433 = n14430 | n14432 ;
  assign n14434 = ( n7929 & ~n10968 ) | ( n7929 & n14430 ) | ( ~n10968 & n14430 ) ;
  assign n14435 = ( ~n10951 & n10956 ) | ( ~n10951 & n14402 ) | ( n10956 & n14402 ) ;
  assign n14436 = n14435 ^ n10968 ^ n10956 ;
  assign n14437 = n14433 | n14434 ;
  assign n14438 = n7930 & ~n14436 ;
  assign n14439 = n14437 | n14438 ;
  assign n14440 = n14439 ^ x8 ^ 1'b0 ;
  assign n14441 = n14440 ^ n14409 ^ n14347 ;
  assign n14442 = ( n14347 & ~n14409 ) | ( n14347 & n14440 ) | ( ~n14409 & n14440 ) ;
  assign n14443 = n7829 & n10951 ;
  assign n14444 = ( n7833 & ~n10959 ) | ( n7833 & n14443 ) | ( ~n10959 & n14443 ) ;
  assign n14445 = n14443 | n14444 ;
  assign n14446 = ( n7834 & ~n10956 ) | ( n7834 & n14443 ) | ( ~n10956 & n14443 ) ;
  assign n14447 = n14445 | n14446 ;
  assign n14448 = n7838 & n14425 ;
  assign n14449 = n14447 | n14448 ;
  assign n14450 = n14449 ^ x11 ^ 1'b0 ;
  assign n14451 = n14450 ^ n14293 ^ n14264 ;
  assign n14452 = ( n14264 & ~n14293 ) | ( n14264 & n14450 ) | ( ~n14293 & n14450 ) ;
  assign n14453 = n8086 & ~n10959 ;
  assign n14454 = ( n8088 & n10951 ) | ( n8088 & n14453 ) | ( n10951 & n14453 ) ;
  assign n14455 = n14453 | n14454 ;
  assign n14456 = ( n8090 & ~n10956 ) | ( n8090 & n14453 ) | ( ~n10956 & n14453 ) ;
  assign n14457 = n14455 | n14456 ;
  assign n14458 = ( n8089 & n14425 ) | ( n8089 & n14457 ) | ( n14425 & n14457 ) ;
  assign n14459 = n14457 | n14458 ;
  assign n14460 = n14459 ^ x2 ^ 1'b0 ;
  assign n14461 = n14460 ^ n14419 ^ n14306 ;
  assign n14462 = ( ~n14306 & n14419 ) | ( ~n14306 & n14460 ) | ( n14419 & n14460 ) ;
  assign n14463 = ( n10956 & n10968 ) | ( n10956 & n14435 ) | ( n10968 & n14435 ) ;
  assign n14464 = ( n10967 & n10968 ) | ( n10967 & n14463 ) | ( n10968 & n14463 ) ;
  assign n14465 = ( n10967 & ~n10969 ) | ( n10967 & n14464 ) | ( ~n10969 & n14464 ) ;
  assign n14466 = n14464 ^ n10969 ^ n10967 ;
  assign n14467 = n7932 & ~n10967 ;
  assign n14468 = n14465 ^ n10963 ^ 1'b0 ;
  assign n14469 = ( n7943 & ~n10968 ) | ( n7943 & n14467 ) | ( ~n10968 & n14467 ) ;
  assign n14470 = n14467 | n14469 ;
  assign n14471 = ( n7929 & n10969 ) | ( n7929 & n14467 ) | ( n10969 & n14467 ) ;
  assign n14472 = n14470 | n14471 ;
  assign n14473 = n7930 & n14466 ;
  assign n14474 = n14472 | n14473 ;
  assign n14475 = n14474 ^ x8 ^ 1'b0 ;
  assign n14476 = ( n14397 & ~n14451 ) | ( n14397 & n14475 ) | ( ~n14451 & n14475 ) ;
  assign n14477 = n14475 ^ n14451 ^ n14397 ;
  assign n14478 = n14463 ^ n10968 ^ n10967 ;
  assign n14479 = n7932 & ~n10968 ;
  assign n14480 = ( n7943 & ~n10956 ) | ( n7943 & n14479 ) | ( ~n10956 & n14479 ) ;
  assign n14481 = n14479 | n14480 ;
  assign n14482 = ( n7929 & ~n10967 ) | ( n7929 & n14479 ) | ( ~n10967 & n14479 ) ;
  assign n14483 = n14481 | n14482 ;
  assign n14484 = n7930 & ~n14478 ;
  assign n14485 = n14483 | n14484 ;
  assign n14486 = n14485 ^ x8 ^ 1'b0 ;
  assign n14487 = n14486 ^ n14408 ^ n14398 ;
  assign n14488 = ( n14398 & n14408 ) | ( n14398 & n14486 ) | ( n14408 & n14486 ) ;
  assign n14489 = ( n8029 & n8033 ) | ( n8029 & n10969 ) | ( n8033 & n10969 ) ;
  assign n14490 = n8033 | n14489 ;
  assign n14491 = ( n8033 & n8037 ) | ( n8033 & ~n10967 ) | ( n8037 & ~n10967 ) ;
  assign n14492 = n14490 | n14491 ;
  assign n14493 = n8034 & n14468 ;
  assign n14494 = n14492 | n14493 ;
  assign n14495 = ( n12655 & ~n14477 ) | ( n12655 & n14488 ) | ( ~n14477 & n14488 ) ;
  assign n14496 = n14488 ^ n14477 ^ n12655 ;
  assign n14497 = n8029 & ~n10967 ;
  assign n14498 = ( n8037 & ~n10968 ) | ( n8037 & n14497 ) | ( ~n10968 & n14497 ) ;
  assign n14499 = n14497 | n14498 ;
  assign n14500 = ( n8033 & n10969 ) | ( n8033 & n14497 ) | ( n10969 & n14497 ) ;
  assign n14501 = n14499 | n14500 ;
  assign n14502 = n8034 & n14466 ;
  assign n14503 = n14501 | n14502 ;
  assign n14504 = n14494 ^ x5 ^ 1'b0 ;
  assign n14505 = n14503 ^ x5 ^ 1'b0 ;
  assign n14506 = ( n12257 & n14429 ) | ( n12257 & n14505 ) | ( n14429 & n14505 ) ;
  assign n14507 = n14505 ^ n14429 ^ n12257 ;
  assign n14508 = n14504 ^ n14441 ^ n14431 ;
  assign n14509 = ( n14431 & ~n14441 ) | ( n14431 & n14504 ) | ( ~n14441 & n14504 ) ;
  assign n14510 = n8029 & n10951 ;
  assign n14511 = ( n8037 & ~n10959 ) | ( n8037 & n14510 ) | ( ~n10959 & n14510 ) ;
  assign n14512 = n14510 | n14511 ;
  assign n14513 = ( n8033 & ~n10956 ) | ( n8033 & n14510 ) | ( ~n10956 & n14510 ) ;
  assign n14514 = n14512 | n14513 ;
  assign n14515 = n8034 & n14425 ;
  assign n14516 = n14514 | n14515 ;
  assign n14517 = n14516 ^ x5 ^ 1'b0 ;
  assign n14518 = n14517 ^ n14387 ^ n14314 ;
  assign n14519 = ( n14314 & n14387 ) | ( n14314 & n14517 ) | ( n14387 & n14517 ) ;
  assign n14520 = n8029 & ~n10956 ;
  assign n14521 = ( n8037 & n10951 ) | ( n8037 & n14520 ) | ( n10951 & n14520 ) ;
  assign n14522 = n14520 | n14521 ;
  assign n14523 = ( n8033 & ~n10968 ) | ( n8033 & n14520 ) | ( ~n10968 & n14520 ) ;
  assign n14524 = n14522 | n14523 ;
  assign n14525 = n8034 & ~n14436 ;
  assign n14526 = n14524 | n14525 ;
  assign n14527 = n14526 ^ x5 ^ 1'b0 ;
  assign n14528 = ( n14337 & n14519 ) | ( n14337 & n14527 ) | ( n14519 & n14527 ) ;
  assign n14529 = n14527 ^ n14519 ^ n14337 ;
  assign n14530 = n8029 & ~n10968 ;
  assign n14531 = ( n8037 & ~n10956 ) | ( n8037 & n14530 ) | ( ~n10956 & n14530 ) ;
  assign n14532 = n14530 | n14531 ;
  assign n14533 = ( n8033 & ~n10967 ) | ( n8033 & n14530 ) | ( ~n10967 & n14530 ) ;
  assign n14534 = n14532 | n14533 ;
  assign n14535 = n8034 & ~n14478 ;
  assign n14536 = n14534 | n14535 ;
  assign n14537 = n14536 ^ x5 ^ 1'b0 ;
  assign n14538 = n14537 ^ n14528 ^ n14367 ;
  assign n14539 = ( n14367 & n14528 ) | ( n14367 & n14537 ) | ( n14528 & n14537 ) ;
  assign n14540 = n8086 & n10951 ;
  assign n14541 = ( n8088 & ~n10956 ) | ( n8088 & n14540 ) | ( ~n10956 & n14540 ) ;
  assign n14542 = n14540 | n14541 ;
  assign n14543 = ( n8090 & ~n10968 ) | ( n8090 & n14540 ) | ( ~n10968 & n14540 ) ;
  assign n14544 = n14542 | n14543 ;
  assign n14545 = n8089 & ~n14436 ;
  assign n14546 = n14544 & ~n14545 ;
  assign n14547 = n14546 ^ n14545 ^ x2 ;
  assign n14548 = ( ~n14361 & n14462 ) | ( ~n14361 & n14547 ) | ( n14462 & n14547 ) ;
  assign n14549 = n14547 ^ n14462 ^ n14361 ;
  assign n14550 = n8086 & ~n10956 ;
  assign n14551 = ( n8088 & ~n10968 ) | ( n8088 & n14550 ) | ( ~n10968 & n14550 ) ;
  assign n14552 = n14550 | n14551 ;
  assign n14553 = ( n8090 & ~n10967 ) | ( n8090 & n14550 ) | ( ~n10967 & n14550 ) ;
  assign n14554 = n14552 | n14553 ;
  assign n14555 = n8089 & ~n14478 ;
  assign n14556 = n14554 & ~n14555 ;
  assign n14557 = n14556 ^ n14555 ^ x2 ;
  assign n14558 = ( n14388 & n14548 ) | ( n14388 & n14557 ) | ( n14548 & n14557 ) ;
  assign n14559 = n14557 ^ n14548 ^ n14388 ;
  assign n14560 = n8086 & ~n10968 ;
  assign n14561 = ( n8088 & ~n10967 ) | ( n8088 & n14560 ) | ( ~n10967 & n14560 ) ;
  assign n14562 = n14560 | n14561 ;
  assign n14563 = ( n8090 & n10969 ) | ( n8090 & n14560 ) | ( n10969 & n14560 ) ;
  assign n14564 = n14562 | n14563 ;
  assign n14565 = ( n8089 & n14466 ) | ( n8089 & n14564 ) | ( n14466 & n14564 ) ;
  assign n14566 = n14564 | n14565 ;
  assign n14567 = n14566 ^ x2 ^ 1'b0 ;
  assign n14568 = ( n14518 & n14558 ) | ( n14518 & n14567 ) | ( n14558 & n14567 ) ;
  assign n14569 = n14567 ^ n14558 ^ n14518 ;
  assign n14570 = ( n8086 & n8090 ) | ( n8086 & ~n10967 ) | ( n8090 & ~n10967 ) ;
  assign n14571 = n8090 | n14570 ;
  assign n14572 = ( n8088 & n8090 ) | ( n8088 & n10969 ) | ( n8090 & n10969 ) ;
  assign n14573 = n14571 | n14572 ;
  assign n14574 = ( n8089 & n14468 ) | ( n8089 & n14573 ) | ( n14468 & n14573 ) ;
  assign n14575 = n14573 | n14574 ;
  assign n14576 = n14575 ^ x2 ^ 1'b0 ;
  assign n14577 = ( n14529 & n14568 ) | ( n14529 & n14576 ) | ( n14568 & n14576 ) ;
  assign n14578 = n14576 ^ n14568 ^ n14529 ;
  assign n14579 = ( n14332 & n14538 ) | ( n14332 & n14577 ) | ( n14538 & n14577 ) ;
  assign n14580 = n14577 ^ n14538 ^ n14332 ;
  assign n14581 = ( n14507 & n14539 ) | ( n14507 & n14579 ) | ( n14539 & n14579 ) ;
  assign n14582 = ( n14506 & ~n14508 ) | ( n14506 & n14581 ) | ( ~n14508 & n14581 ) ;
  assign n14583 = n14581 ^ n14508 ^ n14506 ;
  assign n14584 = n14579 ^ n14539 ^ n14507 ;
  assign n14585 = n8029 | n8034 ;
  assign n14586 = n8033 | n14585 ;
  assign n14587 = ( n8033 & n8037 ) | ( n8033 & n10969 ) | ( n8037 & n10969 ) ;
  assign n14588 = n14586 | n14587 ;
  assign n14589 = n14588 ^ x5 ^ 1'b0 ;
  assign n14590 = n14589 ^ n14487 ^ n14442 ;
  assign n14591 = ( n14442 & n14487 ) | ( n14442 & n14589 ) | ( n14487 & n14589 ) ;
  assign n14592 = n7669 & ~n10954 ;
  assign n14593 = ( n7674 & n10957 ) | ( n7674 & n14592 ) | ( n10957 & n14592 ) ;
  assign n14594 = n14592 | n14593 ;
  assign n14595 = ( n7667 & ~n10959 ) | ( n7667 & n14592 ) | ( ~n10959 & n14592 ) ;
  assign n14596 = n14594 | n14595 ;
  assign n14597 = n7666 & n14327 ;
  assign n14598 = n14596 | n14597 ;
  assign n14599 = n14590 ^ n14582 ^ n14509 ;
  assign n14600 = n14598 ^ x14 ^ 1'b0 ;
  assign n14601 = ( n14509 & n14582 ) | ( n14509 & n14590 ) | ( n14582 & n14590 ) ;
  assign n14602 = n14600 ^ n14292 ^ n14207 ;
  assign n14603 = ( ~n14207 & n14292 ) | ( ~n14207 & n14600 ) | ( n14292 & n14600 ) ;
  assign n14604 = n7669 & ~n10959 ;
  assign n14605 = ( n7674 & ~n10954 ) | ( n7674 & n14604 ) | ( ~n10954 & n14604 ) ;
  assign n14606 = n14604 | n14605 ;
  assign n14607 = ( n7667 & n10951 ) | ( n7667 & n14604 ) | ( n10951 & n14604 ) ;
  assign n14608 = n14606 | n14607 ;
  assign n14609 = ( ~n14496 & n14591 ) | ( ~n14496 & n14601 ) | ( n14591 & n14601 ) ;
  assign n14610 = n14601 ^ n14591 ^ n14496 ;
  assign n14611 = ( n7929 & n7932 ) | ( n7929 & n10969 ) | ( n7932 & n10969 ) ;
  assign n14612 = n7929 | n14611 ;
  assign n14613 = ( n7929 & n7943 ) | ( n7929 & ~n10967 ) | ( n7943 & ~n10967 ) ;
  assign n14614 = n14612 | n14613 ;
  assign n14615 = n7930 & n14468 ;
  assign n14616 = n14614 | n14615 ;
  assign n14617 = n7666 & n14363 ;
  assign n14618 = n14608 | n14617 ;
  assign n14619 = n7829 & ~n10956 ;
  assign n14620 = ( n7833 & n10951 ) | ( n7833 & n14619 ) | ( n10951 & n14619 ) ;
  assign n14621 = n14619 | n14620 ;
  assign n14622 = ( n7834 & ~n10968 ) | ( n7834 & n14619 ) | ( ~n10968 & n14619 ) ;
  assign n14623 = n14621 | n14622 ;
  assign n14624 = n14616 ^ x8 ^ 1'b0 ;
  assign n14625 = n7838 & ~n14436 ;
  assign n14626 = n14618 ^ x14 ^ 1'b0 ;
  assign n14627 = n14623 | n14625 ;
  assign n14628 = n14627 ^ x11 ^ 1'b0 ;
  assign n14629 = ( n14206 & n14253 ) | ( n14206 & n14626 ) | ( n14253 & n14626 ) ;
  assign n14630 = n14626 ^ n14253 ^ n14206 ;
  assign n14631 = ( n14452 & ~n14602 ) | ( n14452 & n14628 ) | ( ~n14602 & n14628 ) ;
  assign n14632 = n14628 ^ n14602 ^ n14452 ;
  assign n14633 = n7838 & ~n14478 ;
  assign n14634 = n14632 ^ n14624 ^ n14476 ;
  assign n14635 = n7829 & ~n10968 ;
  assign n14636 = ( n14476 & n14624 ) | ( n14476 & ~n14632 ) | ( n14624 & ~n14632 ) ;
  assign n14637 = ( n7932 & n7943 ) | ( n7932 & n10969 ) | ( n7943 & n10969 ) ;
  assign n14638 = n7929 | n14637 ;
  assign n14639 = ( n7833 & ~n10956 ) | ( n7833 & n14635 ) | ( ~n10956 & n14635 ) ;
  assign n14640 = n14635 | n14639 ;
  assign n14641 = ( n7834 & ~n10967 ) | ( n7834 & n14635 ) | ( ~n10967 & n14635 ) ;
  assign n14642 = n14640 | n14641 ;
  assign n14643 = n14634 ^ n14609 ^ n14495 ;
  assign n14644 = ( n14495 & n14609 ) | ( n14495 & ~n14634 ) | ( n14609 & ~n14634 ) ;
  assign n14645 = n7930 | n7932 ;
  assign n14646 = n14638 | n14645 ;
  assign n14647 = n14646 ^ x8 ^ 1'b0 ;
  assign n14648 = n14633 | n14642 ;
  assign n14649 = n14648 ^ x11 ^ 1'b0 ;
  assign n14650 = n14649 ^ n14630 ^ n14603 ;
  assign n14651 = ( n14603 & n14630 ) | ( n14603 & n14649 ) | ( n14630 & n14649 ) ;
  assign n14652 = n14650 ^ n14647 ^ n14631 ;
  assign n14653 = ( n14631 & n14647 ) | ( n14631 & n14650 ) | ( n14647 & n14650 ) ;
  assign n14654 = ( n14636 & n14644 ) | ( n14636 & n14652 ) | ( n14644 & n14652 ) ;
  assign n14655 = n14652 ^ n14644 ^ n14636 ;
  assign n14656 = n7485 & n10957 ;
  assign n14657 = ( n7486 & ~n10954 ) | ( n7486 & n14656 ) | ( ~n10954 & n14656 ) ;
  assign n14658 = n14656 | n14657 ;
  assign n14659 = ( n7493 & n10965 ) | ( n7493 & n14656 ) | ( n10965 & n14656 ) ;
  assign n14660 = n14658 | n14659 ;
  assign n14661 = n7487 & ~n14281 ;
  assign n14662 = n14660 | n14661 ;
  assign n14663 = n14662 ^ x17 ^ 1'b0 ;
  assign n14664 = n14663 ^ n14039 ^ n13864 ;
  assign n14665 = ( n13864 & ~n14039 ) | ( n13864 & n14663 ) | ( ~n14039 & n14663 ) ;
  assign n14666 = n7669 & n10951 ;
  assign n14667 = ( n7674 & ~n10959 ) | ( n7674 & n14666 ) | ( ~n10959 & n14666 ) ;
  assign n14668 = n14666 | n14667 ;
  assign n14669 = ( n7667 & ~n10956 ) | ( n7667 & n14666 ) | ( ~n10956 & n14666 ) ;
  assign n14670 = n14668 | n14669 ;
  assign n14671 = n7666 & n14425 ;
  assign n14672 = n14670 | n14671 ;
  assign n14673 = n14672 ^ x14 ^ 1'b0 ;
  assign n14674 = n14673 ^ n14664 ^ n14254 ;
  assign n14675 = ( n14254 & ~n14664 ) | ( n14254 & n14673 ) | ( ~n14664 & n14673 ) ;
  assign n14676 = n7829 & ~n10967 ;
  assign n14677 = ( n7833 & ~n10968 ) | ( n7833 & n14676 ) | ( ~n10968 & n14676 ) ;
  assign n14678 = n14676 | n14677 ;
  assign n14679 = ( n7834 & n10969 ) | ( n7834 & n14676 ) | ( n10969 & n14676 ) ;
  assign n14680 = n14678 | n14679 ;
  assign n14681 = n7838 & n14466 ;
  assign n14682 = n14680 | n14681 ;
  assign n14683 = n14682 ^ x11 ^ 1'b0 ;
  assign n14684 = ( n14629 & ~n14674 ) | ( n14629 & n14683 ) | ( ~n14674 & n14683 ) ;
  assign n14685 = n14683 ^ n14674 ^ n14629 ;
  assign n14686 = ( n12883 & n14651 ) | ( n12883 & ~n14685 ) | ( n14651 & ~n14685 ) ;
  assign n14687 = n7669 & ~n10956 ;
  assign n14688 = n14685 ^ n14651 ^ n12883 ;
  assign n14689 = ( n7674 & n10951 ) | ( n7674 & n14687 ) | ( n10951 & n14687 ) ;
  assign n14690 = n14687 | n14689 ;
  assign n14691 = ( n7667 & ~n10968 ) | ( n7667 & n14687 ) | ( ~n10968 & n14687 ) ;
  assign n14692 = n14688 ^ n14654 ^ n14653 ;
  assign n14693 = ( n14653 & n14654 ) | ( n14653 & ~n14688 ) | ( n14654 & ~n14688 ) ;
  assign n14694 = n7485 & ~n10954 ;
  assign n14695 = ( n7829 & n7834 ) | ( n7829 & n10969 ) | ( n7834 & n10969 ) ;
  assign n14696 = n14690 | n14691 ;
  assign n14697 = n7666 & ~n14436 ;
  assign n14698 = n7834 | n14695 ;
  assign n14699 = n14696 | n14697 ;
  assign n14700 = ( n7833 & n7834 ) | ( n7833 & ~n10967 ) | ( n7834 & ~n10967 ) ;
  assign n14701 = n14698 | n14700 ;
  assign n14702 = ( n7486 & ~n10959 ) | ( n7486 & n14694 ) | ( ~n10959 & n14694 ) ;
  assign n14703 = n14694 | n14702 ;
  assign n14704 = ( n7493 & n10957 ) | ( n7493 & n14694 ) | ( n10957 & n14694 ) ;
  assign n14705 = n14703 | n14704 ;
  assign n14706 = n7487 & n14327 ;
  assign n14707 = n14705 | n14706 ;
  assign n14708 = n14707 ^ x17 ^ 1'b0 ;
  assign n14709 = ( ~n14127 & n14665 ) | ( ~n14127 & n14708 ) | ( n14665 & n14708 ) ;
  assign n14710 = n14708 ^ n14665 ^ n14127 ;
  assign n14711 = n7838 & n14468 ;
  assign n14712 = n14699 ^ x14 ^ 1'b0 ;
  assign n14713 = ( n14675 & ~n14710 ) | ( n14675 & n14712 ) | ( ~n14710 & n14712 ) ;
  assign n14714 = n14701 | n14711 ;
  assign n14715 = n14712 ^ n14710 ^ n14675 ;
  assign n14716 = n14714 ^ x11 ^ 1'b0 ;
  assign n14717 = ( n14684 & ~n14715 ) | ( n14684 & n14716 ) | ( ~n14715 & n14716 ) ;
  assign n14718 = n14716 ^ n14715 ^ n14684 ;
  assign n14719 = ( n14686 & n14693 ) | ( n14686 & ~n14718 ) | ( n14693 & ~n14718 ) ;
  assign n14720 = n14718 ^ n14693 ^ n14686 ;
  assign n14721 = n7485 & ~n10959 ;
  assign n14722 = ( n7486 & n10951 ) | ( n7486 & n14721 ) | ( n10951 & n14721 ) ;
  assign n14723 = n14721 | n14722 ;
  assign n14724 = ( n7493 & ~n10954 ) | ( n7493 & n14721 ) | ( ~n10954 & n14721 ) ;
  assign n14725 = n14723 | n14724 ;
  assign n14726 = n7487 & n14363 ;
  assign n14727 = n14725 | n14726 ;
  assign n14728 = n14727 ^ x17 ^ 1'b0 ;
  assign n14729 = ( n14126 & ~n14243 ) | ( n14126 & n14728 ) | ( ~n14243 & n14728 ) ;
  assign n14730 = n14728 ^ n14243 ^ n14126 ;
  assign n14731 = n7339 & n10957 ;
  assign n14732 = ( n7337 & ~n10954 ) | ( n7337 & n14731 ) | ( ~n10954 & n14731 ) ;
  assign n14733 = n14731 | n14732 ;
  assign n14734 = ( n7338 & n10965 ) | ( n7338 & n14731 ) | ( n10965 & n14731 ) ;
  assign n14735 = n14733 | n14734 ;
  assign n14736 = n7340 & ~n14281 ;
  assign n14737 = n14735 | n14736 ;
  assign n14738 = n14737 ^ x20 ^ 1'b0 ;
  assign n14739 = ( n13874 & ~n14030 ) | ( n13874 & n14738 ) | ( ~n14030 & n14738 ) ;
  assign n14740 = n14738 ^ n14030 ^ n13874 ;
  assign n14741 = n7669 & ~n10968 ;
  assign n14742 = ( n7674 & ~n10956 ) | ( n7674 & n14741 ) | ( ~n10956 & n14741 ) ;
  assign n14743 = n14741 | n14742 ;
  assign n14744 = ( n7667 & ~n10967 ) | ( n7667 & n14741 ) | ( ~n10967 & n14741 ) ;
  assign n14745 = n14743 | n14744 ;
  assign n14746 = n7666 & ~n14478 ;
  assign n14747 = n14745 | n14746 ;
  assign n14748 = n14747 ^ x14 ^ 1'b0 ;
  assign n14749 = n14748 ^ n14730 ^ n14709 ;
  assign n14750 = ( n14709 & ~n14730 ) | ( n14709 & n14748 ) | ( ~n14730 & n14748 ) ;
  assign n14751 = n7485 & n10951 ;
  assign n14752 = ( n7486 & ~n10956 ) | ( n7486 & n14751 ) | ( ~n10956 & n14751 ) ;
  assign n14753 = n14751 | n14752 ;
  assign n14754 = ( n7493 & ~n10959 ) | ( n7493 & n14751 ) | ( ~n10959 & n14751 ) ;
  assign n14755 = n14753 | n14754 ;
  assign n14756 = n7487 & n14425 ;
  assign n14757 = n14755 | n14756 ;
  assign n14758 = n14757 ^ x17 ^ 1'b0 ;
  assign n14759 = n14758 ^ n14740 ^ n14244 ;
  assign n14760 = ( n14244 & ~n14740 ) | ( n14244 & n14758 ) | ( ~n14740 & n14758 ) ;
  assign n14761 = n7829 | n7838 ;
  assign n14762 = ( n7829 & n7833 ) | ( n7829 & n10969 ) | ( n7833 & n10969 ) ;
  assign n14763 = n7834 | n14762 ;
  assign n14764 = n14761 | n14763 ;
  assign n14765 = n14764 ^ x11 ^ 1'b0 ;
  assign n14766 = n14765 ^ n14749 ^ n14713 ;
  assign n14767 = ( n14713 & ~n14749 ) | ( n14713 & n14765 ) | ( ~n14749 & n14765 ) ;
  assign n14768 = ( n14717 & n14719 ) | ( n14717 & ~n14766 ) | ( n14719 & ~n14766 ) ;
  assign n14769 = n7669 & ~n10967 ;
  assign n14770 = n14766 ^ n14719 ^ n14717 ;
  assign n14771 = ( n7674 & ~n10968 ) | ( n7674 & n14769 ) | ( ~n10968 & n14769 ) ;
  assign n14772 = n7666 & n14466 ;
  assign n14773 = n14769 | n14771 ;
  assign n14774 = ( n7667 & n10969 ) | ( n7667 & n14769 ) | ( n10969 & n14769 ) ;
  assign n14775 = n14773 | n14774 ;
  assign n14776 = n14772 | n14775 ;
  assign n14777 = n14776 ^ x14 ^ 1'b0 ;
  assign n14778 = ( n14729 & ~n14759 ) | ( n14729 & n14777 ) | ( ~n14759 & n14777 ) ;
  assign n14779 = n14777 ^ n14759 ^ n14729 ;
  assign n14780 = n14779 ^ n14750 ^ n13159 ;
  assign n14781 = n14780 ^ n14768 ^ n14767 ;
  assign n14782 = ( n14767 & n14768 ) | ( n14767 & ~n14780 ) | ( n14768 & ~n14780 ) ;
  assign n14783 = ( n13159 & n14750 ) | ( n13159 & ~n14779 ) | ( n14750 & ~n14779 ) ;
  assign n14784 = n7339 & ~n10954 ;
  assign n14785 = ( n7337 & ~n10959 ) | ( n7337 & n14784 ) | ( ~n10959 & n14784 ) ;
  assign n14786 = n14784 | n14785 ;
  assign n14787 = ( n7338 & n10957 ) | ( n7338 & n14784 ) | ( n10957 & n14784 ) ;
  assign n14788 = n14786 | n14787 ;
  assign n14789 = n7340 & n14327 ;
  assign n14790 = n14788 | n14789 ;
  assign n14791 = n14790 ^ x20 ^ 1'b0 ;
  assign n14792 = ( ~n14117 & n14739 ) | ( ~n14117 & n14791 ) | ( n14739 & n14791 ) ;
  assign n14793 = n14791 ^ n14739 ^ n14117 ;
  assign n14794 = n7485 & ~n10956 ;
  assign n14795 = ( n7486 & ~n10968 ) | ( n7486 & n14794 ) | ( ~n10968 & n14794 ) ;
  assign n14796 = n14794 | n14795 ;
  assign n14797 = ( n7493 & n10951 ) | ( n7493 & n14794 ) | ( n10951 & n14794 ) ;
  assign n14798 = n14796 | n14797 ;
  assign n14799 = n7487 & ~n14436 ;
  assign n14800 = n14798 | n14799 ;
  assign n14801 = n14800 ^ x17 ^ 1'b0 ;
  assign n14802 = ( n14760 & ~n14793 ) | ( n14760 & n14801 ) | ( ~n14793 & n14801 ) ;
  assign n14803 = n14801 ^ n14793 ^ n14760 ;
  assign n14804 = ( n7667 & n7669 ) | ( n7667 & n10969 ) | ( n7669 & n10969 ) ;
  assign n14805 = ( n7667 & n7674 ) | ( n7667 & ~n10967 ) | ( n7674 & ~n10967 ) ;
  assign n14806 = n7667 | n14804 ;
  assign n14807 = n14805 | n14806 ;
  assign n14808 = n7666 & n14468 ;
  assign n14809 = n14807 | n14808 ;
  assign n14810 = n14809 ^ x14 ^ 1'b0 ;
  assign n14811 = n14810 ^ n14803 ^ n14778 ;
  assign n14812 = ( n14778 & ~n14803 ) | ( n14778 & n14810 ) | ( ~n14803 & n14810 ) ;
  assign n14813 = ( n14782 & n14783 ) | ( n14782 & ~n14811 ) | ( n14783 & ~n14811 ) ;
  assign n14814 = n14811 ^ n14783 ^ n14782 ;
  assign n14815 = n7485 & ~n10968 ;
  assign n14816 = ( n7486 & ~n10967 ) | ( n7486 & n14815 ) | ( ~n10967 & n14815 ) ;
  assign n14817 = n14815 | n14816 ;
  assign n14818 = n7487 & ~n14478 ;
  assign n14819 = ( n7493 & ~n10956 ) | ( n7493 & n14815 ) | ( ~n10956 & n14815 ) ;
  assign n14820 = n14817 | n14819 ;
  assign n14821 = n7339 & ~n10959 ;
  assign n14822 = n14818 | n14820 ;
  assign n14823 = ( n7337 & n10951 ) | ( n7337 & n14821 ) | ( n10951 & n14821 ) ;
  assign n14824 = n14822 ^ x17 ^ 1'b0 ;
  assign n14825 = n14821 | n14823 ;
  assign n14826 = ( n7338 & ~n10954 ) | ( n7338 & n14821 ) | ( ~n10954 & n14821 ) ;
  assign n14827 = n14825 | n14826 ;
  assign n14828 = n7340 & n14363 ;
  assign n14829 = n14827 | n14828 ;
  assign n14830 = n14829 ^ x20 ^ 1'b0 ;
  assign n14831 = n14830 ^ n14234 ^ n14116 ;
  assign n14832 = ( n14116 & n14234 ) | ( n14116 & n14830 ) | ( n14234 & n14830 ) ;
  assign n14833 = n7666 | n7669 ;
  assign n14834 = ( n7669 & n7674 ) | ( n7669 & n10969 ) | ( n7674 & n10969 ) ;
  assign n14835 = n7667 | n14834 ;
  assign n14836 = n14833 | n14835 ;
  assign n14837 = n14836 ^ x14 ^ 1'b0 ;
  assign n14838 = ( n14792 & n14824 ) | ( n14792 & n14831 ) | ( n14824 & n14831 ) ;
  assign n14839 = n14831 ^ n14824 ^ n14792 ;
  assign n14840 = ( n14802 & n14837 ) | ( n14802 & n14839 ) | ( n14837 & n14839 ) ;
  assign n14841 = n14839 ^ n14837 ^ n14802 ;
  assign n14842 = ( n14812 & n14813 ) | ( n14812 & n14841 ) | ( n14813 & n14841 ) ;
  assign n14843 = n14841 ^ n14813 ^ n14812 ;
  assign n14844 = n7188 & ~n10954 ;
  assign n14845 = ( n7190 & n10965 ) | ( n7190 & n14844 ) | ( n10965 & n14844 ) ;
  assign n14846 = n14844 | n14845 ;
  assign n14847 = ( n7192 & n10957 ) | ( n7192 & n14844 ) | ( n10957 & n14844 ) ;
  assign n14848 = n14846 | n14847 ;
  assign n14849 = n7196 & ~n14281 ;
  assign n14850 = n14848 | n14849 ;
  assign n14851 = n14850 ^ x23 ^ 1'b0 ;
  assign n14852 = ( n13913 & n14009 ) | ( n13913 & n14851 ) | ( n14009 & n14851 ) ;
  assign n14853 = n14851 ^ n14009 ^ n13913 ;
  assign n14854 = n7339 & n10951 ;
  assign n14855 = ( n7337 & ~n10956 ) | ( n7337 & n14854 ) | ( ~n10956 & n14854 ) ;
  assign n14856 = n14854 | n14855 ;
  assign n14857 = ( n7338 & ~n10959 ) | ( n7338 & n14854 ) | ( ~n10959 & n14854 ) ;
  assign n14858 = n14856 | n14857 ;
  assign n14859 = n7340 & n14425 ;
  assign n14860 = n14858 | n14859 ;
  assign n14861 = n14860 ^ x20 ^ 1'b0 ;
  assign n14862 = n14861 ^ n14853 ^ n14233 ;
  assign n14863 = ( n14233 & n14853 ) | ( n14233 & n14861 ) | ( n14853 & n14861 ) ;
  assign n14864 = n7485 & ~n10967 ;
  assign n14865 = ( n7486 & n10969 ) | ( n7486 & n14864 ) | ( n10969 & n14864 ) ;
  assign n14866 = n14864 | n14865 ;
  assign n14867 = ( n7493 & ~n10968 ) | ( n7493 & n14864 ) | ( ~n10968 & n14864 ) ;
  assign n14868 = n14866 | n14867 ;
  assign n14869 = n7487 & n14466 ;
  assign n14870 = n14868 | n14869 ;
  assign n14871 = n14870 ^ x17 ^ 1'b0 ;
  assign n14872 = n14871 ^ n14862 ^ n14832 ;
  assign n14873 = ( n14832 & n14862 ) | ( n14832 & n14871 ) | ( n14862 & n14871 ) ;
  assign n14874 = n7188 & ~n10959 ;
  assign n14875 = ( n13523 & n14838 ) | ( n13523 & n14872 ) | ( n14838 & n14872 ) ;
  assign n14876 = n14872 ^ n14838 ^ n13523 ;
  assign n14877 = ( n7190 & n10957 ) | ( n7190 & n14874 ) | ( n10957 & n14874 ) ;
  assign n14878 = ( n7192 & ~n10954 ) | ( n7192 & n14874 ) | ( ~n10954 & n14874 ) ;
  assign n14879 = n14874 | n14877 ;
  assign n14880 = n14878 | n14879 ;
  assign n14881 = n7196 & n14327 ;
  assign n14882 = n14880 | n14881 ;
  assign n14883 = n14882 ^ x23 ^ 1'b0 ;
  assign n14884 = ( ~n14196 & n14852 ) | ( ~n14196 & n14883 ) | ( n14852 & n14883 ) ;
  assign n14885 = n14883 ^ n14852 ^ n14196 ;
  assign n14886 = ( n7485 & n7486 ) | ( n7485 & n10969 ) | ( n7486 & n10969 ) ;
  assign n14887 = n7486 | n14886 ;
  assign n14888 = n14876 ^ n14842 ^ n14840 ;
  assign n14889 = n7487 & n14468 ;
  assign n14890 = ( n14840 & n14842 ) | ( n14840 & n14876 ) | ( n14842 & n14876 ) ;
  assign n14891 = n7340 & ~n14436 ;
  assign n14892 = ( n7486 & n7493 ) | ( n7486 & ~n10967 ) | ( n7493 & ~n10967 ) ;
  assign n14893 = n14887 | n14892 ;
  assign n14894 = n7339 & ~n10956 ;
  assign n14895 = n14889 | n14893 ;
  assign n14896 = ( n7337 & ~n10968 ) | ( n7337 & n14894 ) | ( ~n10968 & n14894 ) ;
  assign n14897 = n14894 | n14896 ;
  assign n14898 = ( n7338 & n10951 ) | ( n7338 & n14894 ) | ( n10951 & n14894 ) ;
  assign n14899 = n14895 ^ x17 ^ 1'b0 ;
  assign n14900 = n14897 | n14898 ;
  assign n14901 = n14891 | n14900 ;
  assign n14902 = n14901 ^ x20 ^ 1'b0 ;
  assign n14903 = ( n14863 & ~n14885 ) | ( n14863 & n14902 ) | ( ~n14885 & n14902 ) ;
  assign n14904 = n14902 ^ n14885 ^ n14863 ;
  assign n14905 = ( n14873 & n14899 ) | ( n14873 & ~n14904 ) | ( n14899 & ~n14904 ) ;
  assign n14906 = n14904 ^ n14899 ^ n14873 ;
  assign n14907 = n14906 ^ n14890 ^ n14875 ;
  assign n14908 = ( n14875 & n14890 ) | ( n14875 & ~n14906 ) | ( n14890 & ~n14906 ) ;
  assign n14909 = n7037 & ~n10954 ;
  assign n14910 = ( n7036 & n10957 ) | ( n7036 & n14909 ) | ( n10957 & n14909 ) ;
  assign n14911 = n14909 | n14910 ;
  assign n14912 = ( n7052 & n10965 ) | ( n7052 & n14909 ) | ( n10965 & n14909 ) ;
  assign n14913 = n14911 | n14912 ;
  assign n14914 = n7035 & ~n14281 ;
  assign n14915 = n14913 | n14914 ;
  assign n14916 = n14915 ^ x26 ^ 1'b0 ;
  assign n14917 = ( n13933 & ~n13987 ) | ( n13933 & n14916 ) | ( ~n13987 & n14916 ) ;
  assign n14918 = n14916 ^ n13987 ^ n13933 ;
  assign n14919 = n7188 & ~n10956 ;
  assign n14920 = ( n7190 & ~n10959 ) | ( n7190 & n14919 ) | ( ~n10959 & n14919 ) ;
  assign n14921 = n14919 | n14920 ;
  assign n14922 = ( n7192 & n10951 ) | ( n7192 & n14919 ) | ( n10951 & n14919 ) ;
  assign n14923 = n14921 | n14922 ;
  assign n14924 = n7196 & n14425 ;
  assign n14925 = n14923 | n14924 ;
  assign n14926 = n14925 ^ x23 ^ 1'b0 ;
  assign n14927 = n14926 ^ n14918 ^ n14167 ;
  assign n14928 = ( n14167 & ~n14918 ) | ( n14167 & n14926 ) | ( ~n14918 & n14926 ) ;
  assign n14929 = n7188 & n10951 ;
  assign n14930 = ( n7190 & ~n10954 ) | ( n7190 & n14929 ) | ( ~n10954 & n14929 ) ;
  assign n14931 = n14929 | n14930 ;
  assign n14932 = ( n7192 & ~n10959 ) | ( n7192 & n14929 ) | ( ~n10959 & n14929 ) ;
  assign n14933 = n14931 | n14932 ;
  assign n14934 = n7196 & n14363 ;
  assign n14935 = n14933 | n14934 ;
  assign n14936 = n14935 ^ x23 ^ 1'b0 ;
  assign n14937 = n14936 ^ n14197 ^ n14166 ;
  assign n14938 = ( n14166 & n14197 ) | ( n14166 & n14936 ) | ( n14197 & n14936 ) ;
  assign n14939 = n7339 & ~n10968 ;
  assign n14940 = ( n7337 & ~n10967 ) | ( n7337 & n14939 ) | ( ~n10967 & n14939 ) ;
  assign n14941 = n14939 | n14940 ;
  assign n14942 = ( n7338 & ~n10956 ) | ( n7338 & n14939 ) | ( ~n10956 & n14939 ) ;
  assign n14943 = n14941 | n14942 ;
  assign n14944 = n7340 & ~n14478 ;
  assign n14945 = n14943 | n14944 ;
  assign n14946 = n14945 ^ x20 ^ 1'b0 ;
  assign n14947 = ( n14884 & n14937 ) | ( n14884 & n14946 ) | ( n14937 & n14946 ) ;
  assign n14948 = n14946 ^ n14937 ^ n14884 ;
  assign n14949 = n7339 & ~n10967 ;
  assign n14950 = ( n7337 & n10969 ) | ( n7337 & n14949 ) | ( n10969 & n14949 ) ;
  assign n14951 = n14949 | n14950 ;
  assign n14952 = ( n7338 & ~n10968 ) | ( n7338 & n14949 ) | ( ~n10968 & n14949 ) ;
  assign n14953 = n14951 | n14952 ;
  assign n14954 = n7340 & n14466 ;
  assign n14955 = n14953 | n14954 ;
  assign n14956 = n14955 ^ x20 ^ 1'b0 ;
  assign n14957 = n14956 ^ n14938 ^ n14927 ;
  assign n14958 = ( ~n14927 & n14938 ) | ( ~n14927 & n14956 ) | ( n14938 & n14956 ) ;
  assign n14959 = n7485 | n7487 ;
  assign n14960 = ( n7486 & n7493 ) | ( n7486 & n10969 ) | ( n7493 & n10969 ) ;
  assign n14961 = n7486 | n14959 ;
  assign n14962 = n14960 | n14961 ;
  assign n14963 = n14962 ^ x17 ^ 1'b0 ;
  assign n14964 = n14963 ^ n14948 ^ n14903 ;
  assign n14965 = ( n14903 & n14948 ) | ( n14903 & n14963 ) | ( n14948 & n14963 ) ;
  assign n14966 = ( n14905 & n14908 ) | ( n14905 & n14964 ) | ( n14908 & n14964 ) ;
  assign n14967 = n14957 ^ n14947 ^ n13644 ;
  assign n14968 = ( n13644 & n14947 ) | ( n13644 & ~n14957 ) | ( n14947 & ~n14957 ) ;
  assign n14969 = n14964 ^ n14908 ^ n14905 ;
  assign n14970 = n14967 ^ n14966 ^ n14965 ;
  assign n14971 = ( n14965 & n14966 ) | ( n14965 & ~n14967 ) | ( n14966 & ~n14967 ) ;
  assign n14972 = n7037 & ~n10959 ;
  assign n14973 = ( n7036 & ~n10954 ) | ( n7036 & n14972 ) | ( ~n10954 & n14972 ) ;
  assign n14974 = n14972 | n14973 ;
  assign n14975 = ( n7052 & n10957 ) | ( n7052 & n14972 ) | ( n10957 & n14972 ) ;
  assign n14976 = n14974 | n14975 ;
  assign n14977 = n7035 & n14327 ;
  assign n14978 = n14976 | n14977 ;
  assign n14979 = n14978 ^ x26 ^ 1'b0 ;
  assign n14980 = ( n14157 & n14917 ) | ( n14157 & n14979 ) | ( n14917 & n14979 ) ;
  assign n14981 = n14979 ^ n14917 ^ n14157 ;
  assign n14982 = n7188 & ~n10968 ;
  assign n14983 = ( n7190 & n10951 ) | ( n7190 & n14982 ) | ( n10951 & n14982 ) ;
  assign n14984 = n14982 | n14983 ;
  assign n14985 = ( n7192 & ~n10956 ) | ( n7192 & n14982 ) | ( ~n10956 & n14982 ) ;
  assign n14986 = n14984 | n14985 ;
  assign n14987 = n7196 & ~n14436 ;
  assign n14988 = n14986 | n14987 ;
  assign n14989 = n14988 ^ x23 ^ 1'b0 ;
  assign n14990 = ( n14928 & n14981 ) | ( n14928 & n14989 ) | ( n14981 & n14989 ) ;
  assign n14991 = n14989 ^ n14981 ^ n14928 ;
  assign n14992 = ( n7337 & n7339 ) | ( n7337 & n10969 ) | ( n7339 & n10969 ) ;
  assign n14993 = ( n7337 & n7338 ) | ( n7337 & ~n10967 ) | ( n7338 & ~n10967 ) ;
  assign n14994 = n7337 | n14992 ;
  assign n14995 = n14993 | n14994 ;
  assign n14996 = n7340 & n14468 ;
  assign n14997 = n14995 | n14996 ;
  assign n14998 = n14997 ^ x20 ^ 1'b0 ;
  assign n14999 = n14998 ^ n14991 ^ n14958 ;
  assign n15000 = ( n14958 & n14991 ) | ( n14958 & n14998 ) | ( n14991 & n14998 ) ;
  assign n15001 = n14999 ^ n14971 ^ n14968 ;
  assign n15002 = n7339 | n7340 ;
  assign n15003 = n7337 | n15002 ;
  assign n15004 = ( n14968 & n14971 ) | ( n14968 & n14999 ) | ( n14971 & n14999 ) ;
  assign n15005 = n7037 & n10951 ;
  assign n15006 = ( n7036 & ~n10959 ) | ( n7036 & n15005 ) | ( ~n10959 & n15005 ) ;
  assign n15007 = n15005 | n15006 ;
  assign n15008 = ( n7052 & ~n10954 ) | ( n7052 & n15005 ) | ( ~n10954 & n15005 ) ;
  assign n15009 = n7190 ^ n7189 ^ x23 ;
  assign n15010 = n15007 | n15008 ;
  assign n15011 = ( n7337 & n7338 ) | ( n7337 & n10969 ) | ( n7338 & n10969 ) ;
  assign n15012 = n15003 | n15011 ;
  assign n15013 = n7035 & n14363 ;
  assign n15014 = n15012 ^ x20 ^ 1'b0 ;
  assign n15015 = n15010 | n15013 ;
  assign n15016 = n15015 ^ x26 ^ 1'b0 ;
  assign n15017 = n15016 ^ n14156 ^ n14104 ;
  assign n15018 = ( ~n14104 & n14156 ) | ( ~n14104 & n15016 ) | ( n14156 & n15016 ) ;
  assign n15019 = n7188 & ~n10967 ;
  assign n15020 = ( n7190 & ~n10956 ) | ( n7190 & n15019 ) | ( ~n10956 & n15019 ) ;
  assign n15021 = n15019 | n15020 ;
  assign n15022 = ( n7192 & ~n10968 ) | ( n7192 & n15019 ) | ( ~n10968 & n15019 ) ;
  assign n15023 = n15021 | n15022 ;
  assign n15024 = n7196 & ~n14478 ;
  assign n15025 = n15023 | n15024 ;
  assign n15026 = n15025 ^ x23 ^ 1'b0 ;
  assign n15027 = ( n14980 & ~n15017 ) | ( n14980 & n15026 ) | ( ~n15017 & n15026 ) ;
  assign n15028 = n15026 ^ n15017 ^ n14980 ;
  assign n15029 = n15028 ^ n15014 ^ n14990 ;
  assign n15030 = ( n15000 & n15004 ) | ( n15000 & ~n15029 ) | ( n15004 & ~n15029 ) ;
  assign n15031 = ( n14990 & n15014 ) | ( n14990 & ~n15028 ) | ( n15014 & ~n15028 ) ;
  assign n15032 = n15029 ^ n15004 ^ n15000 ;
  assign n15033 = n7339 ^ n7338 ^ n7333 ;
  assign n15034 = n15033 ^ x20 ^ 1'b0 ;
  assign n15035 = n15034 ^ n6827 ^ n6342 ;
  assign n15036 = n15035 ^ n14224 ^ n14099 ;
  assign n15037 = ( n14099 & n14224 ) | ( n14099 & ~n15035 ) | ( n14224 & ~n15035 ) ;
  assign n15038 = n6901 & ~n10954 ;
  assign n15039 = ( n6906 & n10957 ) | ( n6906 & n15038 ) | ( n10957 & n15038 ) ;
  assign n15040 = n15038 | n15039 ;
  assign n15041 = ( n6907 & ~n10959 ) | ( n6907 & n15038 ) | ( ~n10959 & n15038 ) ;
  assign n15042 = n15040 | n15041 ;
  assign n15043 = n6918 & n14327 ;
  assign n15044 = n15042 | n15043 ;
  assign n15045 = n15044 ^ x29 ^ 1'b0 ;
  assign n15046 = n15045 ^ n15036 ^ n14109 ;
  assign n15047 = ( n14109 & ~n15036 ) | ( n14109 & n15045 ) | ( ~n15036 & n15045 ) ;
  assign n15048 = n6901 & n10957 ;
  assign n15049 = n6791 & n10957 ;
  assign n15050 = ( n6342 & n6827 ) | ( n6342 & n15034 ) | ( n6827 & n15034 ) ;
  assign n15051 = ( n6790 & n10965 ) | ( n6790 & n15049 ) | ( n10965 & n15049 ) ;
  assign n15052 = ( n6906 & n10965 ) | ( n6906 & n15048 ) | ( n10965 & n15048 ) ;
  assign n15053 = n15048 | n15052 ;
  assign n15054 = ( n6907 & ~n10954 ) | ( n6907 & n15048 ) | ( ~n10954 & n15048 ) ;
  assign n15055 = n15053 | n15054 ;
  assign n15056 = ( n6788 & ~n10954 ) | ( n6788 & n15049 ) | ( ~n10954 & n15049 ) ;
  assign n15057 = n15049 | n15056 ;
  assign n15058 = n15051 | n15057 ;
  assign n15059 = n7037 & ~n10956 ;
  assign n15060 = ( n7036 & n10951 ) | ( n7036 & n15059 ) | ( n10951 & n15059 ) ;
  assign n15061 = n15059 | n15060 ;
  assign n15062 = ( n7052 & ~n10959 ) | ( n7052 & n15059 ) | ( ~n10959 & n15059 ) ;
  assign n15063 = n15061 | n15062 ;
  assign n15064 = n6918 & ~n14281 ;
  assign n15065 = n15055 | n15064 ;
  assign n15066 = n7035 & n14425 ;
  assign n15067 = n15063 | n15066 ;
  assign n15068 = n15067 ^ x26 ^ 1'b0 ;
  assign n15069 = n15065 ^ x29 ^ 1'b0 ;
  assign n15070 = ( ~n14108 & n15068 ) | ( ~n14108 & n15069 ) | ( n15068 & n15069 ) ;
  assign n15071 = n6789 & ~n14281 ;
  assign n15072 = n15069 ^ n15068 ^ n14108 ;
  assign n15073 = n6788 & ~n10957 ;
  assign n15074 = n15058 | n15071 ;
  assign n15075 = n7188 & n10969 ;
  assign n15076 = ( n7190 & ~n10968 ) | ( n7190 & n15075 ) | ( ~n10968 & n15075 ) ;
  assign n15077 = n15075 | n15076 ;
  assign n15078 = ( n7192 & ~n10967 ) | ( n7192 & n15075 ) | ( ~n10967 & n15075 ) ;
  assign n15079 = n15077 | n15078 ;
  assign n15080 = n7196 & n14466 ;
  assign n15081 = n15079 | n15080 ;
  assign n15082 = n15081 ^ x23 ^ 1'b0 ;
  assign n15083 = ( n15018 & ~n15072 ) | ( n15018 & n15082 ) | ( ~n15072 & n15082 ) ;
  assign n15084 = n15082 ^ n15072 ^ n15018 ;
  assign n15085 = n6791 & ~n10954 ;
  assign n15086 = ( n6790 & n10957 ) | ( n6790 & n15085 ) | ( n10957 & n15085 ) ;
  assign n15087 = n15084 ^ n15034 ^ n15027 ;
  assign n15088 = ( n15027 & n15034 ) | ( n15027 & ~n15084 ) | ( n15034 & ~n15084 ) ;
  assign n15089 = ( n6788 & ~n10959 ) | ( n6788 & n15085 ) | ( ~n10959 & n15085 ) ;
  assign n15090 = ( n6788 & n14279 ) | ( n6788 & ~n15073 ) | ( n14279 & ~n15073 ) ;
  assign n15091 = n15090 ^ n15050 ^ n5160 ;
  assign n15092 = n6789 & ~n14327 ;
  assign n15093 = n15085 | n15089 ;
  assign n15094 = ( n6505 & n6780 ) | ( n6505 & ~n15009 ) | ( n6780 & ~n15009 ) ;
  assign n15095 = n15087 ^ n15031 ^ n15030 ;
  assign n15096 = n15086 | n15093 ;
  assign n15097 = n15009 ^ n6780 ^ n6505 ;
  assign n15098 = ( n15030 & n15031 ) | ( n15030 & ~n15087 ) | ( n15031 & ~n15087 ) ;
  assign n15099 = ( n6789 & ~n15092 ) | ( n6789 & n15096 ) | ( ~n15092 & n15096 ) ;
  assign n15100 = ( n5160 & n15050 ) | ( n5160 & ~n15090 ) | ( n15050 & ~n15090 ) ;
  assign n15101 = ( ~n5160 & n6505 ) | ( ~n5160 & n15100 ) | ( n6505 & n15100 ) ;
  assign n15102 = n15101 ^ n15099 ^ n15097 ;
  assign n15103 = n15100 ^ n6505 ^ n5160 ;
  assign n15104 = ( n15097 & ~n15099 ) | ( n15097 & n15101 ) | ( ~n15099 & n15101 ) ;
  assign n15105 = n6901 & n10951 ;
  assign n15106 = ( n6906 & ~n10959 ) | ( n6906 & n15105 ) | ( ~n10959 & n15105 ) ;
  assign n15107 = n15105 | n15106 ;
  assign n15108 = ( n6907 & ~n10956 ) | ( n6907 & n15105 ) | ( ~n10956 & n15105 ) ;
  assign n15109 = n15107 | n15108 ;
  assign n15110 = ( n6918 & n14425 ) | ( n6918 & n15109 ) | ( n14425 & n15109 ) ;
  assign n15111 = n15109 | n15110 ;
  assign n15112 = n15111 ^ x29 ^ 1'b0 ;
  assign n15113 = ( n15074 & n15103 ) | ( n15074 & n15112 ) | ( n15103 & n15112 ) ;
  assign n15114 = n15112 ^ n15103 ^ n15074 ;
  assign n15115 = n6789 & n14363 ;
  assign n15116 = ( n6791 & ~n10959 ) | ( n6791 & n15115 ) | ( ~n10959 & n15115 ) ;
  assign n15117 = n15115 | n15116 ;
  assign n15118 = ( n6790 & ~n10954 ) | ( n6790 & n15115 ) | ( ~n10954 & n15115 ) ;
  assign n15119 = n15117 | n15118 ;
  assign n15120 = n6901 & ~n10959 ;
  assign n15121 = ( n6906 & ~n10954 ) | ( n6906 & n15120 ) | ( ~n10954 & n15120 ) ;
  assign n15122 = n15120 | n15121 ;
  assign n15123 = ( n6907 & n10951 ) | ( n6907 & n15120 ) | ( n10951 & n15120 ) ;
  assign n15124 = n15122 | n15123 ;
  assign n15125 = n7037 & ~n10967 ;
  assign n15126 = n6789 & ~n14425 ;
  assign n15127 = ( n6918 & n14363 ) | ( n6918 & n15124 ) | ( n14363 & n15124 ) ;
  assign n15128 = n15124 | n15127 ;
  assign n15129 = n15128 ^ x29 ^ 1'b0 ;
  assign n15130 = ( n7036 & ~n10968 ) | ( n7036 & n15125 ) | ( ~n10968 & n15125 ) ;
  assign n15131 = n15125 | n15130 ;
  assign n15132 = ( n7052 & ~n10956 ) | ( n7052 & n15125 ) | ( ~n10956 & n15125 ) ;
  assign n15133 = n15131 | n15132 ;
  assign n15134 = ( n15037 & n15091 ) | ( n15037 & n15129 ) | ( n15091 & n15129 ) ;
  assign n15135 = n15129 ^ n15091 ^ n15037 ;
  assign n15136 = n6791 & n10951 ;
  assign n15137 = ( n6788 & ~n10956 ) | ( n6788 & n15136 ) | ( ~n10956 & n15136 ) ;
  assign n15138 = n15136 | n15137 ;
  assign n15139 = ( n6790 & ~n10959 ) | ( n6790 & n15136 ) | ( ~n10959 & n15136 ) ;
  assign n15140 = n7037 & n10969 ;
  assign n15141 = n15138 | n15139 ;
  assign n15142 = ( n7036 & ~n10967 ) | ( n7036 & n15140 ) | ( ~n10967 & n15140 ) ;
  assign n15143 = n15140 | n15142 ;
  assign n15144 = ( n7052 & ~n10968 ) | ( n7052 & n15140 ) | ( ~n10968 & n15140 ) ;
  assign n15145 = n15143 | n15144 ;
  assign n15146 = n7035 & n14466 ;
  assign n15147 = n15145 | n15146 ;
  assign n15148 = n7035 & ~n14478 ;
  assign n15149 = n15133 | n15148 ;
  assign n15150 = n15149 ^ x26 ^ 1'b0 ;
  assign n15151 = n15150 ^ n15135 ^ n15047 ;
  assign n15152 = ( n15047 & n15135 ) | ( n15047 & n15150 ) | ( n15135 & n15150 ) ;
  assign n15153 = n15147 ^ x26 ^ 1'b0 ;
  assign n15154 = n15153 ^ n15134 ^ n15114 ;
  assign n15155 = ( n15009 & n15152 ) | ( n15009 & n15154 ) | ( n15152 & n15154 ) ;
  assign n15156 = n15154 ^ n15152 ^ n15009 ;
  assign n15157 = ( n15114 & n15134 ) | ( n15114 & n15153 ) | ( n15134 & n15153 ) ;
  assign n15158 = ( n6789 & ~n15126 ) | ( n6789 & n15141 ) | ( ~n15126 & n15141 ) ;
  assign n15159 = n7037 & ~n10968 ;
  assign n15160 = ( n7036 & ~n10956 ) | ( n7036 & n15159 ) | ( ~n10956 & n15159 ) ;
  assign n15161 = n15159 | n15160 ;
  assign n15162 = ( n7052 & n10951 ) | ( n7052 & n15159 ) | ( n10951 & n15159 ) ;
  assign n15163 = n15161 | n15162 ;
  assign n15164 = n7035 & ~n14436 ;
  assign n15165 = n15163 | n15164 ;
  assign n15166 = n15165 ^ x26 ^ 1'b0 ;
  assign n15167 = ( ~n15046 & n15070 ) | ( ~n15046 & n15166 ) | ( n15070 & n15166 ) ;
  assign n15168 = n15166 ^ n15070 ^ n15046 ;
  assign n15169 = n6791 & ~n10956 ;
  assign n15170 = ( n6788 & ~n10968 ) | ( n6788 & n15169 ) | ( ~n10968 & n15169 ) ;
  assign n15171 = n15169 | n15170 ;
  assign n15172 = ( n6790 & n10951 ) | ( n6790 & n15169 ) | ( n10951 & n15169 ) ;
  assign n15173 = n15171 | n15172 ;
  assign n15174 = n15158 ^ n6690 ^ n6440 ;
  assign n15175 = ( n6440 & n6690 ) | ( n6440 & n15158 ) | ( n6690 & n15158 ) ;
  assign n15176 = n7034 ^ x26 ^ 1'b0 ;
  assign n15177 = n6788 & ~n10951 ;
  assign n15178 = ( n6788 & n15119 ) | ( n6788 & ~n15177 ) | ( n15119 & ~n15177 ) ;
  assign n15179 = n6789 & ~n14436 ;
  assign n15180 = n15173 | n15179 ;
  assign n15181 = n6901 & ~n10956 ;
  assign n15182 = ( n6906 & n10951 ) | ( n6906 & n15181 ) | ( n10951 & n15181 ) ;
  assign n15183 = n6918 & ~n14436 ;
  assign n15184 = n15181 | n15182 ;
  assign n15185 = ( n6907 & ~n10968 ) | ( n6907 & n15181 ) | ( ~n10968 & n15181 ) ;
  assign n15186 = n15184 | n15185 ;
  assign n15187 = n7188 | n7196 ;
  assign n15188 = n15183 | n15186 ;
  assign n15189 = n15188 ^ x29 ^ 1'b0 ;
  assign n15190 = n15189 ^ n15113 ^ n15102 ;
  assign n15191 = ( n15102 & n15113 ) | ( n15102 & n15189 ) | ( n15113 & n15189 ) ;
  assign n15192 = ( n7188 & n7190 ) | ( n7188 & n10969 ) | ( n7190 & n10969 ) ;
  assign n15193 = ( n6573 & n6690 ) | ( n6573 & n15176 ) | ( n6690 & n15176 ) ;
  assign n15194 = n7192 | n15192 ;
  assign n15195 = n15187 | n15194 ;
  assign n15196 = n15176 ^ n6690 ^ n6573 ;
  assign n15197 = n15196 ^ n15180 ^ n15175 ;
  assign n15198 = ( n15175 & n15180 ) | ( n15175 & ~n15196 ) | ( n15180 & ~n15196 ) ;
  assign n15199 = n15094 ^ n6690 ^ 1'b0 ;
  assign n15200 = ( n7188 & n7192 ) | ( n7188 & n10969 ) | ( n7192 & n10969 ) ;
  assign n15201 = n15199 ^ n15178 ^ 1'b0 ;
  assign n15202 = ( n6690 & n15094 ) | ( n6690 & n15178 ) | ( n15094 & n15178 ) ;
  assign n15203 = n7196 & n14468 ;
  assign n15204 = ( n7188 & n7190 ) | ( n7188 & ~n10967 ) | ( n7190 & ~n10967 ) ;
  assign n15205 = n7188 | n15204 ;
  assign n15206 = n15200 | n15205 ;
  assign n15207 = n15203 | n15206 ;
  assign n15208 = n15195 ^ x23 ^ 1'b0 ;
  assign n15209 = n15207 ^ x23 ^ 1'b0 ;
  assign n15210 = n15209 ^ n15168 ^ n15083 ;
  assign n15211 = ( n15151 & n15167 ) | ( n15151 & n15208 ) | ( n15167 & n15208 ) ;
  assign n15212 = ( n15083 & ~n15168 ) | ( n15083 & n15209 ) | ( ~n15168 & n15209 ) ;
  assign n15213 = ( n15088 & n15098 ) | ( n15088 & ~n15210 ) | ( n15098 & ~n15210 ) ;
  assign n15214 = n15208 ^ n15167 ^ n15151 ;
  assign n15215 = ( n15212 & n15213 ) | ( n15212 & n15214 ) | ( n15213 & n15214 ) ;
  assign n15216 = n15210 ^ n15098 ^ n15088 ;
  assign n15217 = ( n15156 & n15211 ) | ( n15156 & n15215 ) | ( n15211 & n15215 ) ;
  assign n15218 = n15214 ^ n15213 ^ n15212 ;
  assign n15219 = n15215 ^ n15211 ^ n15156 ;
  assign n15220 = n6901 & ~n10968 ;
  assign n15221 = ( n6906 & ~n10956 ) | ( n6906 & n15220 ) | ( ~n10956 & n15220 ) ;
  assign n15222 = n15220 | n15221 ;
  assign n15223 = ( n6907 & ~n10967 ) | ( n6907 & n15220 ) | ( ~n10967 & n15220 ) ;
  assign n15224 = n15222 | n15223 ;
  assign n15225 = n14478 & ~n15224 ;
  assign n15226 = ( n6918 & n15224 ) | ( n6918 & ~n15225 ) | ( n15224 & ~n15225 ) ;
  assign n15227 = n15226 ^ x29 ^ 1'b0 ;
  assign n15228 = ( ~n15104 & n15201 ) | ( ~n15104 & n15227 ) | ( n15201 & n15227 ) ;
  assign n15229 = n15227 ^ n15201 ^ n15104 ;
  assign n15230 = ( n7036 & n7037 ) | ( n7036 & n10969 ) | ( n7037 & n10969 ) ;
  assign n15231 = n7037 | n15230 ;
  assign n15232 = ( n7037 & n7052 ) | ( n7037 & ~n10967 ) | ( n7052 & ~n10967 ) ;
  assign n15233 = n15231 | n15232 ;
  assign n15234 = n7035 & n14468 ;
  assign n15235 = n15233 | n15234 ;
  assign n15236 = n15235 ^ x26 ^ 1'b0 ;
  assign n15237 = ( n15157 & n15190 ) | ( n15157 & n15236 ) | ( n15190 & n15236 ) ;
  assign n15238 = n15236 ^ n15190 ^ n15157 ;
  assign n15239 = n15238 ^ n15217 ^ n15155 ;
  assign n15240 = n7036 | n7037 ;
  assign n15241 = n7035 | n15240 ;
  assign n15242 = ( n15155 & n15217 ) | ( n15155 & n15238 ) | ( n15217 & n15238 ) ;
  assign n15243 = ( n7035 & n7052 ) | ( n7035 & n10969 ) | ( n7052 & n10969 ) ;
  assign n15244 = n15241 | n15243 ;
  assign n15245 = n15244 ^ x26 ^ 1'b0 ;
  assign n15246 = n15245 ^ n15229 ^ n15191 ;
  assign n15247 = ( n15237 & n15242 ) | ( n15237 & ~n15246 ) | ( n15242 & ~n15246 ) ;
  assign n15248 = n15246 ^ n15242 ^ n15237 ;
  assign n15249 = ( n6901 & n6918 ) | ( n6901 & n14468 ) | ( n6918 & n14468 ) ;
  assign n15250 = ( n6901 & n6906 ) | ( n6901 & ~n10967 ) | ( n6906 & ~n10967 ) ;
  assign n15251 = n15249 | n15250 ;
  assign n15252 = ( n15174 & n15202 ) | ( n15174 & n15228 ) | ( n15202 & n15228 ) ;
  assign n15253 = n15228 ^ n15202 ^ n15174 ;
  assign n15254 = n6901 | n6907 ;
  assign n15255 = n15251 | n15254 ;
  assign n15256 = n6901 & ~n10967 ;
  assign n15257 = ( n6906 & ~n10968 ) | ( n6906 & n15256 ) | ( ~n10968 & n15256 ) ;
  assign n15258 = n15256 | n15257 ;
  assign n15259 = ( n6907 & n10969 ) | ( n6907 & n15256 ) | ( n10969 & n15256 ) ;
  assign n15260 = n15255 ^ x29 ^ 1'b0 ;
  assign n15261 = n15258 | n15259 ;
  assign n15262 = n15260 ^ n15252 ^ n15197 ;
  assign n15263 = ( ~n15197 & n15252 ) | ( ~n15197 & n15260 ) | ( n15252 & n15260 ) ;
  assign n15264 = n6789 & ~n14478 ;
  assign n15265 = ~n6918 & n14466 ;
  assign n15266 = ( n14466 & n15261 ) | ( n14466 & ~n15265 ) | ( n15261 & ~n15265 ) ;
  assign n15267 = n15266 ^ x29 ^ 1'b0 ;
  assign n15268 = n15267 ^ n15253 ^ n15176 ;
  assign n15269 = ( n15191 & ~n15229 ) | ( n15191 & n15245 ) | ( ~n15229 & n15245 ) ;
  assign n15270 = ( n15247 & n15268 ) | ( n15247 & n15269 ) | ( n15268 & n15269 ) ;
  assign n15271 = n15269 ^ n15268 ^ n15247 ;
  assign n15272 = ( n15176 & n15253 ) | ( n15176 & n15267 ) | ( n15253 & n15267 ) ;
  assign n15273 = ( ~n15262 & n15270 ) | ( ~n15262 & n15272 ) | ( n15270 & n15272 ) ;
  assign n15274 = n15272 ^ n15262 ^ 1'b0 ;
  assign n15275 = n15274 ^ n15270 ^ 1'b0 ;
  assign n15276 = ( n6788 & n6791 ) | ( n6788 & n10969 ) | ( n6791 & n10969 ) ;
  assign n15277 = ( n6788 & n6789 ) | ( n6788 & n14468 ) | ( n6789 & n14468 ) ;
  assign n15278 = n15276 | n15277 ;
  assign n15279 = n6791 & ~n10967 ;
  assign n15280 = ( n6788 & n10969 ) | ( n6788 & n15279 ) | ( n10969 & n15279 ) ;
  assign n15281 = n15279 | n15280 ;
  assign n15282 = ( n6790 & ~n10968 ) | ( n6790 & n15279 ) | ( ~n10968 & n15279 ) ;
  assign n15283 = n6791 & ~n10968 ;
  assign n15284 = ( n6788 & ~n10967 ) | ( n6788 & n15283 ) | ( ~n10967 & n15283 ) ;
  assign n15285 = n15283 | n15284 ;
  assign n15286 = ( n6790 & ~n10956 ) | ( n6790 & n15283 ) | ( ~n10956 & n15283 ) ;
  assign n15287 = n15285 | n15286 ;
  assign n15288 = n15193 ^ n6575 ^ 1'b0 ;
  assign n15289 = n6788 | n6790 ;
  assign n15290 = n15278 | n15289 ;
  assign n15291 = n6903 ^ x29 ^ 1'b0 ;
  assign n15292 = n15264 | n15287 ;
  assign n15293 = n15292 ^ n15288 ^ 1'b0 ;
  assign n15294 = n15293 ^ n15291 ^ n15198 ;
  assign n15295 = n15281 | n15282 ;
  assign n15296 = n15294 ^ n15263 ^ 1'b0 ;
  assign n15297 = ( n15263 & n15273 ) | ( n15263 & n15294 ) | ( n15273 & n15294 ) ;
  assign n15298 = n6791 ^ n6790 ^ n6787 ;
  assign n15299 = ( n15198 & n15291 ) | ( n15198 & n15293 ) | ( n15291 & n15293 ) ;
  assign n15300 = ( n6237 & n9904 ) | ( n6237 & ~n15291 ) | ( n9904 & ~n15291 ) ;
  assign n15301 = ( n6575 & n15193 ) | ( n6575 & ~n15292 ) | ( n15193 & ~n15292 ) ;
  assign n15302 = n6789 & ~n14466 ;
  assign n15303 = ( n6789 & n15295 ) | ( n6789 & ~n15302 ) | ( n15295 & ~n15302 ) ;
  assign n15304 = n15301 ^ n9904 ^ n6575 ;
  assign n15305 = n15304 ^ n15303 ^ n15291 ;
  assign n15306 = n15305 ^ n15299 ^ 1'b0 ;
  assign n15307 = ( n15297 & n15299 ) | ( n15297 & n15305 ) | ( n15299 & n15305 ) ;
  assign n15308 = n15306 ^ n15297 ^ 1'b0 ;
  assign n15309 = n15291 ^ n9904 ^ n6237 ;
  assign n15310 = n15300 ^ n15298 ^ n6035 ;
  assign n15311 = ( ~n6575 & n9904 ) | ( ~n6575 & n15301 ) | ( n9904 & n15301 ) ;
  assign n15312 = n15296 ^ n15273 ^ 1'b0 ;
  assign n15313 = ( ~n15290 & n15309 ) | ( ~n15290 & n15311 ) | ( n15309 & n15311 ) ;
  assign n15314 = n15313 ^ n15310 ^ 1'b0 ;
  assign n15315 = n15311 ^ n15309 ^ n15290 ;
  assign n15316 = ( n15291 & n15303 ) | ( n15291 & n15304 ) | ( n15303 & n15304 ) ;
  assign n15317 = n15316 ^ n15315 ^ 1'b0 ;
  assign n15318 = ( n15307 & n15315 ) | ( n15307 & n15316 ) | ( n15315 & n15316 ) ;
  assign n15319 = n15317 ^ n15307 ^ 1'b0 ;
  assign n15320 = n15318 ^ n15314 ^ 1'b0 ;
  assign n15321 = ( n15310 & ~n15313 ) | ( n15310 & n15318 ) | ( ~n15313 & n15318 ) ;
  assign n15322 = n15321 ^ n15298 ^ 1'b0 ;
  assign n15323 = n6791 & ~n14378 ;
  assign n15324 = ( n6788 & n14418 ) | ( n6788 & n15323 ) | ( n14418 & n15323 ) ;
  assign n15325 = ( n6790 & ~n14324 ) | ( n6790 & n15323 ) | ( ~n14324 & n15323 ) ;
  assign n15326 = n14378 ^ n14324 ^ 1'b0 ;
  assign n15327 = ( x2 & ~n8113 ) | ( x2 & n14324 ) | ( ~n8113 & n14324 ) ;
  assign n15328 = n15323 | n15324 ;
  assign n15329 = n15325 | n15328 ;
  assign n15330 = x2 & n15327 ;
  assign n15331 = n6789 & n15326 ;
  assign n15332 = ( n6788 & ~n14378 ) | ( n6788 & n15331 ) | ( ~n14378 & n15331 ) ;
  assign n15333 = ( n14324 & n14378 ) | ( n14324 & ~n14418 ) | ( n14378 & ~n14418 ) ;
  assign n15334 = ( n6791 & ~n14324 ) | ( n6791 & n15331 ) | ( ~n14324 & n15331 ) ;
  assign n15335 = n15331 | n15334 ;
  assign n15336 = ( x2 & ~n8090 ) | ( x2 & n14378 ) | ( ~n8090 & n14378 ) ;
  assign n15337 = n15332 | n15335 ;
  assign n15338 = n15337 ^ n6561 ^ 1'b0 ;
  assign n15339 = ~n6561 & n15337 ;
  assign n15340 = n15330 & n15336 ;
  assign n15341 = n14324 & ~n14378 ;
  assign n15342 = n15341 ^ n14418 ^ 1'b0 ;
  assign n15343 = n6789 & ~n15342 ;
  assign n15344 = ( n6789 & n15329 ) | ( n6789 & ~n15343 ) | ( n15329 & ~n15343 ) ;
  assign n15345 = n15344 ^ n15339 ^ n6682 ;
  assign n15346 = ( ~n6682 & n15339 ) | ( ~n6682 & n15344 ) | ( n15339 & n15344 ) ;
  assign n15347 = n8086 & ~n14324 ;
  assign n15348 = n7483 & ~n14324 ;
  assign n15349 = n7187 & ~n14324 ;
  assign n15350 = n8120 & n15342 ;
  assign n15351 = n7827 & ~n14324 ;
  assign n15352 = n14378 | n15333 ;
  assign n15353 = n8025 & ~n14324 ;
  assign n15354 = n7333 & ~n14324 ;
  assign n15355 = n7927 & ~n14324 ;
  assign n15356 = n8120 & n15326 ;
  assign n15357 = ( n15340 & ~n15350 ) | ( n15340 & n15356 ) | ( ~n15350 & n15356 ) ;
  assign n15358 = ~n15356 & n15357 ;
  assign n15359 = ( n8088 & ~n14378 ) | ( n8088 & n15347 ) | ( ~n14378 & n15347 ) ;
  assign n15360 = n15347 | n15359 ;
  assign n15361 = ( n8090 & n14418 ) | ( n8090 & n15347 ) | ( n14418 & n15347 ) ;
  assign n15362 = n15360 | n15361 ;
  assign n15363 = ( ~n14418 & n14461 ) | ( ~n14418 & n15352 ) | ( n14461 & n15352 ) ;
  assign n15364 = ( x2 & n15350 ) | ( x2 & n15362 ) | ( n15350 & n15362 ) ;
  assign n15365 = x0 & ~n14324 ;
  assign n15366 = ( n15358 & n15364 ) | ( n15358 & ~n15365 ) | ( n15364 & ~n15365 ) ;
  assign n15367 = ~n15364 & n15366 ;
  assign n15368 = n15352 ^ n14461 ^ n14418 ;
  assign n15369 = n6789 & n15368 ;
  assign n15370 = ( n6791 & n14418 ) | ( n6791 & n15369 ) | ( n14418 & n15369 ) ;
  assign n15371 = n15369 | n15370 ;
  assign n15372 = ( n6790 & ~n14378 ) | ( n6790 & n15369 ) | ( ~n14378 & n15369 ) ;
  assign n15373 = n15371 | n15372 ;
  assign n15374 = n6788 & ~n14461 ;
  assign n15375 = n15373 | n15374 ;
  assign n15376 = n15375 ^ n15346 ^ n6630 ;
  assign n15377 = ( n6630 & n15346 ) | ( n6630 & n15375 ) | ( n15346 & n15375 ) ;
  assign n15378 = n8086 & ~n14378 ;
  assign n15379 = ( n8088 & n14418 ) | ( n8088 & n15378 ) | ( n14418 & n15378 ) ;
  assign n15380 = n15378 | n15379 ;
  assign n15381 = n7030 & ~n14324 ;
  assign n15382 = ( n8090 & ~n14461 ) | ( n8090 & n15378 ) | ( ~n14461 & n15378 ) ;
  assign n15383 = n15380 | n15382 ;
  assign n15384 = ~n8089 & n15368 ;
  assign n15385 = ( n15368 & n15383 ) | ( n15368 & ~n15384 ) | ( n15383 & ~n15384 ) ;
  assign n15386 = n15385 ^ x2 ^ 1'b0 ;
  assign n15387 = ( n15353 & n15367 ) | ( n15353 & n15386 ) | ( n15367 & n15386 ) ;
  assign n15388 = n6787 & ~n14324 ;
  assign n15389 = x5 & ~n15353 ;
  assign n15390 = n7663 & ~n14324 ;
  assign n15391 = n6898 & ~n14324 ;
  assign n15392 = n8034 & n15326 ;
  assign n15393 = n8086 & n14418 ;
  assign n15394 = ( n8033 & ~n14378 ) | ( n8033 & n15392 ) | ( ~n14378 & n15392 ) ;
  assign n15395 = ( n8090 & ~n14549 ) | ( n8090 & n15393 ) | ( ~n14549 & n15393 ) ;
  assign n15396 = ( n8029 & ~n14324 ) | ( n8029 & n15392 ) | ( ~n14324 & n15392 ) ;
  assign n15397 = n15392 | n15396 ;
  assign n15398 = n15394 | n15397 ;
  assign n15399 = ( n14461 & n14549 ) | ( n14461 & n15363 ) | ( n14549 & n15363 ) ;
  assign n15400 = ( n8088 & ~n14461 ) | ( n8088 & n15393 ) | ( ~n14461 & n15393 ) ;
  assign n15401 = n15393 | n15400 ;
  assign n15402 = n15395 | n15401 ;
  assign n15403 = n15398 ^ x5 ^ 1'b0 ;
  assign n15404 = n15389 & n15403 ;
  assign n15405 = n15363 ^ n14549 ^ n14461 ;
  assign n15406 = n15403 ^ n15389 ^ 1'b0 ;
  assign n15407 = ~n15402 & n15405 ;
  assign n15408 = ( n8089 & n15402 ) | ( n8089 & ~n15407 ) | ( n15402 & ~n15407 ) ;
  assign n15409 = n15408 ^ x2 ^ 1'b0 ;
  assign n15410 = ( n14549 & ~n14559 ) | ( n14549 & n15399 ) | ( ~n14559 & n15399 ) ;
  assign n15411 = ( n15387 & n15406 ) | ( n15387 & n15409 ) | ( n15406 & n15409 ) ;
  assign n15412 = n6789 & ~n15405 ;
  assign n15413 = ( n6791 & ~n14461 ) | ( n6791 & n15412 ) | ( ~n14461 & n15412 ) ;
  assign n15414 = n15412 | n15413 ;
  assign n15415 = ( n6790 & n14418 ) | ( n6790 & n15412 ) | ( n14418 & n15412 ) ;
  assign n15416 = n15414 | n15415 ;
  assign n15417 = n15399 ^ n14559 ^ n14549 ;
  assign n15418 = n6789 & n15417 ;
  assign n15419 = ( n6791 & ~n14549 ) | ( n6791 & n15418 ) | ( ~n14549 & n15418 ) ;
  assign n15420 = n15418 | n15419 ;
  assign n15421 = ( n6790 & ~n14461 ) | ( n6790 & n15418 ) | ( ~n14461 & n15418 ) ;
  assign n15422 = n15420 | n15421 ;
  assign n15423 = n6788 & ~n14549 ;
  assign n15424 = n15416 | n15423 ;
  assign n15425 = ( ~n6579 & n15377 ) | ( ~n6579 & n15424 ) | ( n15377 & n15424 ) ;
  assign n15426 = n15424 ^ n15377 ^ n6579 ;
  assign n15427 = n8029 & ~n14378 ;
  assign n15428 = ( n8037 & ~n14324 ) | ( n8037 & n15427 ) | ( ~n14324 & n15427 ) ;
  assign n15429 = n15427 | n15428 ;
  assign n15430 = ( n8033 & n14418 ) | ( n8033 & n15429 ) | ( n14418 & n15429 ) ;
  assign n15431 = n15429 | n15430 ;
  assign n15432 = ( n8034 & n15342 ) | ( n8034 & n15429 ) | ( n15342 & n15429 ) ;
  assign n15433 = n15431 | n15432 ;
  assign n15434 = n6788 & ~n14559 ;
  assign n15435 = ( n6788 & n15422 ) | ( n6788 & ~n15434 ) | ( n15422 & ~n15434 ) ;
  assign n15436 = n15435 ^ n15425 ^ n6443 ;
  assign n15437 = n15433 ^ x5 ^ 1'b0 ;
  assign n15438 = ( ~n6443 & n15425 ) | ( ~n6443 & n15435 ) | ( n15425 & n15435 ) ;
  assign n15439 = n8086 & ~n14461 ;
  assign n15440 = ( n8088 & ~n14549 ) | ( n8088 & n15439 ) | ( ~n14549 & n15439 ) ;
  assign n15441 = n15439 | n15440 ;
  assign n15442 = ( n8090 & n14559 ) | ( n8090 & n15439 ) | ( n14559 & n15439 ) ;
  assign n15443 = n15441 | n15442 ;
  assign n15444 = ~n8089 & n15417 ;
  assign n15445 = ( n15417 & n15443 ) | ( n15417 & ~n15444 ) | ( n15443 & ~n15444 ) ;
  assign n15446 = n15445 ^ x2 ^ 1'b0 ;
  assign n15447 = n15404 & n15437 ;
  assign n15448 = n15437 ^ n15404 ^ 1'b0 ;
  assign n15449 = ( n15411 & n15446 ) | ( n15411 & n15448 ) | ( n15446 & n15448 ) ;
  assign n15450 = ( n14559 & n14569 ) | ( n14559 & ~n15410 ) | ( n14569 & ~n15410 ) ;
  assign n15451 = n8029 & n14418 ;
  assign n15452 = n15410 ^ n14569 ^ n14559 ;
  assign n15453 = n6789 & ~n15452 ;
  assign n15454 = ( n8037 & ~n14378 ) | ( n8037 & n15451 ) | ( ~n14378 & n15451 ) ;
  assign n15455 = ( n6791 & n14559 ) | ( n6791 & n15453 ) | ( n14559 & n15453 ) ;
  assign n15456 = n15453 | n15455 ;
  assign n15457 = ( n6790 & ~n14549 ) | ( n6790 & n15453 ) | ( ~n14549 & n15453 ) ;
  assign n15458 = n15456 | n15457 ;
  assign n15459 = n8086 & ~n14549 ;
  assign n15460 = n15451 | n15454 ;
  assign n15461 = ( n8033 & ~n14461 ) | ( n8033 & n15451 ) | ( ~n14461 & n15451 ) ;
  assign n15462 = n15460 | n15461 ;
  assign n15463 = ( n8088 & n14559 ) | ( n8088 & n15459 ) | ( n14559 & n15459 ) ;
  assign n15464 = n15459 | n15463 ;
  assign n15465 = ( n8090 & n14569 ) | ( n8090 & n15459 ) | ( n14569 & n15459 ) ;
  assign n15466 = n15464 | n15465 ;
  assign n15467 = n15452 & ~n15466 ;
  assign n15468 = ( n8089 & n15466 ) | ( n8089 & ~n15467 ) | ( n15466 & ~n15467 ) ;
  assign n15469 = n15468 ^ x2 ^ 1'b0 ;
  assign n15470 = n8034 & n15368 ;
  assign n15471 = n15462 | n15470 ;
  assign n15472 = n15471 ^ x5 ^ 1'b0 ;
  assign n15473 = n15472 ^ n15447 ^ n15355 ;
  assign n15474 = ( n15449 & n15469 ) | ( n15449 & n15473 ) | ( n15469 & n15473 ) ;
  assign n15475 = n15450 ^ n14578 ^ n14569 ;
  assign n15476 = n6788 & ~n14569 ;
  assign n15477 = ( n6788 & n15458 ) | ( n6788 & ~n15476 ) | ( n15458 & ~n15476 ) ;
  assign n15478 = ( ~n6578 & n15438 ) | ( ~n6578 & n15477 ) | ( n15438 & n15477 ) ;
  assign n15479 = ( n14569 & n14578 ) | ( n14569 & n15450 ) | ( n14578 & n15450 ) ;
  assign n15480 = n15477 ^ n15438 ^ n6578 ;
  assign n15481 = n6789 & n15475 ;
  assign n15482 = ( n6791 & n14569 ) | ( n6791 & n15481 ) | ( n14569 & n15481 ) ;
  assign n15483 = n15481 | n15482 ;
  assign n15484 = ( n6790 & n14559 ) | ( n6790 & n15481 ) | ( n14559 & n15481 ) ;
  assign n15485 = n15483 | n15484 ;
  assign n15486 = n7932 & ~n14324 ;
  assign n15487 = ( n15355 & n15447 ) | ( n15355 & n15472 ) | ( n15447 & n15472 ) ;
  assign n15488 = n6788 & ~n14578 ;
  assign n15489 = ( n6788 & n15485 ) | ( n6788 & ~n15488 ) | ( n15485 & ~n15488 ) ;
  assign n15490 = ( n6722 & n15478 ) | ( n6722 & n15489 ) | ( n15478 & n15489 ) ;
  assign n15491 = n15489 ^ n15478 ^ n6722 ;
  assign n15492 = ( n7930 & n15326 ) | ( n7930 & n15486 ) | ( n15326 & n15486 ) ;
  assign n15493 = n15486 | n15492 ;
  assign n15494 = n8029 & ~n14461 ;
  assign n15495 = ( n7929 & ~n14378 ) | ( n7929 & n15486 ) | ( ~n14378 & n15486 ) ;
  assign n15496 = n15493 | n15495 ;
  assign n15497 = n15496 ^ x8 ^ 1'b0 ;
  assign n15498 = ( n8037 & n14418 ) | ( n8037 & n15494 ) | ( n14418 & n15494 ) ;
  assign n15499 = n15494 | n15498 ;
  assign n15500 = x8 & ~n15355 ;
  assign n15501 = ( n8033 & ~n14549 ) | ( n8033 & n15494 ) | ( ~n14549 & n15494 ) ;
  assign n15502 = n15499 | n15501 ;
  assign n15503 = n15500 ^ n15497 ^ 1'b0 ;
  assign n15504 = n15497 & n15500 ;
  assign n15505 = n8034 & ~n15405 ;
  assign n15506 = n15502 & ~n15505 ;
  assign n15507 = n15506 ^ n15505 ^ x5 ;
  assign n15508 = ( n15487 & n15503 ) | ( n15487 & n15507 ) | ( n15503 & n15507 ) ;
  assign n15509 = n15507 ^ n15503 ^ n15487 ;
  assign n15510 = n8086 & n14559 ;
  assign n15511 = ( n8088 & n14569 ) | ( n8088 & n15510 ) | ( n14569 & n15510 ) ;
  assign n15512 = n15510 | n15511 ;
  assign n15513 = ( n8090 & n14578 ) | ( n8090 & n15510 ) | ( n14578 & n15510 ) ;
  assign n15514 = n15512 | n15513 ;
  assign n15515 = ~n8089 & n15475 ;
  assign n15516 = ( n15475 & n15514 ) | ( n15475 & ~n15515 ) | ( n15514 & ~n15515 ) ;
  assign n15517 = n15516 ^ x2 ^ 1'b0 ;
  assign n15518 = ( n15474 & n15509 ) | ( n15474 & n15517 ) | ( n15509 & n15517 ) ;
  assign n15519 = n7932 & ~n14378 ;
  assign n15520 = n8029 & ~n14549 ;
  assign n15521 = ( n7943 & ~n14324 ) | ( n7943 & n15519 ) | ( ~n14324 & n15519 ) ;
  assign n15522 = ( n8037 & ~n14461 ) | ( n8037 & n15520 ) | ( ~n14461 & n15520 ) ;
  assign n15523 = n15520 | n15522 ;
  assign n15524 = ( n8033 & n14559 ) | ( n8033 & n15520 ) | ( n14559 & n15520 ) ;
  assign n15525 = n15519 | n15521 ;
  assign n15526 = ( n7929 & n14418 ) | ( n7929 & n15525 ) | ( n14418 & n15525 ) ;
  assign n15527 = n15525 | n15526 ;
  assign n15528 = ( n7930 & n15342 ) | ( n7930 & n15525 ) | ( n15342 & n15525 ) ;
  assign n15529 = n15527 | n15528 ;
  assign n15530 = n15529 ^ x8 ^ 1'b0 ;
  assign n15531 = n15504 & n15530 ;
  assign n15532 = n15523 | n15524 ;
  assign n15533 = n8034 & n15417 ;
  assign n15534 = n15532 | n15533 ;
  assign n15535 = n15479 ^ n14580 ^ n14578 ;
  assign n15536 = n15534 ^ x5 ^ 1'b0 ;
  assign n15537 = n15530 ^ n15504 ^ 1'b0 ;
  assign n15538 = ( n15508 & n15536 ) | ( n15508 & n15537 ) | ( n15536 & n15537 ) ;
  assign n15539 = n15537 ^ n15536 ^ n15508 ;
  assign n15540 = ( n14578 & n14580 ) | ( n14578 & n15479 ) | ( n14580 & n15479 ) ;
  assign n15541 = n8086 & n14569 ;
  assign n15542 = ( n8088 & n14578 ) | ( n8088 & n15541 ) | ( n14578 & n15541 ) ;
  assign n15543 = n15541 | n15542 ;
  assign n15544 = ( n8090 & n14580 ) | ( n8090 & n15541 ) | ( n14580 & n15541 ) ;
  assign n15545 = n15543 | n15544 ;
  assign n15546 = ~n8089 & n15535 ;
  assign n15547 = ( n15535 & n15545 ) | ( n15535 & ~n15546 ) | ( n15545 & ~n15546 ) ;
  assign n15548 = n15547 ^ x2 ^ 1'b0 ;
  assign n15549 = ( n15518 & n15539 ) | ( n15518 & n15548 ) | ( n15539 & n15548 ) ;
  assign n15550 = n6789 & n15535 ;
  assign n15551 = n6788 & ~n14580 ;
  assign n15552 = ( n6791 & n14578 ) | ( n6791 & n15550 ) | ( n14578 & n15550 ) ;
  assign n15553 = n15550 | n15552 ;
  assign n15554 = ( n6790 & n14569 ) | ( n6790 & n15550 ) | ( n14569 & n15550 ) ;
  assign n15555 = n15553 | n15554 ;
  assign n15556 = ( n6788 & ~n15551 ) | ( n6788 & n15555 ) | ( ~n15551 & n15555 ) ;
  assign n15557 = ( ~n6580 & n15490 ) | ( ~n6580 & n15556 ) | ( n15490 & n15556 ) ;
  assign n15558 = n15556 ^ n15490 ^ n6580 ;
  assign n15559 = n7932 & n14418 ;
  assign n15560 = ( n7929 & ~n14461 ) | ( n7929 & n15559 ) | ( ~n14461 & n15559 ) ;
  assign n15561 = ( n7943 & ~n14378 ) | ( n7943 & n15559 ) | ( ~n14378 & n15559 ) ;
  assign n15562 = n15559 | n15561 ;
  assign n15563 = n15560 | n15562 ;
  assign n15564 = n8029 & n14559 ;
  assign n15565 = n8034 & ~n15452 ;
  assign n15566 = ( n8037 & ~n14549 ) | ( n8037 & n15564 ) | ( ~n14549 & n15564 ) ;
  assign n15567 = n15564 | n15566 ;
  assign n15568 = ( n8033 & n14569 ) | ( n8033 & n15564 ) | ( n14569 & n15564 ) ;
  assign n15569 = n15567 | n15568 ;
  assign n15570 = n7930 & n15368 ;
  assign n15571 = ~n15565 & n15569 ;
  assign n15572 = n15571 ^ n15565 ^ x5 ;
  assign n15573 = n15563 | n15570 ;
  assign n15574 = n15573 ^ x8 ^ 1'b0 ;
  assign n15575 = n15574 ^ n15531 ^ n15351 ;
  assign n15576 = ( n15538 & n15572 ) | ( n15538 & n15575 ) | ( n15572 & n15575 ) ;
  assign n15577 = n15575 ^ n15572 ^ n15538 ;
  assign n15578 = n8086 & n14578 ;
  assign n15579 = ( n8088 & n14580 ) | ( n8088 & n15578 ) | ( n14580 & n15578 ) ;
  assign n15580 = n15578 | n15579 ;
  assign n15581 = ( n8090 & n14584 ) | ( n8090 & n15578 ) | ( n14584 & n15578 ) ;
  assign n15582 = n15580 | n15581 ;
  assign n15583 = n15540 ^ n14584 ^ n14580 ;
  assign n15584 = ( n15351 & n15531 ) | ( n15351 & n15574 ) | ( n15531 & n15574 ) ;
  assign n15585 = ~n8089 & n15583 ;
  assign n15586 = ( n15582 & n15583 ) | ( n15582 & ~n15585 ) | ( n15583 & ~n15585 ) ;
  assign n15587 = n15586 ^ x2 ^ 1'b0 ;
  assign n15588 = ( n15549 & n15577 ) | ( n15549 & n15587 ) | ( n15577 & n15587 ) ;
  assign n15589 = n6789 & n15583 ;
  assign n15590 = ( n6791 & n14580 ) | ( n6791 & n15589 ) | ( n14580 & n15589 ) ;
  assign n15591 = n15589 | n15590 ;
  assign n15592 = n6788 & ~n14584 ;
  assign n15593 = ( n6790 & n14578 ) | ( n6790 & n15589 ) | ( n14578 & n15589 ) ;
  assign n15594 = n15591 | n15593 ;
  assign n15595 = ( n6788 & ~n15592 ) | ( n6788 & n15594 ) | ( ~n15592 & n15594 ) ;
  assign n15596 = ( n14580 & n14584 ) | ( n14580 & n15540 ) | ( n14584 & n15540 ) ;
  assign n15597 = n15595 ^ n15557 ^ n6510 ;
  assign n15598 = ( ~n6510 & n15557 ) | ( ~n6510 & n15595 ) | ( n15557 & n15595 ) ;
  assign n15599 = x11 & ~n15351 ;
  assign n15600 = n7829 & ~n14324 ;
  assign n15601 = n7932 & ~n14461 ;
  assign n15602 = ( n7943 & n14418 ) | ( n7943 & n15601 ) | ( n14418 & n15601 ) ;
  assign n15603 = ( n7838 & n15326 ) | ( n7838 & n15600 ) | ( n15326 & n15600 ) ;
  assign n15604 = n15601 | n15602 ;
  assign n15605 = ( n7929 & ~n14549 ) | ( n7929 & n15601 ) | ( ~n14549 & n15601 ) ;
  assign n15606 = n15604 | n15605 ;
  assign n15607 = ( n7834 & ~n14378 ) | ( n7834 & n15600 ) | ( ~n14378 & n15600 ) ;
  assign n15608 = n15600 | n15603 ;
  assign n15609 = n15607 | n15608 ;
  assign n15610 = n7930 & ~n15405 ;
  assign n15611 = n7932 & ~n14549 ;
  assign n15612 = n15606 & ~n15610 ;
  assign n15613 = ( n7943 & ~n14461 ) | ( n7943 & n15611 ) | ( ~n14461 & n15611 ) ;
  assign n15614 = n15609 ^ x11 ^ 1'b0 ;
  assign n15615 = n15611 | n15613 ;
  assign n15616 = n15612 ^ n15610 ^ x8 ;
  assign n15617 = ( n7929 & n14559 ) | ( n7929 & n15611 ) | ( n14559 & n15611 ) ;
  assign n15618 = n15599 & n15614 ;
  assign n15619 = n15614 ^ n15599 ^ 1'b0 ;
  assign n15620 = n15615 | n15617 ;
  assign n15621 = n15619 ^ n15616 ^ n15584 ;
  assign n15622 = n8029 & n14569 ;
  assign n15623 = ( n15584 & n15616 ) | ( n15584 & n15619 ) | ( n15616 & n15619 ) ;
  assign n15624 = ( n8033 & n14578 ) | ( n8033 & n15622 ) | ( n14578 & n15622 ) ;
  assign n15625 = ( n8037 & n14559 ) | ( n8037 & n15622 ) | ( n14559 & n15622 ) ;
  assign n15626 = n15622 | n15625 ;
  assign n15627 = n15624 | n15626 ;
  assign n15628 = n8086 & n14580 ;
  assign n15629 = n8034 & n15475 ;
  assign n15630 = n15627 | n15629 ;
  assign n15631 = ( n8088 & n14584 ) | ( n8088 & n15628 ) | ( n14584 & n15628 ) ;
  assign n15632 = n15628 | n15631 ;
  assign n15633 = ( n8090 & ~n14583 ) | ( n8090 & n15628 ) | ( ~n14583 & n15628 ) ;
  assign n15634 = n15632 | n15633 ;
  assign n15635 = n15630 ^ x5 ^ 1'b0 ;
  assign n15636 = n15635 ^ n15621 ^ n15576 ;
  assign n15637 = ( n15576 & n15621 ) | ( n15576 & n15635 ) | ( n15621 & n15635 ) ;
  assign n15638 = n15596 ^ n14584 ^ n14583 ;
  assign n15639 = n7930 & n15417 ;
  assign n15640 = ( ~n14583 & n14584 ) | ( ~n14583 & n15596 ) | ( n14584 & n15596 ) ;
  assign n15641 = n15620 | n15639 ;
  assign n15642 = ~n15634 & n15638 ;
  assign n15643 = ( n8089 & n15634 ) | ( n8089 & ~n15642 ) | ( n15634 & ~n15642 ) ;
  assign n15644 = n7829 & ~n14378 ;
  assign n15645 = n15643 ^ x2 ^ 1'b0 ;
  assign n15646 = ( n15588 & n15636 ) | ( n15588 & n15645 ) | ( n15636 & n15645 ) ;
  assign n15647 = n8029 & n14578 ;
  assign n15648 = ( n8037 & n14569 ) | ( n8037 & n15647 ) | ( n14569 & n15647 ) ;
  assign n15649 = n15647 | n15648 ;
  assign n15650 = ( n8033 & n14580 ) | ( n8033 & n15647 ) | ( n14580 & n15647 ) ;
  assign n15651 = n15649 | n15650 ;
  assign n15652 = ( n7833 & ~n14324 ) | ( n7833 & n15644 ) | ( ~n14324 & n15644 ) ;
  assign n15653 = n15644 | n15652 ;
  assign n15654 = n15641 ^ x8 ^ 1'b0 ;
  assign n15655 = ( n7834 & n14418 ) | ( n7834 & n15653 ) | ( n14418 & n15653 ) ;
  assign n15656 = n15653 | n15655 ;
  assign n15657 = ( n7838 & n15342 ) | ( n7838 & n15653 ) | ( n15342 & n15653 ) ;
  assign n15658 = n15656 | n15657 ;
  assign n15659 = n15658 ^ x11 ^ 1'b0 ;
  assign n15660 = n15659 ^ n15618 ^ 1'b0 ;
  assign n15661 = n15618 & n15659 ;
  assign n15662 = ( n15623 & n15654 ) | ( n15623 & n15660 ) | ( n15654 & n15660 ) ;
  assign n15663 = n15660 ^ n15654 ^ n15623 ;
  assign n15664 = n8086 & n14584 ;
  assign n15665 = ( n8088 & ~n14583 ) | ( n8088 & n15664 ) | ( ~n14583 & n15664 ) ;
  assign n15666 = n15664 | n15665 ;
  assign n15667 = ( n8090 & n14599 ) | ( n8090 & n15664 ) | ( n14599 & n15664 ) ;
  assign n15668 = n15666 | n15667 ;
  assign n15669 = ( n8034 & n15535 ) | ( n8034 & n15651 ) | ( n15535 & n15651 ) ;
  assign n15670 = n15651 | n15669 ;
  assign n15671 = n15670 ^ x5 ^ 1'b0 ;
  assign n15672 = ( n15637 & n15663 ) | ( n15637 & n15671 ) | ( n15663 & n15671 ) ;
  assign n15673 = n15671 ^ n15663 ^ n15637 ;
  assign n15674 = n15640 ^ n14599 ^ n14583 ;
  assign n15675 = ( ~n14583 & n14599 ) | ( ~n14583 & n15640 ) | ( n14599 & n15640 ) ;
  assign n15676 = ~n15668 & n15674 ;
  assign n15677 = ( n8089 & n15668 ) | ( n8089 & ~n15676 ) | ( n15668 & ~n15676 ) ;
  assign n15678 = n15677 ^ x2 ^ 1'b0 ;
  assign n15679 = ( n15646 & n15673 ) | ( n15646 & n15678 ) | ( n15673 & n15678 ) ;
  assign n15680 = n6788 & ~n14583 ;
  assign n15681 = n6789 & ~n15638 ;
  assign n15682 = ( n6791 & n14584 ) | ( n6791 & n15681 ) | ( n14584 & n15681 ) ;
  assign n15683 = ( n6790 & n14580 ) | ( n6790 & n15681 ) | ( n14580 & n15681 ) ;
  assign n15684 = n15681 | n15682 ;
  assign n15685 = n15683 | n15684 ;
  assign n15686 = n15680 | n15685 ;
  assign n15687 = ( ~n6699 & n15598 ) | ( ~n6699 & n15686 ) | ( n15598 & n15686 ) ;
  assign n15688 = n15686 ^ n15598 ^ n6699 ;
  assign n15689 = n7932 & n14559 ;
  assign n15690 = n7829 & n14418 ;
  assign n15691 = ( n7833 & ~n14378 ) | ( n7833 & n15690 ) | ( ~n14378 & n15690 ) ;
  assign n15692 = ( n7834 & ~n14461 ) | ( n7834 & n15690 ) | ( ~n14461 & n15690 ) ;
  assign n15693 = n15690 | n15691 ;
  assign n15694 = ( n7943 & ~n14549 ) | ( n7943 & n15689 ) | ( ~n14549 & n15689 ) ;
  assign n15695 = n15692 | n15693 ;
  assign n15696 = n7838 & n15368 ;
  assign n15697 = n15695 | n15696 ;
  assign n15698 = n15697 ^ x11 ^ 1'b0 ;
  assign n15699 = ( n15390 & n15661 ) | ( n15390 & n15698 ) | ( n15661 & n15698 ) ;
  assign n15700 = n15689 | n15694 ;
  assign n15701 = n15698 ^ n15661 ^ n15390 ;
  assign n15702 = n8029 & n14580 ;
  assign n15703 = ( n7929 & n14569 ) | ( n7929 & n15689 ) | ( n14569 & n15689 ) ;
  assign n15704 = n15700 | n15703 ;
  assign n15705 = n7930 & ~n15452 ;
  assign n15706 = n15704 & ~n15705 ;
  assign n15707 = n15706 ^ n15705 ^ x8 ;
  assign n15708 = n15707 ^ n15701 ^ n15662 ;
  assign n15709 = ( n15662 & n15701 ) | ( n15662 & n15707 ) | ( n15701 & n15707 ) ;
  assign n15710 = ( n8033 & n14584 ) | ( n8033 & n15702 ) | ( n14584 & n15702 ) ;
  assign n15711 = ( n8037 & n14578 ) | ( n8037 & n15702 ) | ( n14578 & n15702 ) ;
  assign n15712 = n15702 | n15711 ;
  assign n15713 = n15710 | n15712 ;
  assign n15714 = ( n8034 & n15583 ) | ( n8034 & n15713 ) | ( n15583 & n15713 ) ;
  assign n15715 = n15713 | n15714 ;
  assign n15716 = n15715 ^ x5 ^ 1'b0 ;
  assign n15717 = n15716 ^ n15708 ^ n15672 ;
  assign n15718 = ( n15672 & n15708 ) | ( n15672 & n15716 ) | ( n15708 & n15716 ) ;
  assign n15719 = n8086 & ~n14583 ;
  assign n15720 = ( n8090 & ~n14610 ) | ( n8090 & n15719 ) | ( ~n14610 & n15719 ) ;
  assign n15721 = ( n8088 & n14599 ) | ( n8088 & n15719 ) | ( n14599 & n15719 ) ;
  assign n15722 = n15719 | n15721 ;
  assign n15723 = n15720 | n15722 ;
  assign n15724 = n15675 ^ n14610 ^ n14599 ;
  assign n15725 = ~n15723 & n15724 ;
  assign n15726 = ( n8089 & n15723 ) | ( n8089 & ~n15725 ) | ( n15723 & ~n15725 ) ;
  assign n15727 = n15726 ^ x2 ^ 1'b0 ;
  assign n15728 = ( n15679 & n15717 ) | ( n15679 & n15727 ) | ( n15717 & n15727 ) ;
  assign n15729 = n7829 & ~n14461 ;
  assign n15730 = ( n7833 & n14418 ) | ( n7833 & n15729 ) | ( n14418 & n15729 ) ;
  assign n15731 = n15729 | n15730 ;
  assign n15732 = x14 & ~n15390 ;
  assign n15733 = ( n7834 & ~n14549 ) | ( n7834 & n15729 ) | ( ~n14549 & n15729 ) ;
  assign n15734 = n15731 | n15733 ;
  assign n15735 = n6789 & ~n15674 ;
  assign n15736 = ( n6791 & ~n14583 ) | ( n6791 & n15735 ) | ( ~n14583 & n15735 ) ;
  assign n15737 = n15735 | n15736 ;
  assign n15738 = ( n6790 & n14584 ) | ( n6790 & n15735 ) | ( n14584 & n15735 ) ;
  assign n15739 = n15737 | n15738 ;
  assign n15740 = n6788 & ~n14599 ;
  assign n15741 = ( n6788 & n15739 ) | ( n6788 & ~n15740 ) | ( n15739 & ~n15740 ) ;
  assign n15742 = n7838 & ~n15405 ;
  assign n15743 = n15734 & ~n15742 ;
  assign n15744 = n15743 ^ n15742 ^ x11 ;
  assign n15745 = ( ~n6781 & n15687 ) | ( ~n6781 & n15741 ) | ( n15687 & n15741 ) ;
  assign n15746 = n15741 ^ n15687 ^ n6781 ;
  assign n15747 = n7669 & ~n14324 ;
  assign n15748 = ( n7666 & n15326 ) | ( n7666 & n15747 ) | ( n15326 & n15747 ) ;
  assign n15749 = n15747 | n15748 ;
  assign n15750 = ( n7667 & ~n14378 ) | ( n7667 & n15747 ) | ( ~n14378 & n15747 ) ;
  assign n15751 = n15749 | n15750 ;
  assign n15752 = n15751 ^ x14 ^ 1'b0 ;
  assign n15753 = n15752 ^ n15732 ^ 1'b0 ;
  assign n15754 = n15732 & n15752 ;
  assign n15755 = n15753 ^ n15744 ^ n15699 ;
  assign n15756 = ( n15699 & n15744 ) | ( n15699 & n15753 ) | ( n15744 & n15753 ) ;
  assign n15757 = n7932 & n14569 ;
  assign n15758 = ( n7943 & n14559 ) | ( n7943 & n15757 ) | ( n14559 & n15757 ) ;
  assign n15759 = n15757 | n15758 ;
  assign n15760 = ( n7929 & n14578 ) | ( n7929 & n15757 ) | ( n14578 & n15757 ) ;
  assign n15761 = n7930 & n15475 ;
  assign n15762 = n15759 | n15760 ;
  assign n15763 = n15761 | n15762 ;
  assign n15764 = n15763 ^ x8 ^ 1'b0 ;
  assign n15765 = n15764 ^ n15755 ^ n15709 ;
  assign n15766 = ( n15709 & n15755 ) | ( n15709 & n15764 ) | ( n15755 & n15764 ) ;
  assign n15767 = n6901 & n14418 ;
  assign n15768 = n8029 & n14584 ;
  assign n15769 = ( n6907 & ~n14461 ) | ( n6907 & n15767 ) | ( ~n14461 & n15767 ) ;
  assign n15770 = ( n8037 & n14580 ) | ( n8037 & n15768 ) | ( n14580 & n15768 ) ;
  assign n15771 = n15768 | n15770 ;
  assign n15772 = ( n8033 & ~n14583 ) | ( n8033 & n15768 ) | ( ~n14583 & n15768 ) ;
  assign n15773 = n15771 | n15772 ;
  assign n15774 = n8034 & ~n15638 ;
  assign n15775 = n15773 & ~n15774 ;
  assign n15776 = n15775 ^ n15774 ^ x5 ;
  assign n15777 = ( n15718 & n15765 ) | ( n15718 & n15776 ) | ( n15765 & n15776 ) ;
  assign n15778 = n15776 ^ n15765 ^ n15718 ;
  assign n15779 = n6901 & ~n14549 ;
  assign n15780 = ( n6906 & ~n14378 ) | ( n6906 & n15767 ) | ( ~n14378 & n15767 ) ;
  assign n15781 = n15767 | n15780 ;
  assign n15782 = n15769 | n15781 ;
  assign n15783 = ( n6906 & ~n14461 ) | ( n6906 & n15779 ) | ( ~n14461 & n15779 ) ;
  assign n15784 = ( n6907 & n14559 ) | ( n6907 & n15779 ) | ( n14559 & n15779 ) ;
  assign n15785 = n15779 | n15783 ;
  assign n15786 = n15784 | n15785 ;
  assign n15787 = n6901 & ~n14461 ;
  assign n15788 = ( n6906 & n14418 ) | ( n6906 & n15787 ) | ( n14418 & n15787 ) ;
  assign n15789 = n15787 | n15788 ;
  assign n15790 = ( n6907 & ~n14549 ) | ( n6907 & n15787 ) | ( ~n14549 & n15787 ) ;
  assign n15791 = n15789 | n15790 ;
  assign n15792 = n6918 & n15417 ;
  assign n15793 = n15786 | n15792 ;
  assign n15794 = n15793 ^ x29 ^ 1'b0 ;
  assign n15795 = n6918 & ~n15405 ;
  assign n15796 = n15791 | n15795 ;
  assign n15797 = n6918 & n15368 ;
  assign n15798 = n15782 | n15797 ;
  assign n15799 = n15796 ^ x29 ^ 1'b0 ;
  assign n15800 = n15798 ^ x29 ^ 1'b0 ;
  assign n15801 = n6901 & ~n14378 ;
  assign n15802 = ( n6906 & ~n14324 ) | ( n6906 & n15801 ) | ( ~n14324 & n15801 ) ;
  assign n15803 = n15801 | n15802 ;
  assign n15804 = ( n6907 & n14418 ) | ( n6907 & n15803 ) | ( n14418 & n15803 ) ;
  assign n15805 = n6918 & n15326 ;
  assign n15806 = ( n6918 & n15342 ) | ( n6918 & n15803 ) | ( n15342 & n15803 ) ;
  assign n15807 = n15803 | n15804 ;
  assign n15808 = x29 & ~n15391 ;
  assign n15809 = n15806 | n15807 ;
  assign n15810 = ( n6901 & ~n14324 ) | ( n6901 & n15805 ) | ( ~n14324 & n15805 ) ;
  assign n15811 = n15805 | n15810 ;
  assign n15812 = ( n6907 & ~n14378 ) | ( n6907 & n15805 ) | ( ~n14378 & n15805 ) ;
  assign n15813 = n15811 | n15812 ;
  assign n15814 = n15813 ^ x29 ^ 1'b0 ;
  assign n15815 = n15808 & n15814 ;
  assign n15816 = n15809 ^ x29 ^ 1'b0 ;
  assign n15817 = n15814 ^ n15808 ^ 1'b0 ;
  assign n15818 = n15815 & n15816 ;
  assign n15819 = n15816 ^ n15815 ^ 1'b0 ;
  assign n15820 = ( n15388 & n15800 ) | ( n15388 & n15818 ) | ( n15800 & n15818 ) ;
  assign n15821 = n15818 ^ n15800 ^ n15388 ;
  assign n15822 = n6901 & n14569 ;
  assign n15823 = ( n6906 & n14559 ) | ( n6906 & n15822 ) | ( n14559 & n15822 ) ;
  assign n15824 = n15822 | n15823 ;
  assign n15825 = ( n6907 & n14578 ) | ( n6907 & n15822 ) | ( n14578 & n15822 ) ;
  assign n15826 = n15824 | n15825 ;
  assign n15827 = ( ~n15338 & n15799 ) | ( ~n15338 & n15820 ) | ( n15799 & n15820 ) ;
  assign n15828 = n15820 ^ n15799 ^ n15338 ;
  assign n15829 = ( ~n15345 & n15794 ) | ( ~n15345 & n15827 ) | ( n15794 & n15827 ) ;
  assign n15830 = n6901 & n14559 ;
  assign n15831 = n15827 ^ n15794 ^ n15345 ;
  assign n15832 = ( n6906 & ~n14549 ) | ( n6906 & n15830 ) | ( ~n14549 & n15830 ) ;
  assign n15833 = n15830 | n15832 ;
  assign n15834 = n6918 & n15475 ;
  assign n15835 = ( n6907 & n14569 ) | ( n6907 & n15830 ) | ( n14569 & n15830 ) ;
  assign n15836 = n15833 | n15835 ;
  assign n15837 = n15826 | n15834 ;
  assign n15838 = n6918 & ~n15452 ;
  assign n15839 = n15836 | n15838 ;
  assign n15840 = n15839 ^ x29 ^ 1'b0 ;
  assign n15841 = n15837 ^ x29 ^ 1'b0 ;
  assign n15842 = n15840 ^ n15829 ^ n15376 ;
  assign n15843 = ( n15376 & n15829 ) | ( n15376 & n15840 ) | ( n15829 & n15840 ) ;
  assign n15844 = n15843 ^ n15841 ^ n15426 ;
  assign n15845 = ( ~n15426 & n15841 ) | ( ~n15426 & n15843 ) | ( n15841 & n15843 ) ;
  assign n15846 = n6901 & n14578 ;
  assign n15847 = ( n6906 & n14569 ) | ( n6906 & n15846 ) | ( n14569 & n15846 ) ;
  assign n15848 = n15846 | n15847 ;
  assign n15849 = ( n6907 & n14580 ) | ( n6907 & n15846 ) | ( n14580 & n15846 ) ;
  assign n15850 = n15848 | n15849 ;
  assign n15851 = n6918 & n15535 ;
  assign n15852 = n15850 | n15851 ;
  assign n15853 = n15852 ^ x29 ^ 1'b0 ;
  assign n15854 = n15853 ^ n15845 ^ n15436 ;
  assign n15855 = ( ~n15436 & n15845 ) | ( ~n15436 & n15853 ) | ( n15845 & n15853 ) ;
  assign n15856 = n6901 & n14580 ;
  assign n15857 = ( n6906 & n14578 ) | ( n6906 & n15856 ) | ( n14578 & n15856 ) ;
  assign n15858 = n15856 | n15857 ;
  assign n15859 = ( n6907 & n14584 ) | ( n6907 & n15856 ) | ( n14584 & n15856 ) ;
  assign n15860 = n15858 | n15859 ;
  assign n15861 = ( n6918 & n15583 ) | ( n6918 & n15860 ) | ( n15583 & n15860 ) ;
  assign n15862 = n15860 | n15861 ;
  assign n15863 = n15862 ^ x29 ^ 1'b0 ;
  assign n15864 = ( ~n15480 & n15855 ) | ( ~n15480 & n15863 ) | ( n15855 & n15863 ) ;
  assign n15865 = n15863 ^ n15855 ^ n15480 ;
  assign n15866 = n6901 & n14584 ;
  assign n15867 = ( n6906 & n14580 ) | ( n6906 & n15866 ) | ( n14580 & n15866 ) ;
  assign n15868 = n15866 | n15867 ;
  assign n15869 = ( n6907 & ~n14583 ) | ( n6907 & n15866 ) | ( ~n14583 & n15866 ) ;
  assign n15870 = n15868 | n15869 ;
  assign n15871 = n6918 & ~n15638 ;
  assign n15872 = n15870 & ~n15871 ;
  assign n15873 = n15872 ^ n15871 ^ x29 ;
  assign n15874 = ( n15491 & n15864 ) | ( n15491 & n15873 ) | ( n15864 & n15873 ) ;
  assign n15875 = n15873 ^ n15864 ^ n15491 ;
  assign n15876 = n6901 & ~n14583 ;
  assign n15877 = ( n6906 & n14584 ) | ( n6906 & n15876 ) | ( n14584 & n15876 ) ;
  assign n15878 = n15876 | n15877 ;
  assign n15879 = ( n6907 & n14599 ) | ( n6907 & n15878 ) | ( n14599 & n15878 ) ;
  assign n15880 = n15878 | n15879 ;
  assign n15881 = ( n6918 & ~n15674 ) | ( n6918 & n15878 ) | ( ~n15674 & n15878 ) ;
  assign n15882 = n15880 | n15881 ;
  assign n15883 = n15882 ^ x29 ^ 1'b0 ;
  assign n15884 = ( ~n15558 & n15874 ) | ( ~n15558 & n15883 ) | ( n15874 & n15883 ) ;
  assign n15885 = n15883 ^ n15874 ^ n15558 ;
  assign n15886 = n6901 & n14599 ;
  assign n15887 = ( n6906 & ~n14583 ) | ( n6906 & n15886 ) | ( ~n14583 & n15886 ) ;
  assign n15888 = n15886 | n15887 ;
  assign n15889 = ( n6907 & ~n14610 ) | ( n6907 & n15886 ) | ( ~n14610 & n15886 ) ;
  assign n15890 = n15888 | n15889 ;
  assign n15891 = n6918 & ~n15724 ;
  assign n15892 = n15890 & ~n15891 ;
  assign n15893 = n15892 ^ n15891 ^ x29 ;
  assign n15894 = n7838 & n15417 ;
  assign n15895 = n15893 ^ n15884 ^ n15597 ;
  assign n15896 = ( ~n15597 & n15884 ) | ( ~n15597 & n15893 ) | ( n15884 & n15893 ) ;
  assign n15897 = n7829 & ~n14549 ;
  assign n15898 = ( n7833 & ~n14461 ) | ( n7833 & n15897 ) | ( ~n14461 & n15897 ) ;
  assign n15899 = n15897 | n15898 ;
  assign n15900 = ( n7834 & n14559 ) | ( n7834 & n15897 ) | ( n14559 & n15897 ) ;
  assign n15901 = n15899 | n15900 ;
  assign n15902 = n15894 | n15901 ;
  assign n15903 = n7669 & ~n14378 ;
  assign n15904 = ( n7674 & ~n14324 ) | ( n7674 & n15903 ) | ( ~n14324 & n15903 ) ;
  assign n15905 = n15903 | n15904 ;
  assign n15906 = ( n7667 & n14418 ) | ( n7667 & n15905 ) | ( n14418 & n15905 ) ;
  assign n15907 = n15905 | n15906 ;
  assign n15908 = n15902 ^ x11 ^ 1'b0 ;
  assign n15909 = ( n7666 & n15342 ) | ( n7666 & n15905 ) | ( n15342 & n15905 ) ;
  assign n15910 = n15907 | n15909 ;
  assign n15911 = n15910 ^ x14 ^ 1'b0 ;
  assign n15912 = n15911 ^ n15754 ^ 1'b0 ;
  assign n15913 = n15754 & n15911 ;
  assign n15914 = ( n15756 & n15908 ) | ( n15756 & n15912 ) | ( n15908 & n15912 ) ;
  assign n15915 = n15912 ^ n15908 ^ n15756 ;
  assign n15916 = n7932 & n14578 ;
  assign n15917 = ( n7943 & n14569 ) | ( n7943 & n15916 ) | ( n14569 & n15916 ) ;
  assign n15918 = n15916 | n15917 ;
  assign n15919 = ( n7929 & n14580 ) | ( n7929 & n15916 ) | ( n14580 & n15916 ) ;
  assign n15920 = n15918 | n15919 ;
  assign n15921 = ( n7930 & n15535 ) | ( n7930 & n15920 ) | ( n15535 & n15920 ) ;
  assign n15922 = n15920 | n15921 ;
  assign n15923 = n15922 ^ x8 ^ 1'b0 ;
  assign n15924 = ( n15766 & n15915 ) | ( n15766 & n15923 ) | ( n15915 & n15923 ) ;
  assign n15925 = n15923 ^ n15915 ^ n15766 ;
  assign n15926 = n8029 & ~n14583 ;
  assign n15927 = ( n8037 & n14584 ) | ( n8037 & n15926 ) | ( n14584 & n15926 ) ;
  assign n15928 = n15926 | n15927 ;
  assign n15929 = ( n8033 & n14599 ) | ( n8033 & n15926 ) | ( n14599 & n15926 ) ;
  assign n15930 = n15928 | n15929 ;
  assign n15931 = n8034 & ~n15674 ;
  assign n15932 = n15930 | n15931 ;
  assign n15933 = n15932 ^ x5 ^ 1'b0 ;
  assign n15934 = n15933 ^ n15925 ^ n15777 ;
  assign n15935 = ( n15777 & n15925 ) | ( n15777 & n15933 ) | ( n15925 & n15933 ) ;
  assign n15936 = n7190 & ~n14324 ;
  assign n15937 = n7188 & ~n14378 ;
  assign n15938 = ( n7192 & ~n14378 ) | ( n7192 & n15936 ) | ( ~n14378 & n15936 ) ;
  assign n15939 = ( n7196 & n15326 ) | ( n7196 & n15937 ) | ( n15326 & n15937 ) ;
  assign n15940 = ( n7192 & ~n14324 ) | ( n7192 & n15937 ) | ( ~n14324 & n15937 ) ;
  assign n15941 = n15936 | n15938 ;
  assign n15942 = ( n7196 & n15342 ) | ( n7196 & n15941 ) | ( n15342 & n15941 ) ;
  assign n15943 = ( n7188 & n14418 ) | ( n7188 & n15941 ) | ( n14418 & n15941 ) ;
  assign n15944 = n15941 | n15943 ;
  assign n15945 = n7188 & ~n14549 ;
  assign n15946 = n15942 | n15944 ;
  assign n15947 = x23 & ~n15349 ;
  assign n15948 = n15937 | n15939 ;
  assign n15949 = n15946 ^ x23 ^ 1'b0 ;
  assign n15950 = n15940 | n15948 ;
  assign n15951 = n15950 ^ x23 ^ 1'b0 ;
  assign n15952 = ( n7190 & n14418 ) | ( n7190 & n15945 ) | ( n14418 & n15945 ) ;
  assign n15953 = n15947 & n15951 ;
  assign n15954 = ( n7192 & ~n14461 ) | ( n7192 & n15945 ) | ( ~n14461 & n15945 ) ;
  assign n15955 = n15945 | n15952 ;
  assign n15956 = n15954 | n15955 ;
  assign n15957 = n15953 ^ n15949 ^ 1'b0 ;
  assign n15958 = n7188 & ~n14461 ;
  assign n15959 = n15949 & n15953 ;
  assign n15960 = n7196 & ~n15405 ;
  assign n15961 = n15956 & ~n15960 ;
  assign n15962 = n15961 ^ n15960 ^ x23 ;
  assign n15963 = ( n7190 & ~n14378 ) | ( n7190 & n15958 ) | ( ~n14378 & n15958 ) ;
  assign n15964 = n15958 | n15963 ;
  assign n15965 = ( n7192 & n14418 ) | ( n7192 & n15958 ) | ( n14418 & n15958 ) ;
  assign n15966 = n15964 | n15965 ;
  assign n15967 = n7196 & n15368 ;
  assign n15968 = n15966 | n15967 ;
  assign n15969 = n15968 ^ x23 ^ 1'b0 ;
  assign n15970 = ( n15381 & n15959 ) | ( n15381 & n15969 ) | ( n15959 & n15969 ) ;
  assign n15971 = n15969 ^ n15959 ^ n15381 ;
  assign n15972 = x26 & ~n15381 ;
  assign n15973 = n15951 ^ n15947 ^ 1'b0 ;
  assign n15974 = n7037 & ~n14378 ;
  assign n15975 = ( n7036 & ~n14324 ) | ( n7036 & n15974 ) | ( ~n14324 & n15974 ) ;
  assign n15976 = n15974 | n15975 ;
  assign n15977 = ( n7035 & n15326 ) | ( n7035 & n15974 ) | ( n15326 & n15974 ) ;
  assign n15978 = n15976 | n15977 ;
  assign n15979 = n15978 ^ x26 ^ 1'b0 ;
  assign n15980 = n15979 ^ n15972 ^ 1'b0 ;
  assign n15981 = n15972 & n15979 ;
  assign n15982 = n15980 ^ n15970 ^ n15962 ;
  assign n15983 = ( n15962 & n15970 ) | ( n15962 & n15980 ) | ( n15970 & n15980 ) ;
  assign n15984 = n7340 & n15326 ;
  assign n15985 = ( n7339 & ~n14324 ) | ( n7339 & n15984 ) | ( ~n14324 & n15984 ) ;
  assign n15986 = ( n7337 & ~n14378 ) | ( n7337 & n15984 ) | ( ~n14378 & n15984 ) ;
  assign n15987 = n15984 | n15985 ;
  assign n15988 = n15986 | n15987 ;
  assign n15989 = n7485 & ~n14324 ;
  assign n15990 = n7036 & ~n14378 ;
  assign n15991 = ( n7052 & ~n14324 ) | ( n7052 & n15990 ) | ( ~n14324 & n15990 ) ;
  assign n15992 = n15990 | n15991 ;
  assign n15993 = ( n7037 & n14418 ) | ( n7037 & n15992 ) | ( n14418 & n15992 ) ;
  assign n15994 = ( n7487 & n15326 ) | ( n7487 & n15989 ) | ( n15326 & n15989 ) ;
  assign n15995 = n15989 | n15994 ;
  assign n15996 = ( n7486 & ~n14378 ) | ( n7486 & n15989 ) | ( ~n14378 & n15989 ) ;
  assign n15997 = n15992 | n15993 ;
  assign n15998 = ( n7035 & n15342 ) | ( n7035 & n15992 ) | ( n15342 & n15992 ) ;
  assign n15999 = n15995 | n15996 ;
  assign n16000 = n15997 | n15998 ;
  assign n16001 = n7485 & ~n14378 ;
  assign n16002 = n15988 ^ x20 ^ 1'b0 ;
  assign n16003 = n16000 ^ x26 ^ 1'b0 ;
  assign n16004 = ( n7493 & ~n14324 ) | ( n7493 & n16001 ) | ( ~n14324 & n16001 ) ;
  assign n16005 = n16001 | n16004 ;
  assign n16006 = n7339 & ~n14378 ;
  assign n16007 = ( n7338 & ~n14324 ) | ( n7338 & n16006 ) | ( ~n14324 & n16006 ) ;
  assign n16008 = n16006 | n16007 ;
  assign n16009 = ( n7486 & n14418 ) | ( n7486 & n16005 ) | ( n14418 & n16005 ) ;
  assign n16010 = n16005 | n16009 ;
  assign n16011 = ( n7487 & n15342 ) | ( n7487 & n16005 ) | ( n15342 & n16005 ) ;
  assign n16012 = n16010 | n16011 ;
  assign n16013 = n15981 & n16003 ;
  assign n16014 = n16003 ^ n15981 ^ 1'b0 ;
  assign n16015 = n16012 ^ x17 ^ 1'b0 ;
  assign n16016 = n15999 ^ x17 ^ 1'b0 ;
  assign n16017 = ( n7340 & n15342 ) | ( n7340 & n16008 ) | ( n15342 & n16008 ) ;
  assign n16018 = ( n7337 & n14418 ) | ( n7337 & n16008 ) | ( n14418 & n16008 ) ;
  assign n16019 = n16008 | n16018 ;
  assign n16020 = n7037 & ~n14461 ;
  assign n16021 = n16017 | n16019 ;
  assign n16022 = n16021 ^ x20 ^ 1'b0 ;
  assign n16023 = ( n7036 & n14418 ) | ( n7036 & n16020 ) | ( n14418 & n16020 ) ;
  assign n16024 = n16020 | n16023 ;
  assign n16025 = ( n7052 & ~n14378 ) | ( n7052 & n16020 ) | ( ~n14378 & n16020 ) ;
  assign n16026 = n16024 | n16025 ;
  assign n16027 = n7035 & n15368 ;
  assign n16028 = n16026 | n16027 ;
  assign n16029 = n16028 ^ x26 ^ 1'b0 ;
  assign n16030 = n16029 ^ n16013 ^ n15391 ;
  assign n16031 = ( n15391 & n16013 ) | ( n15391 & n16029 ) | ( n16013 & n16029 ) ;
  assign n16032 = n7037 & ~n14549 ;
  assign n16033 = ( n7036 & ~n14461 ) | ( n7036 & n16032 ) | ( ~n14461 & n16032 ) ;
  assign n16034 = n16032 | n16033 ;
  assign n16035 = ( n7052 & n14418 ) | ( n7052 & n16032 ) | ( n14418 & n16032 ) ;
  assign n16036 = n16034 | n16035 ;
  assign n16037 = n7035 & ~n15405 ;
  assign n16038 = n16036 & ~n16037 ;
  assign n16039 = n16038 ^ n16037 ^ x26 ;
  assign n16040 = n16039 ^ n16031 ^ n15817 ;
  assign n16041 = ( n15817 & n16031 ) | ( n15817 & n16039 ) | ( n16031 & n16039 ) ;
  assign n16042 = n7485 & n14418 ;
  assign n16043 = ( n7493 & ~n14378 ) | ( n7493 & n16042 ) | ( ~n14378 & n16042 ) ;
  assign n16044 = ( n7486 & ~n14461 ) | ( n7486 & n16042 ) | ( ~n14461 & n16042 ) ;
  assign n16045 = n16042 | n16044 ;
  assign n16046 = n7339 & n14418 ;
  assign n16047 = n16043 | n16045 ;
  assign n16048 = ( n7337 & ~n14461 ) | ( n7337 & n16046 ) | ( ~n14461 & n16046 ) ;
  assign n16049 = n16046 | n16048 ;
  assign n16050 = ( n7338 & ~n14378 ) | ( n7338 & n16046 ) | ( ~n14378 & n16046 ) ;
  assign n16051 = n16049 | n16050 ;
  assign n16052 = n7669 & n14418 ;
  assign n16053 = ( n7674 & ~n14378 ) | ( n7674 & n16052 ) | ( ~n14378 & n16052 ) ;
  assign n16054 = n16052 | n16053 ;
  assign n16055 = ( n7667 & ~n14461 ) | ( n7667 & n16052 ) | ( ~n14461 & n16052 ) ;
  assign n16056 = n16054 | n16055 ;
  assign n16057 = n7340 & n15368 ;
  assign n16058 = n16051 | n16057 ;
  assign n16059 = n7666 & n15368 ;
  assign n16060 = n16056 | n16059 ;
  assign n16061 = n16060 ^ x14 ^ 1'b0 ;
  assign n16062 = n16061 ^ n15913 ^ n15348 ;
  assign n16063 = n7487 & n15368 ;
  assign n16064 = ( n15348 & n15913 ) | ( n15348 & n16061 ) | ( n15913 & n16061 ) ;
  assign n16065 = n7485 & ~n14461 ;
  assign n16066 = n16047 | n16063 ;
  assign n16067 = ( n7486 & ~n14549 ) | ( n7486 & n16065 ) | ( ~n14549 & n16065 ) ;
  assign n16068 = n16065 | n16067 ;
  assign n16069 = ( n7493 & n14418 ) | ( n7493 & n16065 ) | ( n14418 & n16065 ) ;
  assign n16070 = n16068 | n16069 ;
  assign n16071 = x17 & ~n15348 ;
  assign n16072 = n16016 & n16071 ;
  assign n16073 = n16066 ^ x17 ^ 1'b0 ;
  assign n16074 = n16058 ^ x20 ^ 1'b0 ;
  assign n16075 = n16071 ^ n16016 ^ 1'b0 ;
  assign n16076 = n16015 & n16072 ;
  assign n16077 = n16072 ^ n16015 ^ 1'b0 ;
  assign n16078 = ( n15354 & n16073 ) | ( n15354 & n16076 ) | ( n16073 & n16076 ) ;
  assign n16079 = n16076 ^ n16073 ^ n15354 ;
  assign n16080 = n7487 & ~n15405 ;
  assign n16081 = n16070 & ~n16080 ;
  assign n16082 = x20 & ~n15354 ;
  assign n16083 = n16081 ^ n16080 ^ x17 ;
  assign n16084 = n16002 & n16082 ;
  assign n16085 = n16082 ^ n16002 ^ 1'b0 ;
  assign n16086 = n16084 ^ n16022 ^ 1'b0 ;
  assign n16087 = n16022 & n16084 ;
  assign n16088 = n16087 ^ n16074 ^ n15349 ;
  assign n16089 = ( n15349 & n16074 ) | ( n15349 & n16087 ) | ( n16074 & n16087 ) ;
  assign n16090 = n16085 ^ n16083 ^ n16078 ;
  assign n16091 = ( n16078 & n16083 ) | ( n16078 & n16085 ) | ( n16083 & n16085 ) ;
  assign n16092 = n7485 & ~n14549 ;
  assign n16093 = ( n7486 & n14559 ) | ( n7486 & n16092 ) | ( n14559 & n16092 ) ;
  assign n16094 = n16092 | n16093 ;
  assign n16095 = ( n7493 & ~n14461 ) | ( n7493 & n16092 ) | ( ~n14461 & n16092 ) ;
  assign n16096 = n16094 | n16095 ;
  assign n16097 = n7487 & n15417 ;
  assign n16098 = n16096 | n16097 ;
  assign n16099 = n16098 ^ x17 ^ 1'b0 ;
  assign n16100 = n16099 ^ n16091 ^ n16086 ;
  assign n16101 = ( n16086 & n16091 ) | ( n16086 & n16099 ) | ( n16091 & n16099 ) ;
  assign n16102 = n7485 & n14559 ;
  assign n16103 = ( n7486 & n14569 ) | ( n7486 & n16102 ) | ( n14569 & n16102 ) ;
  assign n16104 = n16102 | n16103 ;
  assign n16105 = ( n7493 & ~n14549 ) | ( n7493 & n16102 ) | ( ~n14549 & n16102 ) ;
  assign n16106 = n16104 | n16105 ;
  assign n16107 = n7487 & ~n15452 ;
  assign n16108 = n16106 & ~n16107 ;
  assign n16109 = n16108 ^ n16107 ^ x17 ;
  assign n16110 = n16109 ^ n16101 ^ n16088 ;
  assign n16111 = ( n16088 & n16101 ) | ( n16088 & n16109 ) | ( n16101 & n16109 ) ;
  assign n16112 = n7339 & ~n14461 ;
  assign n16113 = ( n7337 & ~n14549 ) | ( n7337 & n16112 ) | ( ~n14549 & n16112 ) ;
  assign n16114 = n16112 | n16113 ;
  assign n16115 = ( n7338 & n14418 ) | ( n7338 & n16112 ) | ( n14418 & n16112 ) ;
  assign n16116 = n16114 | n16115 ;
  assign n16117 = n7669 & ~n14461 ;
  assign n16118 = ( n7674 & n14418 ) | ( n7674 & n16117 ) | ( n14418 & n16117 ) ;
  assign n16119 = n16117 | n16118 ;
  assign n16120 = ( n7667 & ~n14549 ) | ( n7667 & n16117 ) | ( ~n14549 & n16117 ) ;
  assign n16121 = n16119 | n16120 ;
  assign n16122 = n7666 & ~n15405 ;
  assign n16123 = n7340 & ~n15405 ;
  assign n16124 = n16116 & ~n16123 ;
  assign n16125 = n16121 & ~n16122 ;
  assign n16126 = n16125 ^ n16122 ^ x14 ;
  assign n16127 = n16124 ^ n16123 ^ x20 ;
  assign n16128 = n7485 & n14569 ;
  assign n16129 = ( n7486 & n14578 ) | ( n7486 & n16128 ) | ( n14578 & n16128 ) ;
  assign n16130 = n16128 | n16129 ;
  assign n16131 = ( n7493 & n14559 ) | ( n7493 & n16128 ) | ( n14559 & n16128 ) ;
  assign n16132 = n16130 | n16131 ;
  assign n16133 = n16126 ^ n16075 ^ n16064 ;
  assign n16134 = ( n16064 & n16075 ) | ( n16064 & n16126 ) | ( n16075 & n16126 ) ;
  assign n16135 = ( n15973 & n16089 ) | ( n15973 & n16127 ) | ( n16089 & n16127 ) ;
  assign n16136 = n7487 & n15475 ;
  assign n16137 = n16127 ^ n16089 ^ n15973 ;
  assign n16138 = n16132 | n16136 ;
  assign n16139 = n16138 ^ x17 ^ 1'b0 ;
  assign n16140 = n16139 ^ n16137 ^ n16111 ;
  assign n16141 = ( n16111 & n16137 ) | ( n16111 & n16139 ) | ( n16137 & n16139 ) ;
  assign n16142 = n7037 & n14559 ;
  assign n16143 = ( n7036 & ~n14549 ) | ( n7036 & n16142 ) | ( ~n14549 & n16142 ) ;
  assign n16144 = n16142 | n16143 ;
  assign n16145 = ( n7052 & ~n14461 ) | ( n7052 & n16142 ) | ( ~n14461 & n16142 ) ;
  assign n16146 = n16144 | n16145 ;
  assign n16147 = n7035 & n15417 ;
  assign n16148 = n16146 | n16147 ;
  assign n16149 = n16148 ^ x26 ^ 1'b0 ;
  assign n16150 = n16149 ^ n16041 ^ n15819 ;
  assign n16151 = ( n15819 & n16041 ) | ( n15819 & n16149 ) | ( n16041 & n16149 ) ;
  assign n16152 = n7339 & ~n14549 ;
  assign n16153 = ( n7337 & n14559 ) | ( n7337 & n16152 ) | ( n14559 & n16152 ) ;
  assign n16154 = n16152 | n16153 ;
  assign n16155 = ( n7338 & ~n14461 ) | ( n7338 & n16152 ) | ( ~n14461 & n16152 ) ;
  assign n16156 = n16154 | n16155 ;
  assign n16157 = n7340 & n15417 ;
  assign n16158 = n16156 | n16157 ;
  assign n16159 = n16158 ^ x20 ^ 1'b0 ;
  assign n16160 = n16159 ^ n16135 ^ n15957 ;
  assign n16161 = ( n15957 & n16135 ) | ( n15957 & n16159 ) | ( n16135 & n16159 ) ;
  assign n16162 = n7188 & n14559 ;
  assign n16163 = ( n7190 & ~n14461 ) | ( n7190 & n16162 ) | ( ~n14461 & n16162 ) ;
  assign n16164 = n16162 | n16163 ;
  assign n16165 = ( n7192 & ~n14549 ) | ( n7192 & n16162 ) | ( ~n14549 & n16162 ) ;
  assign n16166 = n16164 | n16165 ;
  assign n16167 = n7669 & ~n14549 ;
  assign n16168 = ( n7674 & ~n14461 ) | ( n7674 & n16167 ) | ( ~n14461 & n16167 ) ;
  assign n16169 = n16167 | n16168 ;
  assign n16170 = ( n7667 & n14559 ) | ( n7667 & n16167 ) | ( n14559 & n16167 ) ;
  assign n16171 = n16169 | n16170 ;
  assign n16172 = n7666 & n15417 ;
  assign n16173 = n7196 & n15417 ;
  assign n16174 = n16166 | n16173 ;
  assign n16175 = n7188 & n14569 ;
  assign n16176 = n16171 | n16172 ;
  assign n16177 = n16174 ^ x23 ^ 1'b0 ;
  assign n16178 = n16177 ^ n16014 ^ n15983 ;
  assign n16179 = n16176 ^ x14 ^ 1'b0 ;
  assign n16180 = ( n15983 & n16014 ) | ( n15983 & n16177 ) | ( n16014 & n16177 ) ;
  assign n16181 = ( n16077 & n16134 ) | ( n16077 & n16179 ) | ( n16134 & n16179 ) ;
  assign n16182 = n16179 ^ n16134 ^ n16077 ;
  assign n16183 = ( n7190 & ~n14549 ) | ( n7190 & n16175 ) | ( ~n14549 & n16175 ) ;
  assign n16184 = n16175 | n16183 ;
  assign n16185 = ( n7192 & n14559 ) | ( n7192 & n16175 ) | ( n14559 & n16175 ) ;
  assign n16186 = n16184 | n16185 ;
  assign n16187 = n7196 & ~n15452 ;
  assign n16188 = n16186 & ~n16187 ;
  assign n16189 = n16188 ^ n16187 ^ x23 ;
  assign n16190 = n16189 ^ n16180 ^ n16030 ;
  assign n16191 = ( n16030 & n16180 ) | ( n16030 & n16189 ) | ( n16180 & n16189 ) ;
  assign n16192 = n7339 & n14559 ;
  assign n16193 = ( n7337 & n14569 ) | ( n7337 & n16192 ) | ( n14569 & n16192 ) ;
  assign n16194 = n16192 | n16193 ;
  assign n16195 = ( n7338 & ~n14549 ) | ( n7338 & n16192 ) | ( ~n14549 & n16192 ) ;
  assign n16196 = n16194 | n16195 ;
  assign n16197 = n7340 & ~n15452 ;
  assign n16198 = n16196 & ~n16197 ;
  assign n16199 = n16198 ^ n16197 ^ x20 ;
  assign n16200 = ( n15971 & n16161 ) | ( n15971 & n16199 ) | ( n16161 & n16199 ) ;
  assign n16201 = n16199 ^ n16161 ^ n15971 ;
  assign n16202 = n7037 & n14569 ;
  assign n16203 = ( n7036 & n14559 ) | ( n7036 & n16202 ) | ( n14559 & n16202 ) ;
  assign n16204 = n16202 | n16203 ;
  assign n16205 = ( n7052 & ~n14549 ) | ( n7052 & n16202 ) | ( ~n14549 & n16202 ) ;
  assign n16206 = n16204 | n16205 ;
  assign n16207 = n7035 & ~n15452 ;
  assign n16208 = n16206 | n16207 ;
  assign n16209 = n16208 ^ x26 ^ 1'b0 ;
  assign n16210 = n16209 ^ n16151 ^ n15821 ;
  assign n16211 = ( n15821 & n16151 ) | ( n15821 & n16209 ) | ( n16151 & n16209 ) ;
  assign n16212 = n7829 & n14559 ;
  assign n16213 = ( n7833 & ~n14549 ) | ( n7833 & n16212 ) | ( ~n14549 & n16212 ) ;
  assign n16214 = n16212 | n16213 ;
  assign n16215 = ( n7834 & n14569 ) | ( n7834 & n16212 ) | ( n14569 & n16212 ) ;
  assign n16216 = n16214 | n16215 ;
  assign n16217 = n7838 & ~n15452 ;
  assign n16218 = n16216 & ~n16217 ;
  assign n16219 = n16218 ^ n16217 ^ x11 ;
  assign n16220 = ( n15914 & n16062 ) | ( n15914 & n16219 ) | ( n16062 & n16219 ) ;
  assign n16221 = n16219 ^ n16062 ^ n15914 ;
  assign n16222 = n7669 & n14559 ;
  assign n16223 = ( n7667 & n14569 ) | ( n7667 & n16222 ) | ( n14569 & n16222 ) ;
  assign n16224 = ( n7674 & ~n14549 ) | ( n7674 & n16222 ) | ( ~n14549 & n16222 ) ;
  assign n16225 = n16222 | n16224 ;
  assign n16226 = n16223 | n16225 ;
  assign n16227 = n7666 & ~n15452 ;
  assign n16228 = n16226 & ~n16227 ;
  assign n16229 = n16228 ^ n16227 ^ x14 ;
  assign n16230 = ( n16079 & n16181 ) | ( n16079 & n16229 ) | ( n16181 & n16229 ) ;
  assign n16231 = n16229 ^ n16181 ^ n16079 ;
  assign n16232 = n7669 & n14569 ;
  assign n16233 = n7037 & n14578 ;
  assign n16234 = n7188 & n14578 ;
  assign n16235 = ( n7192 & n14569 ) | ( n7192 & n16234 ) | ( n14569 & n16234 ) ;
  assign n16236 = ( n7674 & n14559 ) | ( n7674 & n16232 ) | ( n14559 & n16232 ) ;
  assign n16237 = n16232 | n16236 ;
  assign n16238 = ( n7667 & n14578 ) | ( n7667 & n16232 ) | ( n14578 & n16232 ) ;
  assign n16239 = n16237 | n16238 ;
  assign n16240 = n7666 & n15475 ;
  assign n16241 = n16239 | n16240 ;
  assign n16242 = ( n7190 & n14559 ) | ( n7190 & n16234 ) | ( n14559 & n16234 ) ;
  assign n16243 = n16234 | n16242 ;
  assign n16244 = n7339 & n14569 ;
  assign n16245 = n16235 | n16243 ;
  assign n16246 = n16241 ^ x14 ^ 1'b0 ;
  assign n16247 = ( n7337 & n14578 ) | ( n7337 & n16244 ) | ( n14578 & n16244 ) ;
  assign n16248 = n16244 | n16247 ;
  assign n16249 = ( n7338 & n14559 ) | ( n7338 & n16244 ) | ( n14559 & n16244 ) ;
  assign n16250 = n16248 | n16249 ;
  assign n16251 = n7340 & n15475 ;
  assign n16252 = n16250 | n16251 ;
  assign n16253 = ( n7036 & n14569 ) | ( n7036 & n16233 ) | ( n14569 & n16233 ) ;
  assign n16254 = n16233 | n16253 ;
  assign n16255 = ( n7052 & n14559 ) | ( n7052 & n16233 ) | ( n14559 & n16233 ) ;
  assign n16256 = n16252 ^ x20 ^ 1'b0 ;
  assign n16257 = n16254 | n16255 ;
  assign n16258 = ( n16090 & n16230 ) | ( n16090 & n16246 ) | ( n16230 & n16246 ) ;
  assign n16259 = n16246 ^ n16230 ^ n16090 ;
  assign n16260 = n16256 ^ n16200 ^ n15982 ;
  assign n16261 = ( n15982 & n16200 ) | ( n15982 & n16256 ) | ( n16200 & n16256 ) ;
  assign n16262 = n7669 & n14578 ;
  assign n16263 = ( n7674 & n14569 ) | ( n7674 & n16262 ) | ( n14569 & n16262 ) ;
  assign n16264 = n16262 | n16263 ;
  assign n16265 = ( n7667 & n14580 ) | ( n7667 & n16262 ) | ( n14580 & n16262 ) ;
  assign n16266 = n16264 | n16265 ;
  assign n16267 = ( n7035 & n15475 ) | ( n7035 & n16257 ) | ( n15475 & n16257 ) ;
  assign n16268 = n7829 & n14569 ;
  assign n16269 = n16257 | n16267 ;
  assign n16270 = ( n7666 & n15535 ) | ( n7666 & n16266 ) | ( n15535 & n16266 ) ;
  assign n16271 = n16266 | n16270 ;
  assign n16272 = ( n7833 & n14559 ) | ( n7833 & n16268 ) | ( n14559 & n16268 ) ;
  assign n16273 = n16268 | n16272 ;
  assign n16274 = ( n7834 & n14578 ) | ( n7834 & n16268 ) | ( n14578 & n16268 ) ;
  assign n16275 = n7838 & n15475 ;
  assign n16276 = n16271 ^ x14 ^ 1'b0 ;
  assign n16277 = n16269 ^ x26 ^ 1'b0 ;
  assign n16278 = n16273 | n16274 ;
  assign n16279 = n7196 & n15475 ;
  assign n16280 = ( ~n15828 & n16211 ) | ( ~n15828 & n16277 ) | ( n16211 & n16277 ) ;
  assign n16281 = n16277 ^ n16211 ^ n15828 ;
  assign n16282 = n7669 & n14580 ;
  assign n16283 = ( n16100 & n16258 ) | ( n16100 & n16276 ) | ( n16258 & n16276 ) ;
  assign n16284 = n16276 ^ n16258 ^ n16100 ;
  assign n16285 = ( n7674 & n14578 ) | ( n7674 & n16282 ) | ( n14578 & n16282 ) ;
  assign n16286 = n16282 | n16285 ;
  assign n16287 = n16245 | n16279 ;
  assign n16288 = ( n7667 & n14584 ) | ( n7667 & n16282 ) | ( n14584 & n16282 ) ;
  assign n16289 = n16287 ^ x23 ^ 1'b0 ;
  assign n16290 = ( n16040 & n16191 ) | ( n16040 & n16289 ) | ( n16191 & n16289 ) ;
  assign n16291 = n16275 | n16278 ;
  assign n16292 = n7669 & n14584 ;
  assign n16293 = ( n7674 & n14580 ) | ( n7674 & n16292 ) | ( n14580 & n16292 ) ;
  assign n16294 = n16292 | n16293 ;
  assign n16295 = n16291 ^ x11 ^ 1'b0 ;
  assign n16296 = n16286 | n16288 ;
  assign n16297 = ( n7666 & n15583 ) | ( n7666 & n16296 ) | ( n15583 & n16296 ) ;
  assign n16298 = n16296 | n16297 ;
  assign n16299 = n16289 ^ n16191 ^ n16040 ;
  assign n16300 = n16298 ^ x14 ^ 1'b0 ;
  assign n16301 = n7666 & ~n15638 ;
  assign n16302 = ( n16133 & n16220 ) | ( n16133 & n16295 ) | ( n16220 & n16295 ) ;
  assign n16303 = n16300 ^ n16283 ^ n16110 ;
  assign n16304 = ( n16110 & n16283 ) | ( n16110 & n16300 ) | ( n16283 & n16300 ) ;
  assign n16305 = ( n7667 & ~n14583 ) | ( n7667 & n16292 ) | ( ~n14583 & n16292 ) ;
  assign n16306 = n16294 | n16305 ;
  assign n16307 = ~n16301 & n16306 ;
  assign n16308 = n16307 ^ n16301 ^ x14 ;
  assign n16309 = ( n16140 & n16304 ) | ( n16140 & n16308 ) | ( n16304 & n16308 ) ;
  assign n16310 = n16308 ^ n16304 ^ n16140 ;
  assign n16311 = n16295 ^ n16220 ^ n16133 ;
  assign n16312 = n7037 & n14580 ;
  assign n16313 = ( n7036 & n14578 ) | ( n7036 & n16312 ) | ( n14578 & n16312 ) ;
  assign n16314 = n16312 | n16313 ;
  assign n16315 = ( n7052 & n14569 ) | ( n7052 & n16312 ) | ( n14569 & n16312 ) ;
  assign n16316 = n16314 | n16315 ;
  assign n16317 = ( n7035 & n15535 ) | ( n7035 & n16316 ) | ( n15535 & n16316 ) ;
  assign n16318 = n16316 | n16317 ;
  assign n16319 = n16318 ^ x26 ^ 1'b0 ;
  assign n16320 = n16319 ^ n16280 ^ n15831 ;
  assign n16321 = ( ~n15831 & n16280 ) | ( ~n15831 & n16319 ) | ( n16280 & n16319 ) ;
  assign n16322 = n7339 & n14578 ;
  assign n16323 = ( n7337 & n14580 ) | ( n7337 & n16322 ) | ( n14580 & n16322 ) ;
  assign n16324 = n16322 | n16323 ;
  assign n16325 = ( n7338 & n14569 ) | ( n7338 & n16322 ) | ( n14569 & n16322 ) ;
  assign n16326 = n16324 | n16325 ;
  assign n16327 = ( n7340 & n15535 ) | ( n7340 & n16326 ) | ( n15535 & n16326 ) ;
  assign n16328 = n16326 | n16327 ;
  assign n16329 = n16328 ^ x20 ^ 1'b0 ;
  assign n16330 = n16329 ^ n16261 ^ n16178 ;
  assign n16331 = ( n16178 & n16261 ) | ( n16178 & n16329 ) | ( n16261 & n16329 ) ;
  assign n16332 = n7485 & n14578 ;
  assign n16333 = ( n7486 & n14580 ) | ( n7486 & n16332 ) | ( n14580 & n16332 ) ;
  assign n16334 = n16332 | n16333 ;
  assign n16335 = ( n7493 & n14569 ) | ( n7493 & n16332 ) | ( n14569 & n16332 ) ;
  assign n16336 = n16334 | n16335 ;
  assign n16337 = ( n7487 & n15535 ) | ( n7487 & n16336 ) | ( n15535 & n16336 ) ;
  assign n16338 = n16336 | n16337 ;
  assign n16339 = n16338 ^ x17 ^ 1'b0 ;
  assign n16340 = n16339 ^ n16160 ^ n16141 ;
  assign n16341 = ( n16141 & n16160 ) | ( n16141 & n16339 ) | ( n16160 & n16339 ) ;
  assign n16342 = n7829 & n14578 ;
  assign n16343 = ( n7833 & n14569 ) | ( n7833 & n16342 ) | ( n14569 & n16342 ) ;
  assign n16344 = n16342 | n16343 ;
  assign n16345 = ( n7834 & n14580 ) | ( n7834 & n16342 ) | ( n14580 & n16342 ) ;
  assign n16346 = n16344 | n16345 ;
  assign n16347 = ( n7838 & n15535 ) | ( n7838 & n16346 ) | ( n15535 & n16346 ) ;
  assign n16348 = n16346 | n16347 ;
  assign n16349 = n16348 ^ x11 ^ 1'b0 ;
  assign n16350 = n7188 & n14580 ;
  assign n16351 = ( n7190 & n14569 ) | ( n7190 & n16350 ) | ( n14569 & n16350 ) ;
  assign n16352 = n16350 | n16351 ;
  assign n16353 = ( n7192 & n14578 ) | ( n7192 & n16350 ) | ( n14578 & n16350 ) ;
  assign n16354 = n16352 | n16353 ;
  assign n16355 = ( n7196 & n15535 ) | ( n7196 & n16354 ) | ( n15535 & n16354 ) ;
  assign n16356 = n16354 | n16355 ;
  assign n16357 = n16356 ^ x23 ^ 1'b0 ;
  assign n16358 = ( n16150 & n16290 ) | ( n16150 & n16357 ) | ( n16290 & n16357 ) ;
  assign n16359 = n16357 ^ n16290 ^ n16150 ;
  assign n16360 = ( n16182 & n16302 ) | ( n16182 & n16349 ) | ( n16302 & n16349 ) ;
  assign n16361 = n16349 ^ n16302 ^ n16182 ;
  assign n16362 = n7829 & n14580 ;
  assign n16363 = ( n7833 & n14578 ) | ( n7833 & n16362 ) | ( n14578 & n16362 ) ;
  assign n16364 = n16362 | n16363 ;
  assign n16365 = ( n7834 & n14584 ) | ( n7834 & n16362 ) | ( n14584 & n16362 ) ;
  assign n16366 = n16364 | n16365 ;
  assign n16367 = ( n7838 & n15583 ) | ( n7838 & n16366 ) | ( n15583 & n16366 ) ;
  assign n16368 = n16366 | n16367 ;
  assign n16369 = n16368 ^ x11 ^ 1'b0 ;
  assign n16370 = ( n16231 & n16360 ) | ( n16231 & n16369 ) | ( n16360 & n16369 ) ;
  assign n16371 = n16369 ^ n16360 ^ n16231 ;
  assign n16372 = n7339 & n14580 ;
  assign n16373 = ( n7337 & n14584 ) | ( n7337 & n16372 ) | ( n14584 & n16372 ) ;
  assign n16374 = n16372 | n16373 ;
  assign n16375 = ( n7338 & n14578 ) | ( n7338 & n16372 ) | ( n14578 & n16372 ) ;
  assign n16376 = n16374 | n16375 ;
  assign n16377 = ( n7340 & n15583 ) | ( n7340 & n16376 ) | ( n15583 & n16376 ) ;
  assign n16378 = n16376 | n16377 ;
  assign n16379 = n16378 ^ x20 ^ 1'b0 ;
  assign n16380 = n16379 ^ n16331 ^ n16190 ;
  assign n16381 = ( n16190 & n16331 ) | ( n16190 & n16379 ) | ( n16331 & n16379 ) ;
  assign n16382 = n7932 & n14580 ;
  assign n16383 = ( n7943 & n14578 ) | ( n7943 & n16382 ) | ( n14578 & n16382 ) ;
  assign n16384 = n16382 | n16383 ;
  assign n16385 = ( n7929 & n14584 ) | ( n7929 & n16382 ) | ( n14584 & n16382 ) ;
  assign n16386 = n16384 | n16385 ;
  assign n16387 = ( n7930 & n15583 ) | ( n7930 & n16386 ) | ( n15583 & n16386 ) ;
  assign n16388 = n16386 | n16387 ;
  assign n16389 = n16388 ^ x8 ^ 1'b0 ;
  assign n16390 = n16389 ^ n16221 ^ n15924 ;
  assign n16391 = ( n15924 & n16221 ) | ( n15924 & n16389 ) | ( n16221 & n16389 ) ;
  assign n16392 = n7037 & n14584 ;
  assign n16393 = ( n7036 & n14580 ) | ( n7036 & n16392 ) | ( n14580 & n16392 ) ;
  assign n16394 = n16392 | n16393 ;
  assign n16395 = ( n7052 & n14578 ) | ( n7052 & n16392 ) | ( n14578 & n16392 ) ;
  assign n16396 = n16394 | n16395 ;
  assign n16397 = ( n7035 & n15583 ) | ( n7035 & n16396 ) | ( n15583 & n16396 ) ;
  assign n16398 = n16396 | n16397 ;
  assign n16399 = n16398 ^ x26 ^ 1'b0 ;
  assign n16400 = ( n15842 & n16321 ) | ( n15842 & n16399 ) | ( n16321 & n16399 ) ;
  assign n16401 = n16399 ^ n16321 ^ n15842 ;
  assign n16402 = n7485 & n14580 ;
  assign n16403 = ( n7486 & n14584 ) | ( n7486 & n16402 ) | ( n14584 & n16402 ) ;
  assign n16404 = n16402 | n16403 ;
  assign n16405 = ( n7493 & n14578 ) | ( n7493 & n16402 ) | ( n14578 & n16402 ) ;
  assign n16406 = n16404 | n16405 ;
  assign n16407 = ( n7487 & n15583 ) | ( n7487 & n16406 ) | ( n15583 & n16406 ) ;
  assign n16408 = n16406 | n16407 ;
  assign n16409 = n16408 ^ x17 ^ 1'b0 ;
  assign n16410 = n7188 & n14584 ;
  assign n16411 = ( n7190 & n14578 ) | ( n7190 & n16410 ) | ( n14578 & n16410 ) ;
  assign n16412 = n16410 | n16411 ;
  assign n16413 = ( n7192 & n14580 ) | ( n7192 & n16410 ) | ( n14580 & n16410 ) ;
  assign n16414 = n16412 | n16413 ;
  assign n16415 = ( n7196 & n15583 ) | ( n7196 & n16414 ) | ( n15583 & n16414 ) ;
  assign n16416 = n16414 | n16415 ;
  assign n16417 = n16416 ^ x23 ^ 1'b0 ;
  assign n16418 = n7188 & ~n14583 ;
  assign n16419 = ( n7190 & n14580 ) | ( n7190 & n16418 ) | ( n14580 & n16418 ) ;
  assign n16420 = n16418 | n16419 ;
  assign n16421 = ( n7192 & n14584 ) | ( n7192 & n16418 ) | ( n14584 & n16418 ) ;
  assign n16422 = n16420 | n16421 ;
  assign n16423 = n7196 & ~n15638 ;
  assign n16424 = n16422 | n16423 ;
  assign n16425 = n16409 ^ n16341 ^ n16201 ;
  assign n16426 = ( n16201 & n16341 ) | ( n16201 & n16409 ) | ( n16341 & n16409 ) ;
  assign n16427 = n16417 ^ n16358 ^ n16210 ;
  assign n16428 = ( n16210 & n16358 ) | ( n16210 & n16417 ) | ( n16358 & n16417 ) ;
  assign n16429 = n7037 & ~n14583 ;
  assign n16430 = ( n7036 & n14584 ) | ( n7036 & n16429 ) | ( n14584 & n16429 ) ;
  assign n16431 = n16429 | n16430 ;
  assign n16432 = n16424 ^ x23 ^ 1'b0 ;
  assign n16433 = ( n7052 & n14580 ) | ( n7052 & n16429 ) | ( n14580 & n16429 ) ;
  assign n16434 = n16431 | n16433 ;
  assign n16435 = n7829 & n14584 ;
  assign n16436 = ( n7833 & n14580 ) | ( n7833 & n16435 ) | ( n14580 & n16435 ) ;
  assign n16437 = n16435 | n16436 ;
  assign n16438 = ( n7834 & ~n14583 ) | ( n7834 & n16435 ) | ( ~n14583 & n16435 ) ;
  assign n16439 = n16437 | n16438 ;
  assign n16440 = n7838 & ~n15638 ;
  assign n16441 = n16439 & ~n16440 ;
  assign n16442 = n16441 ^ n16440 ^ x11 ;
  assign n16443 = n16432 ^ n16428 ^ n16281 ;
  assign n16444 = ( ~n16281 & n16428 ) | ( ~n16281 & n16432 ) | ( n16428 & n16432 ) ;
  assign n16445 = n7035 & ~n15638 ;
  assign n16446 = ( n16259 & n16370 ) | ( n16259 & n16442 ) | ( n16370 & n16442 ) ;
  assign n16447 = n16442 ^ n16370 ^ n16259 ;
  assign n16448 = n7487 & ~n15638 ;
  assign n16449 = n7485 & n14584 ;
  assign n16450 = n16434 & ~n16445 ;
  assign n16451 = n16450 ^ n16445 ^ x26 ;
  assign n16452 = ( n7486 & ~n14583 ) | ( n7486 & n16449 ) | ( ~n14583 & n16449 ) ;
  assign n16453 = n16449 | n16452 ;
  assign n16454 = ( n7493 & n14580 ) | ( n7493 & n16449 ) | ( n14580 & n16449 ) ;
  assign n16455 = n16453 | n16454 ;
  assign n16456 = n16451 ^ n16400 ^ n15844 ;
  assign n16457 = ( ~n15844 & n16400 ) | ( ~n15844 & n16451 ) | ( n16400 & n16451 ) ;
  assign n16458 = n7932 & n14584 ;
  assign n16459 = ( n7943 & n14580 ) | ( n7943 & n16458 ) | ( n14580 & n16458 ) ;
  assign n16460 = n16458 | n16459 ;
  assign n16461 = ( n7929 & ~n14583 ) | ( n7929 & n16458 ) | ( ~n14583 & n16458 ) ;
  assign n16462 = ~n16448 & n16455 ;
  assign n16463 = n16460 | n16461 ;
  assign n16464 = n7930 & ~n15638 ;
  assign n16465 = n16463 & ~n16464 ;
  assign n16466 = n16465 ^ n16464 ^ x8 ;
  assign n16467 = n16466 ^ n16391 ^ n16311 ;
  assign n16468 = ( n16311 & n16391 ) | ( n16311 & n16466 ) | ( n16391 & n16466 ) ;
  assign n16469 = n7339 & n14584 ;
  assign n16470 = ( n7338 & n14580 ) | ( n7338 & n16469 ) | ( n14580 & n16469 ) ;
  assign n16471 = n7340 & ~n15638 ;
  assign n16472 = ( n7337 & ~n14583 ) | ( n7337 & n16469 ) | ( ~n14583 & n16469 ) ;
  assign n16473 = n16462 ^ n16448 ^ x17 ;
  assign n16474 = n16469 | n16472 ;
  assign n16475 = n16470 | n16474 ;
  assign n16476 = n16473 ^ n16426 ^ n16260 ;
  assign n16477 = ( n16260 & n16426 ) | ( n16260 & n16473 ) | ( n16426 & n16473 ) ;
  assign n16478 = ~n16471 & n16475 ;
  assign n16479 = n16478 ^ n16471 ^ x20 ;
  assign n16480 = ( n16299 & n16381 ) | ( n16299 & n16479 ) | ( n16381 & n16479 ) ;
  assign n16481 = n16479 ^ n16381 ^ n16299 ;
  assign n16482 = n7838 & ~n15674 ;
  assign n16483 = n7829 & ~n14583 ;
  assign n16484 = ( n7833 & n14584 ) | ( n7833 & n16483 ) | ( n14584 & n16483 ) ;
  assign n16485 = n16483 | n16484 ;
  assign n16486 = ( n7834 & n14599 ) | ( n7834 & n16483 ) | ( n14599 & n16483 ) ;
  assign n16487 = n16485 | n16486 ;
  assign n16488 = n16482 | n16487 ;
  assign n16489 = n7485 & ~n14583 ;
  assign n16490 = n16488 ^ x11 ^ 1'b0 ;
  assign n16491 = n16490 ^ n16446 ^ n16284 ;
  assign n16492 = ( n16284 & n16446 ) | ( n16284 & n16490 ) | ( n16446 & n16490 ) ;
  assign n16493 = ( n7493 & n14584 ) | ( n7493 & n16489 ) | ( n14584 & n16489 ) ;
  assign n16494 = ( n7486 & n14599 ) | ( n7486 & n16489 ) | ( n14599 & n16489 ) ;
  assign n16495 = n16489 | n16494 ;
  assign n16496 = n7036 & ~n14583 ;
  assign n16497 = n16493 | n16495 ;
  assign n16498 = ( n7052 & n14584 ) | ( n7052 & n16496 ) | ( n14584 & n16496 ) ;
  assign n16499 = n16496 | n16498 ;
  assign n16500 = n7487 & ~n15674 ;
  assign n16501 = n16497 | n16500 ;
  assign n16502 = ( n7037 & n14599 ) | ( n7037 & n16499 ) | ( n14599 & n16499 ) ;
  assign n16503 = n16499 | n16502 ;
  assign n16504 = ( n7035 & ~n15674 ) | ( n7035 & n16499 ) | ( ~n15674 & n16499 ) ;
  assign n16505 = n16503 | n16504 ;
  assign n16506 = n16501 ^ x17 ^ 1'b0 ;
  assign n16507 = n16505 ^ x26 ^ 1'b0 ;
  assign n16508 = n16507 ^ n16457 ^ n15854 ;
  assign n16509 = ( ~n15854 & n16457 ) | ( ~n15854 & n16507 ) | ( n16457 & n16507 ) ;
  assign n16510 = ( n16330 & n16477 ) | ( n16330 & n16506 ) | ( n16477 & n16506 ) ;
  assign n16511 = n16506 ^ n16477 ^ n16330 ;
  assign n16512 = n7188 & n14599 ;
  assign n16513 = ( n7190 & n14584 ) | ( n7190 & n16512 ) | ( n14584 & n16512 ) ;
  assign n16514 = n16512 | n16513 ;
  assign n16515 = n7196 & ~n15674 ;
  assign n16516 = ( n7192 & ~n14583 ) | ( n7192 & n16512 ) | ( ~n14583 & n16512 ) ;
  assign n16517 = n16514 | n16516 ;
  assign n16518 = n16515 | n16517 ;
  assign n16519 = n7037 & ~n14610 ;
  assign n16520 = n16518 ^ x23 ^ 1'b0 ;
  assign n16521 = n16520 ^ n16444 ^ n16320 ;
  assign n16522 = ( ~n16320 & n16444 ) | ( ~n16320 & n16520 ) | ( n16444 & n16520 ) ;
  assign n16523 = n7339 & ~n14583 ;
  assign n16524 = ( n7337 & n14599 ) | ( n7337 & n16523 ) | ( n14599 & n16523 ) ;
  assign n16525 = n16523 | n16524 ;
  assign n16526 = ( n7338 & n14584 ) | ( n7338 & n16523 ) | ( n14584 & n16523 ) ;
  assign n16527 = n16525 | n16526 ;
  assign n16528 = ( n7036 & n14599 ) | ( n7036 & n16519 ) | ( n14599 & n16519 ) ;
  assign n16529 = n16519 | n16528 ;
  assign n16530 = ( n7052 & ~n14583 ) | ( n7052 & n16519 ) | ( ~n14583 & n16519 ) ;
  assign n16531 = n16529 | n16530 ;
  assign n16532 = n7340 & ~n15674 ;
  assign n16533 = n16527 | n16532 ;
  assign n16534 = n7035 & ~n15724 ;
  assign n16535 = n16531 & ~n16534 ;
  assign n16536 = n16533 ^ x20 ^ 1'b0 ;
  assign n16537 = n16535 ^ n16534 ^ x26 ;
  assign n16538 = ( ~n15865 & n16509 ) | ( ~n15865 & n16537 ) | ( n16509 & n16537 ) ;
  assign n16539 = n16537 ^ n16509 ^ n15865 ;
  assign n16540 = n7932 & ~n14583 ;
  assign n16541 = ( n7943 & n14584 ) | ( n7943 & n16540 ) | ( n14584 & n16540 ) ;
  assign n16542 = n16540 | n16541 ;
  assign n16543 = ( n7929 & n14599 ) | ( n7929 & n16540 ) | ( n14599 & n16540 ) ;
  assign n16544 = n16542 | n16543 ;
  assign n16545 = n7930 & ~n15674 ;
  assign n16546 = n16544 | n16545 ;
  assign n16547 = n16546 ^ x8 ^ 1'b0 ;
  assign n16548 = n16547 ^ n16468 ^ n16361 ;
  assign n16549 = ( n16361 & n16468 ) | ( n16361 & n16547 ) | ( n16468 & n16547 ) ;
  assign n16550 = n7669 & ~n14583 ;
  assign n16551 = ( n7674 & n14584 ) | ( n7674 & n16550 ) | ( n14584 & n16550 ) ;
  assign n16552 = n16536 ^ n16480 ^ n16359 ;
  assign n16553 = n7666 & ~n15674 ;
  assign n16554 = n16550 | n16551 ;
  assign n16555 = ( n7667 & n14599 ) | ( n7667 & n16550 ) | ( n14599 & n16550 ) ;
  assign n16556 = n16554 | n16555 ;
  assign n16557 = n16553 | n16556 ;
  assign n16558 = n16557 ^ x14 ^ 1'b0 ;
  assign n16559 = n16558 ^ n16340 ^ n16309 ;
  assign n16560 = ( n16359 & n16480 ) | ( n16359 & n16536 ) | ( n16480 & n16536 ) ;
  assign n16561 = ( n16309 & n16340 ) | ( n16309 & n16558 ) | ( n16340 & n16558 ) ;
  assign n16562 = n7829 & n14599 ;
  assign n16563 = ( n7834 & ~n14610 ) | ( n7834 & n16562 ) | ( ~n14610 & n16562 ) ;
  assign n16564 = ( n7833 & ~n14583 ) | ( n7833 & n16562 ) | ( ~n14583 & n16562 ) ;
  assign n16565 = n16562 | n16564 ;
  assign n16566 = n16563 | n16565 ;
  assign n16567 = n7838 & ~n15724 ;
  assign n16568 = n16566 | n16567 ;
  assign n16569 = n16568 ^ x11 ^ 1'b0 ;
  assign n16570 = n16569 ^ n16492 ^ n16303 ;
  assign n16571 = ( n16303 & n16492 ) | ( n16303 & n16569 ) | ( n16492 & n16569 ) ;
  assign n16572 = n7188 & ~n14610 ;
  assign n16573 = ( n7190 & ~n14583 ) | ( n7190 & n16572 ) | ( ~n14583 & n16572 ) ;
  assign n16574 = n16572 | n16573 ;
  assign n16575 = ( n7192 & n14599 ) | ( n7192 & n16572 ) | ( n14599 & n16572 ) ;
  assign n16576 = n16574 | n16575 ;
  assign n16577 = n7196 & ~n15724 ;
  assign n16578 = n16576 | n16577 ;
  assign n16579 = n7932 & n14599 ;
  assign n16580 = ( n7943 & ~n14583 ) | ( n7943 & n16579 ) | ( ~n14583 & n16579 ) ;
  assign n16581 = n16579 | n16580 ;
  assign n16582 = ( n7929 & ~n14610 ) | ( n7929 & n16579 ) | ( ~n14610 & n16579 ) ;
  assign n16583 = n16581 | n16582 ;
  assign n16584 = n16578 ^ x23 ^ 1'b0 ;
  assign n16585 = n16584 ^ n16522 ^ n16401 ;
  assign n16586 = ( n16401 & n16522 ) | ( n16401 & n16584 ) | ( n16522 & n16584 ) ;
  assign n16587 = n7669 & n14599 ;
  assign n16588 = ( n7674 & ~n14583 ) | ( n7674 & n16587 ) | ( ~n14583 & n16587 ) ;
  assign n16589 = n16587 | n16588 ;
  assign n16590 = ( n7667 & ~n14610 ) | ( n7667 & n16587 ) | ( ~n14610 & n16587 ) ;
  assign n16591 = n16589 | n16590 ;
  assign n16592 = n7930 & ~n15724 ;
  assign n16593 = n16583 | n16592 ;
  assign n16594 = n16593 ^ x8 ^ 1'b0 ;
  assign n16595 = n16594 ^ n16549 ^ n16371 ;
  assign n16596 = ( n16371 & n16549 ) | ( n16371 & n16594 ) | ( n16549 & n16594 ) ;
  assign n16597 = n7666 & ~n15724 ;
  assign n16598 = n16591 | n16597 ;
  assign n16599 = n7339 & n14599 ;
  assign n16600 = ( n7337 & ~n14610 ) | ( n7337 & n16599 ) | ( ~n14610 & n16599 ) ;
  assign n16601 = n16599 | n16600 ;
  assign n16602 = ( n7338 & ~n14583 ) | ( n7338 & n16599 ) | ( ~n14583 & n16599 ) ;
  assign n16603 = n16601 | n16602 ;
  assign n16604 = n7340 & ~n15724 ;
  assign n16605 = n16603 | n16604 ;
  assign n16606 = n16598 ^ x14 ^ 1'b0 ;
  assign n16607 = n16605 ^ x20 ^ 1'b0 ;
  assign n16608 = ( n16427 & n16560 ) | ( n16427 & n16607 ) | ( n16560 & n16607 ) ;
  assign n16609 = n16607 ^ n16560 ^ n16427 ;
  assign n16610 = n6791 & n14599 ;
  assign n16611 = ( n6788 & ~n14610 ) | ( n6788 & n16610 ) | ( ~n14610 & n16610 ) ;
  assign n16612 = n16610 | n16611 ;
  assign n16613 = ( n6790 & ~n14583 ) | ( n6790 & n16610 ) | ( ~n14583 & n16610 ) ;
  assign n16614 = n16612 | n16613 ;
  assign n16615 = ( n16425 & n16561 ) | ( n16425 & n16606 ) | ( n16561 & n16606 ) ;
  assign n16616 = n16606 ^ n16561 ^ n16425 ;
  assign n16617 = n6789 & ~n15724 ;
  assign n16618 = n7485 & n14599 ;
  assign n16619 = n16614 | n16617 ;
  assign n16620 = ( n7486 & ~n14610 ) | ( n7486 & n16618 ) | ( ~n14610 & n16618 ) ;
  assign n16621 = n16618 | n16620 ;
  assign n16622 = ( n7493 & ~n14583 ) | ( n7493 & n16618 ) | ( ~n14583 & n16618 ) ;
  assign n16623 = n16621 | n16622 ;
  assign n16624 = n7487 & ~n15724 ;
  assign n16625 = n16623 | n16624 ;
  assign n16626 = n16625 ^ x17 ^ 1'b0 ;
  assign n16627 = n16626 ^ n16510 ^ n16380 ;
  assign n16628 = n8034 & ~n15724 ;
  assign n16629 = ( n16380 & n16510 ) | ( n16380 & n16626 ) | ( n16510 & n16626 ) ;
  assign n16630 = n8029 & n14599 ;
  assign n16631 = ( n8033 & ~n14610 ) | ( n8033 & n16630 ) | ( ~n14610 & n16630 ) ;
  assign n16632 = ( n8037 & ~n14583 ) | ( n8037 & n16630 ) | ( ~n14583 & n16630 ) ;
  assign n16633 = n16630 | n16632 ;
  assign n16634 = n16631 | n16633 ;
  assign n16635 = n16628 | n16634 ;
  assign n16636 = n16635 ^ x5 ^ 1'b0 ;
  assign n16637 = ( n15935 & n16390 ) | ( n15935 & n16636 ) | ( n16390 & n16636 ) ;
  assign n16638 = n16636 ^ n16390 ^ n15935 ;
  assign n16639 = n7669 & ~n14610 ;
  assign n16640 = ( n14599 & ~n14610 ) | ( n14599 & n15675 ) | ( ~n14610 & n15675 ) ;
  assign n16641 = ( n7674 & n14599 ) | ( n7674 & n16639 ) | ( n14599 & n16639 ) ;
  assign n16642 = n16640 ^ n14643 ^ n14610 ;
  assign n16643 = n16639 | n16641 ;
  assign n16644 = ( n7667 & ~n14643 ) | ( n7667 & n16639 ) | ( ~n14643 & n16639 ) ;
  assign n16645 = n16643 | n16644 ;
  assign n16646 = n7666 & n16642 ;
  assign n16647 = n16645 | n16646 ;
  assign n16648 = n16647 ^ x14 ^ 1'b0 ;
  assign n16649 = ( n16476 & n16615 ) | ( n16476 & n16648 ) | ( n16615 & n16648 ) ;
  assign n16650 = n16648 ^ n16615 ^ n16476 ;
  assign n16651 = ( n14610 & n14643 ) | ( n14610 & ~n16640 ) | ( n14643 & ~n16640 ) ;
  assign n16652 = n7188 & ~n14643 ;
  assign n16653 = ( n7190 & n14599 ) | ( n7190 & n16652 ) | ( n14599 & n16652 ) ;
  assign n16654 = n16652 | n16653 ;
  assign n16655 = ( n7192 & ~n14610 ) | ( n7192 & n16652 ) | ( ~n14610 & n16652 ) ;
  assign n16656 = n16654 | n16655 ;
  assign n16657 = n7196 & n16642 ;
  assign n16658 = n16656 | n16657 ;
  assign n16659 = n16658 ^ x23 ^ 1'b0 ;
  assign n16660 = ( ~n16456 & n16586 ) | ( ~n16456 & n16659 ) | ( n16586 & n16659 ) ;
  assign n16661 = n16659 ^ n16586 ^ n16456 ;
  assign n16662 = n8086 & n14599 ;
  assign n16663 = ( n8088 & ~n14610 ) | ( n8088 & n16662 ) | ( ~n14610 & n16662 ) ;
  assign n16664 = n16662 | n16663 ;
  assign n16665 = ( n8090 & ~n14643 ) | ( n8090 & n16662 ) | ( ~n14643 & n16662 ) ;
  assign n16666 = n16664 | n16665 ;
  assign n16667 = ~n8089 & n16642 ;
  assign n16668 = ( n16642 & n16666 ) | ( n16642 & ~n16667 ) | ( n16666 & ~n16667 ) ;
  assign n16669 = n8034 & n16642 ;
  assign n16670 = n16668 ^ x2 ^ 1'b0 ;
  assign n16671 = ( n15728 & n15778 ) | ( n15728 & n16670 ) | ( n15778 & n16670 ) ;
  assign n16672 = n8029 & ~n14610 ;
  assign n16673 = ( n8037 & n14599 ) | ( n8037 & n16672 ) | ( n14599 & n16672 ) ;
  assign n16674 = n16672 | n16673 ;
  assign n16675 = ( n8033 & ~n14643 ) | ( n8033 & n16672 ) | ( ~n14643 & n16672 ) ;
  assign n16676 = n16674 | n16675 ;
  assign n16677 = n16669 | n16676 ;
  assign n16678 = n16677 ^ x5 ^ 1'b0 ;
  assign n16679 = n16678 ^ n16637 ^ n16467 ;
  assign n16680 = ( n16467 & n16637 ) | ( n16467 & n16678 ) | ( n16637 & n16678 ) ;
  assign n16681 = n7932 & ~n14610 ;
  assign n16682 = ( n7943 & n14599 ) | ( n7943 & n16681 ) | ( n14599 & n16681 ) ;
  assign n16683 = n16681 | n16682 ;
  assign n16684 = ( n7929 & ~n14643 ) | ( n7929 & n16681 ) | ( ~n14643 & n16681 ) ;
  assign n16685 = n16683 | n16684 ;
  assign n16686 = n8086 & ~n14610 ;
  assign n16687 = n7930 & n16642 ;
  assign n16688 = n16685 | n16687 ;
  assign n16689 = n16688 ^ x8 ^ 1'b0 ;
  assign n16690 = ( n16447 & n16596 ) | ( n16447 & n16689 ) | ( n16596 & n16689 ) ;
  assign n16691 = n16689 ^ n16596 ^ n16447 ;
  assign n16692 = ( n8090 & n14655 ) | ( n8090 & n16686 ) | ( n14655 & n16686 ) ;
  assign n16693 = ( n8088 & ~n14643 ) | ( n8088 & n16686 ) | ( ~n14643 & n16686 ) ;
  assign n16694 = n16686 | n16693 ;
  assign n16695 = n16692 | n16694 ;
  assign n16696 = n16651 ^ n14655 ^ n14643 ;
  assign n16697 = ~n8089 & n16696 ;
  assign n16698 = ( n16695 & n16696 ) | ( n16695 & ~n16697 ) | ( n16696 & ~n16697 ) ;
  assign n16699 = n16698 ^ x2 ^ 1'b0 ;
  assign n16700 = ( n15934 & n16671 ) | ( n15934 & n16699 ) | ( n16671 & n16699 ) ;
  assign n16701 = n7829 & ~n14610 ;
  assign n16702 = n7485 & ~n14610 ;
  assign n16703 = ( n7833 & n14599 ) | ( n7833 & n16701 ) | ( n14599 & n16701 ) ;
  assign n16704 = n16701 | n16703 ;
  assign n16705 = ( n7834 & ~n14643 ) | ( n7834 & n16701 ) | ( ~n14643 & n16701 ) ;
  assign n16706 = n16704 | n16705 ;
  assign n16707 = n7838 & n16642 ;
  assign n16708 = n16706 | n16707 ;
  assign n16709 = n16708 ^ x11 ^ 1'b0 ;
  assign n16710 = ( n14643 & ~n14655 ) | ( n14643 & n16651 ) | ( ~n14655 & n16651 ) ;
  assign n16711 = n16709 ^ n16571 ^ n16310 ;
  assign n16712 = ( n16310 & n16571 ) | ( n16310 & n16709 ) | ( n16571 & n16709 ) ;
  assign n16713 = n7339 & ~n14610 ;
  assign n16714 = ( n7337 & ~n14643 ) | ( n7337 & n16713 ) | ( ~n14643 & n16713 ) ;
  assign n16715 = n16713 | n16714 ;
  assign n16716 = ( n7338 & n14599 ) | ( n7338 & n16713 ) | ( n14599 & n16713 ) ;
  assign n16717 = n16715 | n16716 ;
  assign n16718 = ( n7486 & ~n14643 ) | ( n7486 & n16702 ) | ( ~n14643 & n16702 ) ;
  assign n16719 = n16702 | n16718 ;
  assign n16720 = ( n7493 & n14599 ) | ( n7493 & n16702 ) | ( n14599 & n16702 ) ;
  assign n16721 = n16719 | n16720 ;
  assign n16722 = n7487 & n16642 ;
  assign n16723 = n16721 | n16722 ;
  assign n16724 = ( n7340 & n16642 ) | ( n7340 & n16717 ) | ( n16642 & n16717 ) ;
  assign n16725 = n16717 | n16724 ;
  assign n16726 = n16723 ^ x17 ^ 1'b0 ;
  assign n16727 = ( n16481 & n16629 ) | ( n16481 & n16726 ) | ( n16629 & n16726 ) ;
  assign n16728 = n16725 ^ x20 ^ 1'b0 ;
  assign n16729 = n16726 ^ n16629 ^ n16481 ;
  assign n16730 = n16728 ^ n16608 ^ n16443 ;
  assign n16731 = ( ~n16443 & n16608 ) | ( ~n16443 & n16728 ) | ( n16608 & n16728 ) ;
  assign n16732 = n6901 & ~n14610 ;
  assign n16733 = ( n6906 & n14599 ) | ( n6906 & n16732 ) | ( n14599 & n16732 ) ;
  assign n16734 = n16732 | n16733 ;
  assign n16735 = ( n6907 & ~n14643 ) | ( n6907 & n16732 ) | ( ~n14643 & n16732 ) ;
  assign n16736 = n16734 | n16735 ;
  assign n16737 = ( n6918 & n16642 ) | ( n6918 & n16736 ) | ( n16642 & n16736 ) ;
  assign n16738 = n16736 | n16737 ;
  assign n16739 = n16738 ^ x29 ^ 1'b0 ;
  assign n16740 = ( ~n15688 & n15896 ) | ( ~n15688 & n16739 ) | ( n15896 & n16739 ) ;
  assign n16741 = n16739 ^ n15896 ^ n15688 ;
  assign n16742 = n6901 & ~n14643 ;
  assign n16743 = ( n6906 & ~n14610 ) | ( n6906 & n16742 ) | ( ~n14610 & n16742 ) ;
  assign n16744 = n16742 | n16743 ;
  assign n16745 = ( n6907 & n14655 ) | ( n6907 & n16742 ) | ( n14655 & n16742 ) ;
  assign n16746 = n16744 | n16745 ;
  assign n16747 = ( n6918 & n16696 ) | ( n6918 & n16746 ) | ( n16696 & n16746 ) ;
  assign n16748 = n16746 | n16747 ;
  assign n16749 = n16748 ^ x29 ^ 1'b0 ;
  assign n16750 = ( x2 & ~n6647 ) | ( x2 & n16619 ) | ( ~n6647 & n16619 ) ;
  assign n16751 = n16619 ^ n6647 ^ x2 ;
  assign n16752 = ( ~n15746 & n16740 ) | ( ~n15746 & n16749 ) | ( n16740 & n16749 ) ;
  assign n16753 = n16749 ^ n16740 ^ n15746 ;
  assign n16754 = n7037 & ~n14643 ;
  assign n16755 = ( n7036 & ~n14610 ) | ( n7036 & n16754 ) | ( ~n14610 & n16754 ) ;
  assign n16756 = n16754 | n16755 ;
  assign n16757 = ( n7052 & n14599 ) | ( n7052 & n16754 ) | ( n14599 & n16754 ) ;
  assign n16758 = n16756 | n16757 ;
  assign n16759 = n16750 ^ n6586 ^ x2 ;
  assign n16760 = ( x2 & n6586 ) | ( x2 & n16750 ) | ( n6586 & n16750 ) ;
  assign n16761 = ( n7035 & n16642 ) | ( n7035 & n16758 ) | ( n16642 & n16758 ) ;
  assign n16762 = n16758 | n16761 ;
  assign n16763 = n6789 & ~n16642 ;
  assign n16764 = ( x2 & n6782 ) | ( x2 & n16760 ) | ( n6782 & n16760 ) ;
  assign n16765 = n16760 ^ n6782 ^ x2 ;
  assign n16766 = n16762 ^ x26 ^ 1'b0 ;
  assign n16767 = ( n15875 & n16538 ) | ( n15875 & n16766 ) | ( n16538 & n16766 ) ;
  assign n16768 = n16766 ^ n16538 ^ n15875 ;
  assign n16769 = n6791 & ~n14610 ;
  assign n16770 = ( n6790 & n14599 ) | ( n6790 & n16769 ) | ( n14599 & n16769 ) ;
  assign n16771 = ( n6788 & ~n14643 ) | ( n6788 & n16769 ) | ( ~n14643 & n16769 ) ;
  assign n16772 = n16769 | n16771 ;
  assign n16773 = n16770 | n16772 ;
  assign n16774 = ( n6789 & ~n16763 ) | ( n6789 & n16773 ) | ( ~n16763 & n16773 ) ;
  assign n16775 = n6901 & n14655 ;
  assign n16776 = ( n6906 & ~n14643 ) | ( n6906 & n16775 ) | ( ~n14643 & n16775 ) ;
  assign n16777 = n16775 | n16776 ;
  assign n16778 = ( n6907 & ~n14692 ) | ( n6907 & n16775 ) | ( ~n14692 & n16775 ) ;
  assign n16779 = n16777 | n16778 ;
  assign n16780 = n16710 ^ n14692 ^ n14655 ;
  assign n16781 = ( n6918 & n16779 ) | ( n6918 & n16780 ) | ( n16779 & n16780 ) ;
  assign n16782 = n16779 | n16781 ;
  assign n16783 = n16782 ^ x29 ^ 1'b0 ;
  assign n16784 = ( n15745 & ~n16751 ) | ( n15745 & n16783 ) | ( ~n16751 & n16783 ) ;
  assign n16785 = n16783 ^ n16751 ^ n15745 ;
  assign n16786 = n6791 & ~n14643 ;
  assign n16787 = ( n6788 & n14655 ) | ( n6788 & n16786 ) | ( n14655 & n16786 ) ;
  assign n16788 = n16786 | n16787 ;
  assign n16789 = ( n6790 & ~n14610 ) | ( n6790 & n16786 ) | ( ~n14610 & n16786 ) ;
  assign n16790 = n16788 | n16789 ;
  assign n16791 = n6789 & ~n16696 ;
  assign n16792 = ( n6789 & n16790 ) | ( n6789 & ~n16791 ) | ( n16790 & ~n16791 ) ;
  assign n16793 = ( n16759 & n16774 ) | ( n16759 & n16784 ) | ( n16774 & n16784 ) ;
  assign n16794 = n16784 ^ n16774 ^ n16759 ;
  assign n16795 = n7339 & ~n14643 ;
  assign n16796 = ( n16765 & n16792 ) | ( n16765 & n16793 ) | ( n16792 & n16793 ) ;
  assign n16797 = n16793 ^ n16792 ^ n16765 ;
  assign n16798 = ( n7337 & n14655 ) | ( n7337 & n16795 ) | ( n14655 & n16795 ) ;
  assign n16799 = n16795 | n16798 ;
  assign n16800 = ~n8089 & n16780 ;
  assign n16801 = ( n7338 & ~n14610 ) | ( n7338 & n16795 ) | ( ~n14610 & n16795 ) ;
  assign n16802 = n16799 | n16801 ;
  assign n16803 = ( n7340 & n16696 ) | ( n7340 & n16802 ) | ( n16696 & n16802 ) ;
  assign n16804 = n16802 | n16803 ;
  assign n16805 = n16804 ^ x20 ^ 1'b0 ;
  assign n16806 = n16805 ^ n16731 ^ n16521 ;
  assign n16807 = ( ~n16521 & n16731 ) | ( ~n16521 & n16805 ) | ( n16731 & n16805 ) ;
  assign n16808 = n8086 & ~n14643 ;
  assign n16809 = ( n8088 & n14655 ) | ( n8088 & n16808 ) | ( n14655 & n16808 ) ;
  assign n16810 = n16808 | n16809 ;
  assign n16811 = ( n8090 & ~n14692 ) | ( n8090 & n16808 ) | ( ~n14692 & n16808 ) ;
  assign n16812 = n16810 | n16811 ;
  assign n16813 = ( n16780 & ~n16800 ) | ( n16780 & n16812 ) | ( ~n16800 & n16812 ) ;
  assign n16814 = n16813 ^ x2 ^ 1'b0 ;
  assign n16815 = ( n16638 & n16700 ) | ( n16638 & n16814 ) | ( n16700 & n16814 ) ;
  assign n16816 = n8029 & ~n14643 ;
  assign n16817 = ( n8037 & ~n14610 ) | ( n8037 & n16816 ) | ( ~n14610 & n16816 ) ;
  assign n16818 = n16816 | n16817 ;
  assign n16819 = ( n8033 & n14655 ) | ( n8033 & n16816 ) | ( n14655 & n16816 ) ;
  assign n16820 = n16818 | n16819 ;
  assign n16821 = ( n8034 & n16696 ) | ( n8034 & n16820 ) | ( n16696 & n16820 ) ;
  assign n16822 = n16820 | n16821 ;
  assign n16823 = n16822 ^ x5 ^ 1'b0 ;
  assign n16824 = ( n16548 & n16680 ) | ( n16548 & n16823 ) | ( n16680 & n16823 ) ;
  assign n16825 = n16823 ^ n16680 ^ n16548 ;
  assign n16826 = n7669 & ~n14643 ;
  assign n16827 = ( n7674 & ~n14610 ) | ( n7674 & n16826 ) | ( ~n14610 & n16826 ) ;
  assign n16828 = n16826 | n16827 ;
  assign n16829 = ( n7667 & n14655 ) | ( n7667 & n16826 ) | ( n14655 & n16826 ) ;
  assign n16830 = n16828 | n16829 ;
  assign n16831 = ( n7666 & n16696 ) | ( n7666 & n16830 ) | ( n16696 & n16830 ) ;
  assign n16832 = n16830 | n16831 ;
  assign n16833 = n16832 ^ x14 ^ 1'b0 ;
  assign n16834 = n16833 ^ n16649 ^ n16511 ;
  assign n16835 = ( n16511 & n16649 ) | ( n16511 & n16833 ) | ( n16649 & n16833 ) ;
  assign n16836 = n7932 & ~n14643 ;
  assign n16837 = ( n7943 & ~n14610 ) | ( n7943 & n16836 ) | ( ~n14610 & n16836 ) ;
  assign n16838 = n16836 | n16837 ;
  assign n16839 = ( n7929 & n14655 ) | ( n7929 & n16836 ) | ( n14655 & n16836 ) ;
  assign n16840 = n16838 | n16839 ;
  assign n16841 = ( n7930 & n16696 ) | ( n7930 & n16840 ) | ( n16696 & n16840 ) ;
  assign n16842 = n16840 | n16841 ;
  assign n16843 = n16842 ^ x8 ^ 1'b0 ;
  assign n16844 = n16843 ^ n16690 ^ n16491 ;
  assign n16845 = ( n16491 & n16690 ) | ( n16491 & n16843 ) | ( n16690 & n16843 ) ;
  assign n16846 = n7188 & n14655 ;
  assign n16847 = ( n7190 & ~n14610 ) | ( n7190 & n16846 ) | ( ~n14610 & n16846 ) ;
  assign n16848 = n16846 | n16847 ;
  assign n16849 = ( n7192 & ~n14643 ) | ( n7192 & n16846 ) | ( ~n14643 & n16846 ) ;
  assign n16850 = n16848 | n16849 ;
  assign n16851 = n7196 & n16696 ;
  assign n16852 = n16850 | n16851 ;
  assign n16853 = n16852 ^ x23 ^ 1'b0 ;
  assign n16854 = ( ~n16508 & n16660 ) | ( ~n16508 & n16853 ) | ( n16660 & n16853 ) ;
  assign n16855 = n16853 ^ n16660 ^ n16508 ;
  assign n16856 = n7829 & ~n14643 ;
  assign n16857 = ( n7833 & ~n14610 ) | ( n7833 & n16856 ) | ( ~n14610 & n16856 ) ;
  assign n16858 = n16856 | n16857 ;
  assign n16859 = ( n7834 & n14655 ) | ( n7834 & n16856 ) | ( n14655 & n16856 ) ;
  assign n16860 = n16858 | n16859 ;
  assign n16861 = ( n7838 & n16696 ) | ( n7838 & n16860 ) | ( n16696 & n16860 ) ;
  assign n16862 = n16860 | n16861 ;
  assign n16863 = n16862 ^ x11 ^ 1'b0 ;
  assign n16864 = n16863 ^ n16712 ^ n16559 ;
  assign n16865 = ( n16559 & n16712 ) | ( n16559 & n16863 ) | ( n16712 & n16863 ) ;
  assign n16866 = n7188 & ~n14692 ;
  assign n16867 = ( n7190 & ~n14643 ) | ( n7190 & n16866 ) | ( ~n14643 & n16866 ) ;
  assign n16868 = n16866 | n16867 ;
  assign n16869 = ( n7192 & n14655 ) | ( n7192 & n16866 ) | ( n14655 & n16866 ) ;
  assign n16870 = n16868 | n16869 ;
  assign n16871 = n7196 & n16780 ;
  assign n16872 = n16870 | n16871 ;
  assign n16873 = n16872 ^ x23 ^ 1'b0 ;
  assign n16874 = ( ~n16539 & n16854 ) | ( ~n16539 & n16873 ) | ( n16854 & n16873 ) ;
  assign n16875 = n16873 ^ n16854 ^ n16539 ;
  assign n16876 = n7037 & n14655 ;
  assign n16877 = ( n7036 & ~n14643 ) | ( n7036 & n16876 ) | ( ~n14643 & n16876 ) ;
  assign n16878 = n16876 | n16877 ;
  assign n16879 = ( n7052 & ~n14610 ) | ( n7052 & n16876 ) | ( ~n14610 & n16876 ) ;
  assign n16880 = n16878 | n16879 ;
  assign n16881 = ( n7035 & n16696 ) | ( n7035 & n16880 ) | ( n16696 & n16880 ) ;
  assign n16882 = n16880 | n16881 ;
  assign n16883 = n16882 ^ x26 ^ 1'b0 ;
  assign n16884 = n16883 ^ n16767 ^ n15885 ;
  assign n16885 = ( ~n15885 & n16767 ) | ( ~n15885 & n16883 ) | ( n16767 & n16883 ) ;
  assign n16886 = n7485 & ~n14643 ;
  assign n16887 = ( n7486 & n14655 ) | ( n7486 & n16886 ) | ( n14655 & n16886 ) ;
  assign n16888 = n16886 | n16887 ;
  assign n16889 = ( n7493 & ~n14610 ) | ( n7493 & n16886 ) | ( ~n14610 & n16886 ) ;
  assign n16890 = n16888 | n16889 ;
  assign n16891 = ( n7487 & n16696 ) | ( n7487 & n16890 ) | ( n16696 & n16890 ) ;
  assign n16892 = n16890 | n16891 ;
  assign n16893 = n16892 ^ x17 ^ 1'b0 ;
  assign n16894 = ( n16552 & n16727 ) | ( n16552 & n16893 ) | ( n16727 & n16893 ) ;
  assign n16895 = n16893 ^ n16727 ^ n16552 ;
  assign n16896 = n7485 & n14655 ;
  assign n16897 = ( n7486 & ~n14692 ) | ( n7486 & n16896 ) | ( ~n14692 & n16896 ) ;
  assign n16898 = n16896 | n16897 ;
  assign n16899 = ( n7493 & ~n14643 ) | ( n7493 & n16896 ) | ( ~n14643 & n16896 ) ;
  assign n16900 = n16898 | n16899 ;
  assign n16901 = ( n7487 & n16780 ) | ( n7487 & n16900 ) | ( n16780 & n16900 ) ;
  assign n16902 = n16900 | n16901 ;
  assign n16903 = n16902 ^ x17 ^ 1'b0 ;
  assign n16904 = n16903 ^ n16894 ^ n16609 ;
  assign n16905 = ( n16609 & n16894 ) | ( n16609 & n16903 ) | ( n16894 & n16903 ) ;
  assign n16906 = n8029 & n14655 ;
  assign n16907 = ( n8037 & ~n14643 ) | ( n8037 & n16906 ) | ( ~n14643 & n16906 ) ;
  assign n16908 = n16906 | n16907 ;
  assign n16909 = ( n8033 & ~n14692 ) | ( n8033 & n16906 ) | ( ~n14692 & n16906 ) ;
  assign n16910 = n16908 | n16909 ;
  assign n16911 = ( n8034 & n16780 ) | ( n8034 & n16910 ) | ( n16780 & n16910 ) ;
  assign n16912 = n16910 | n16911 ;
  assign n16913 = n16912 ^ x5 ^ 1'b0 ;
  assign n16914 = n16913 ^ n16824 ^ n16595 ;
  assign n16915 = ( n16595 & n16824 ) | ( n16595 & n16913 ) | ( n16824 & n16913 ) ;
  assign n16916 = n7932 & n14655 ;
  assign n16917 = ( n7943 & ~n14643 ) | ( n7943 & n16916 ) | ( ~n14643 & n16916 ) ;
  assign n16918 = n16916 | n16917 ;
  assign n16919 = ( n7929 & ~n14692 ) | ( n7929 & n16916 ) | ( ~n14692 & n16916 ) ;
  assign n16920 = n16918 | n16919 ;
  assign n16921 = ( n7930 & n16780 ) | ( n7930 & n16920 ) | ( n16780 & n16920 ) ;
  assign n16922 = n16920 | n16921 ;
  assign n16923 = n16922 ^ x8 ^ 1'b0 ;
  assign n16924 = n16923 ^ n16845 ^ n16570 ;
  assign n16925 = ( n16570 & n16845 ) | ( n16570 & n16923 ) | ( n16845 & n16923 ) ;
  assign n16926 = n7339 & n14655 ;
  assign n16927 = ( n7337 & ~n14692 ) | ( n7337 & n16926 ) | ( ~n14692 & n16926 ) ;
  assign n16928 = n16926 | n16927 ;
  assign n16929 = ( n7338 & ~n14643 ) | ( n7338 & n16926 ) | ( ~n14643 & n16926 ) ;
  assign n16930 = n16928 | n16929 ;
  assign n16931 = ( n7340 & n16780 ) | ( n7340 & n16930 ) | ( n16780 & n16930 ) ;
  assign n16932 = n16930 | n16931 ;
  assign n16933 = n16932 ^ x20 ^ 1'b0 ;
  assign n16934 = n16933 ^ n16807 ^ n16585 ;
  assign n16935 = ( n16585 & n16807 ) | ( n16585 & n16933 ) | ( n16807 & n16933 ) ;
  assign n16936 = n7829 & n14655 ;
  assign n16937 = ( n7833 & ~n14643 ) | ( n7833 & n16936 ) | ( ~n14643 & n16936 ) ;
  assign n16938 = n16936 | n16937 ;
  assign n16939 = ( n7834 & ~n14692 ) | ( n7834 & n16936 ) | ( ~n14692 & n16936 ) ;
  assign n16940 = n16938 | n16939 ;
  assign n16941 = ( n7838 & n16780 ) | ( n7838 & n16940 ) | ( n16780 & n16940 ) ;
  assign n16942 = n16940 | n16941 ;
  assign n16943 = n16942 ^ x11 ^ 1'b0 ;
  assign n16944 = n16943 ^ n16865 ^ n16616 ;
  assign n16945 = ( n16616 & n16865 ) | ( n16616 & n16943 ) | ( n16865 & n16943 ) ;
  assign n16946 = n7037 & ~n14692 ;
  assign n16947 = ( n7036 & n14655 ) | ( n7036 & n16946 ) | ( n14655 & n16946 ) ;
  assign n16948 = n16946 | n16947 ;
  assign n16949 = ( n7052 & ~n14643 ) | ( n7052 & n16946 ) | ( ~n14643 & n16946 ) ;
  assign n16950 = n16948 | n16949 ;
  assign n16951 = ( n7035 & n16780 ) | ( n7035 & n16950 ) | ( n16780 & n16950 ) ;
  assign n16952 = n16950 | n16951 ;
  assign n16953 = n16952 ^ x26 ^ 1'b0 ;
  assign n16954 = ( ~n15895 & n16885 ) | ( ~n15895 & n16953 ) | ( n16885 & n16953 ) ;
  assign n16955 = n16953 ^ n16885 ^ n15895 ;
  assign n16956 = n7669 & n14655 ;
  assign n16957 = ( n7674 & ~n14643 ) | ( n7674 & n16956 ) | ( ~n14643 & n16956 ) ;
  assign n16958 = n16956 | n16957 ;
  assign n16959 = ( n7667 & ~n14692 ) | ( n7667 & n16956 ) | ( ~n14692 & n16956 ) ;
  assign n16960 = n16958 | n16959 ;
  assign n16961 = ( n7666 & n16780 ) | ( n7666 & n16960 ) | ( n16780 & n16960 ) ;
  assign n16962 = n16960 | n16961 ;
  assign n16963 = n16962 ^ x14 ^ 1'b0 ;
  assign n16964 = ( n16627 & n16835 ) | ( n16627 & n16963 ) | ( n16835 & n16963 ) ;
  assign n16965 = n16963 ^ n16835 ^ n16627 ;
  assign n16966 = n6791 & n14655 ;
  assign n16967 = ( n6790 & ~n14643 ) | ( n6790 & n16966 ) | ( ~n14643 & n16966 ) ;
  assign n16968 = ( n6788 & ~n14692 ) | ( n6788 & n16966 ) | ( ~n14692 & n16966 ) ;
  assign n16969 = n16966 | n16968 ;
  assign n16970 = n8086 & n14655 ;
  assign n16971 = n16967 | n16969 ;
  assign n16972 = ( n8088 & ~n14692 ) | ( n8088 & n16970 ) | ( ~n14692 & n16970 ) ;
  assign n16973 = n16970 | n16972 ;
  assign n16974 = ( n8090 & ~n14720 ) | ( n8090 & n16970 ) | ( ~n14720 & n16970 ) ;
  assign n16975 = n16973 | n16974 ;
  assign n16976 = ( ~n14655 & n14692 ) | ( ~n14655 & n16710 ) | ( n14692 & n16710 ) ;
  assign n16977 = n16976 ^ n14720 ^ n14692 ;
  assign n16978 = n6789 & ~n16780 ;
  assign n16979 = ( n6789 & n16971 ) | ( n6789 & ~n16978 ) | ( n16971 & ~n16978 ) ;
  assign n16980 = ~n16975 & n16977 ;
  assign n16981 = ( n8089 & n16975 ) | ( n8089 & ~n16980 ) | ( n16975 & ~n16980 ) ;
  assign n16982 = n16981 ^ x2 ^ 1'b0 ;
  assign n16983 = n8029 & ~n14692 ;
  assign n16984 = ( n16679 & n16815 ) | ( n16679 & n16982 ) | ( n16815 & n16982 ) ;
  assign n16985 = n7669 & ~n14692 ;
  assign n16986 = ( n8037 & n14655 ) | ( n8037 & n16983 ) | ( n14655 & n16983 ) ;
  assign n16987 = n16983 | n16986 ;
  assign n16988 = ( n8033 & ~n14720 ) | ( n8033 & n16983 ) | ( ~n14720 & n16983 ) ;
  assign n16989 = n16987 | n16988 ;
  assign n16990 = n8034 & ~n16977 ;
  assign n16991 = n16989 & ~n16990 ;
  assign n16992 = n16991 ^ n16990 ^ x5 ;
  assign n16993 = ( n16691 & n16915 ) | ( n16691 & n16992 ) | ( n16915 & n16992 ) ;
  assign n16994 = n16992 ^ n16915 ^ n16691 ;
  assign n16995 = ( n7667 & ~n14720 ) | ( n7667 & n16985 ) | ( ~n14720 & n16985 ) ;
  assign n16996 = ( n7674 & n14655 ) | ( n7674 & n16985 ) | ( n14655 & n16985 ) ;
  assign n16997 = n16985 | n16996 ;
  assign n16998 = n7485 & ~n14692 ;
  assign n16999 = n16995 | n16997 ;
  assign n17000 = ( n7486 & ~n14720 ) | ( n7486 & n16998 ) | ( ~n14720 & n16998 ) ;
  assign n17001 = n16998 | n17000 ;
  assign n17002 = ( n7493 & n14655 ) | ( n7493 & n16998 ) | ( n14655 & n16998 ) ;
  assign n17003 = n17001 | n17002 ;
  assign n17004 = n7487 & ~n16977 ;
  assign n17005 = n17003 | n17004 ;
  assign n17006 = n7666 & ~n16977 ;
  assign n17007 = n16999 & ~n17006 ;
  assign n17008 = n17007 ^ n17006 ^ x14 ;
  assign n17009 = n17008 ^ n16964 ^ n16729 ;
  assign n17010 = ( n16729 & n16964 ) | ( n16729 & n17008 ) | ( n16964 & n17008 ) ;
  assign n17011 = n7188 & ~n14720 ;
  assign n17012 = ( n7190 & n14655 ) | ( n7190 & n17011 ) | ( n14655 & n17011 ) ;
  assign n17013 = n17011 | n17012 ;
  assign n17014 = ( n7192 & ~n14692 ) | ( n7192 & n17011 ) | ( ~n14692 & n17011 ) ;
  assign n17015 = n17013 | n17014 ;
  assign n17016 = n17005 ^ x17 ^ 1'b0 ;
  assign n17017 = ( ~n16730 & n16905 ) | ( ~n16730 & n17016 ) | ( n16905 & n17016 ) ;
  assign n17018 = n17016 ^ n16905 ^ n16730 ;
  assign n17019 = n7932 & ~n14692 ;
  assign n17020 = n7196 & ~n16977 ;
  assign n17021 = n17015 | n17020 ;
  assign n17022 = ( n7943 & n14655 ) | ( n7943 & n17019 ) | ( n14655 & n17019 ) ;
  assign n17023 = n17019 | n17022 ;
  assign n17024 = ( n7929 & ~n14720 ) | ( n7929 & n17019 ) | ( ~n14720 & n17019 ) ;
  assign n17025 = n17021 ^ x23 ^ 1'b0 ;
  assign n17026 = n17023 | n17024 ;
  assign n17027 = n7930 & ~n16977 ;
  assign n17028 = n17026 & ~n17027 ;
  assign n17029 = n17028 ^ n17027 ^ x8 ;
  assign n17030 = ( n16711 & n16925 ) | ( n16711 & n17029 ) | ( n16925 & n17029 ) ;
  assign n17031 = n17029 ^ n16925 ^ n16711 ;
  assign n17032 = n7339 & ~n14692 ;
  assign n17033 = ( n7337 & ~n14720 ) | ( n7337 & n17032 ) | ( ~n14720 & n17032 ) ;
  assign n17034 = n17032 | n17033 ;
  assign n17035 = ( n7338 & n14655 ) | ( n7338 & n17032 ) | ( n14655 & n17032 ) ;
  assign n17036 = n17034 | n17035 ;
  assign n17037 = n7340 & ~n16977 ;
  assign n17038 = n17036 & ~n17037 ;
  assign n17039 = n17038 ^ n17037 ^ x20 ;
  assign n17040 = n17039 ^ n16935 ^ n16661 ;
  assign n17041 = ( ~n16661 & n16935 ) | ( ~n16661 & n17039 ) | ( n16935 & n17039 ) ;
  assign n17042 = ( n16768 & n16874 ) | ( n16768 & n17025 ) | ( n16874 & n17025 ) ;
  assign n17043 = n17025 ^ n16874 ^ n16768 ;
  assign n17044 = ( n14692 & n14720 ) | ( n14692 & n16976 ) | ( n14720 & n16976 ) ;
  assign n17045 = n7037 & ~n14720 ;
  assign n17046 = ( n7036 & ~n14692 ) | ( n7036 & n17045 ) | ( ~n14692 & n17045 ) ;
  assign n17047 = n17045 | n17046 ;
  assign n17048 = ( n7052 & n14655 ) | ( n7052 & n17045 ) | ( n14655 & n17045 ) ;
  assign n17049 = n17047 | n17048 ;
  assign n17050 = n7035 & ~n16977 ;
  assign n17051 = n17049 & ~n17050 ;
  assign n17052 = n17051 ^ n17050 ^ x26 ;
  assign n17053 = n17052 ^ n16954 ^ n16741 ;
  assign n17054 = ( ~n16741 & n16954 ) | ( ~n16741 & n17052 ) | ( n16954 & n17052 ) ;
  assign n17055 = n7339 & ~n14720 ;
  assign n17056 = ( n7337 & ~n14770 ) | ( n7337 & n17055 ) | ( ~n14770 & n17055 ) ;
  assign n17057 = n17044 ^ n14770 ^ n14720 ;
  assign n17058 = n17055 | n17056 ;
  assign n17059 = ( n7338 & ~n14692 ) | ( n7338 & n17055 ) | ( ~n14692 & n17055 ) ;
  assign n17060 = n17058 | n17059 ;
  assign n17061 = n7340 & ~n17057 ;
  assign n17062 = n17060 & ~n17061 ;
  assign n17063 = n17062 ^ n17061 ^ x20 ;
  assign n17064 = n17063 ^ n17041 ^ n16855 ;
  assign n17065 = ( ~n16855 & n17041 ) | ( ~n16855 & n17063 ) | ( n17041 & n17063 ) ;
  assign n17066 = n7829 & ~n14692 ;
  assign n17067 = ( n7833 & n14655 ) | ( n7833 & n17066 ) | ( n14655 & n17066 ) ;
  assign n17068 = n17066 | n17067 ;
  assign n17069 = ( n7834 & ~n14720 ) | ( n7834 & n17066 ) | ( ~n14720 & n17066 ) ;
  assign n17070 = n17068 | n17069 ;
  assign n17071 = n7838 & ~n16977 ;
  assign n17072 = n17070 & ~n17071 ;
  assign n17073 = n17072 ^ n17071 ^ x11 ;
  assign n17074 = n17073 ^ n16945 ^ n16650 ;
  assign n17075 = ( n16650 & n16945 ) | ( n16650 & n17073 ) | ( n16945 & n17073 ) ;
  assign n17076 = n8086 & ~n14692 ;
  assign n17077 = ( n8088 & ~n14720 ) | ( n8088 & n17076 ) | ( ~n14720 & n17076 ) ;
  assign n17078 = n17076 | n17077 ;
  assign n17079 = ( n8090 & ~n14770 ) | ( n8090 & n17076 ) | ( ~n14770 & n17076 ) ;
  assign n17080 = n17078 | n17079 ;
  assign n17081 = n17057 & ~n17080 ;
  assign n17082 = ( n8089 & n17080 ) | ( n8089 & ~n17081 ) | ( n17080 & ~n17081 ) ;
  assign n17083 = n17082 ^ x2 ^ 1'b0 ;
  assign n17084 = n6901 & ~n14692 ;
  assign n17085 = ( n16825 & n16984 ) | ( n16825 & n17083 ) | ( n16984 & n17083 ) ;
  assign n17086 = ( n6906 & n14655 ) | ( n6906 & n17084 ) | ( n14655 & n17084 ) ;
  assign n17087 = ( n6907 & ~n14720 ) | ( n6907 & n17084 ) | ( ~n14720 & n17084 ) ;
  assign n17088 = n17084 | n17086 ;
  assign n17089 = n6791 & ~n14692 ;
  assign n17090 = n17087 | n17088 ;
  assign n17091 = ( n6788 & ~n14720 ) | ( n6788 & n17089 ) | ( ~n14720 & n17089 ) ;
  assign n17092 = ( n6790 & n14655 ) | ( n6790 & n17089 ) | ( n14655 & n17089 ) ;
  assign n17093 = n17089 | n17091 ;
  assign n17094 = n17092 | n17093 ;
  assign n17095 = n8029 & ~n14720 ;
  assign n17096 = n6789 & ~n16977 ;
  assign n17097 = n17094 | n17096 ;
  assign n17098 = ( n8033 & ~n14770 ) | ( n8033 & n17095 ) | ( ~n14770 & n17095 ) ;
  assign n17099 = n6918 & ~n16977 ;
  assign n17100 = n17090 | n17099 ;
  assign n17101 = ( n8037 & ~n14692 ) | ( n8037 & n17095 ) | ( ~n14692 & n17095 ) ;
  assign n17102 = n17095 | n17101 ;
  assign n17103 = n17098 | n17102 ;
  assign n17104 = n8034 & ~n17057 ;
  assign n17105 = n17103 | n17104 ;
  assign n17106 = n17105 ^ x5 ^ 1'b0 ;
  assign n17107 = ( n16844 & n16993 ) | ( n16844 & n17106 ) | ( n16993 & n17106 ) ;
  assign n17108 = n17106 ^ n16993 ^ n16844 ;
  assign n17109 = n6588 ^ x5 ^ x2 ;
  assign n17110 = n17109 ^ n16979 ^ n16764 ;
  assign n17111 = ( n16764 & n16979 ) | ( n16764 & n17109 ) | ( n16979 & n17109 ) ;
  assign n17112 = n8086 & ~n14720 ;
  assign n17113 = ( n8090 & ~n14781 ) | ( n8090 & n17112 ) | ( ~n14781 & n17112 ) ;
  assign n17114 = ( n8088 & ~n14770 ) | ( n8088 & n17112 ) | ( ~n14770 & n17112 ) ;
  assign n17115 = n17112 | n17114 ;
  assign n17116 = n17113 | n17115 ;
  assign n17117 = ( n14720 & n14770 ) | ( n14720 & n17044 ) | ( n14770 & n17044 ) ;
  assign n17118 = n17117 ^ n14781 ^ n14770 ;
  assign n17119 = ~n17116 & n17118 ;
  assign n17120 = ( n8089 & n17116 ) | ( n8089 & ~n17119 ) | ( n17116 & ~n17119 ) ;
  assign n17121 = n17120 ^ x2 ^ 1'b0 ;
  assign n17122 = ( n16914 & n17085 ) | ( n16914 & n17121 ) | ( n17085 & n17121 ) ;
  assign n17123 = ( n14770 & n14781 ) | ( n14770 & n17117 ) | ( n14781 & n17117 ) ;
  assign n17124 = n17123 ^ n14814 ^ n14781 ;
  assign n17125 = n6901 & ~n14781 ;
  assign n17126 = ( n6906 & ~n14770 ) | ( n6906 & n17125 ) | ( ~n14770 & n17125 ) ;
  assign n17127 = n17125 | n17126 ;
  assign n17128 = ( n6907 & ~n14814 ) | ( n6907 & n17125 ) | ( ~n14814 & n17125 ) ;
  assign n17129 = ( x2 & x5 ) | ( x2 & ~n6588 ) | ( x5 & ~n6588 ) ;
  assign n17130 = n17127 | n17128 ;
  assign n17131 = ( n6648 & ~n17097 ) | ( n6648 & n17129 ) | ( ~n17097 & n17129 ) ;
  assign n17132 = n17129 ^ n17097 ^ n6648 ;
  assign n17133 = n6918 & ~n17124 ;
  assign n17134 = n17130 & ~n17133 ;
  assign n17135 = n17134 ^ n17133 ^ x29 ;
  assign n17136 = n17135 ^ n17132 ^ n17111 ;
  assign n17137 = ( n17111 & n17132 ) | ( n17111 & n17135 ) | ( n17132 & n17135 ) ;
  assign n17138 = n6791 & ~n14720 ;
  assign n17139 = ( n6788 & ~n14770 ) | ( n6788 & n17138 ) | ( ~n14770 & n17138 ) ;
  assign n17140 = n17138 | n17139 ;
  assign n17141 = ( n6790 & ~n14692 ) | ( n6790 & n17138 ) | ( ~n14692 & n17138 ) ;
  assign n17142 = n17140 | n17141 ;
  assign n17143 = n6789 & ~n17057 ;
  assign n17144 = n17142 | n17143 ;
  assign n17145 = ( n5960 & n6648 ) | ( n5960 & n17131 ) | ( n6648 & n17131 ) ;
  assign n17146 = n17131 ^ n6648 ^ n5960 ;
  assign n17147 = ( n17137 & n17144 ) | ( n17137 & ~n17146 ) | ( n17144 & ~n17146 ) ;
  assign n17148 = n17146 ^ n17144 ^ n17137 ;
  assign n17149 = n7485 & ~n14720 ;
  assign n17150 = ( n7486 & ~n14770 ) | ( n7486 & n17149 ) | ( ~n14770 & n17149 ) ;
  assign n17151 = n17149 | n17150 ;
  assign n17152 = ( n7493 & ~n14692 ) | ( n7493 & n17149 ) | ( ~n14692 & n17149 ) ;
  assign n17153 = n17151 | n17152 ;
  assign n17154 = n7487 & ~n17057 ;
  assign n17155 = n17153 | n17154 ;
  assign n17156 = n17155 ^ x17 ^ 1'b0 ;
  assign n17157 = ( ~n16806 & n17017 ) | ( ~n16806 & n17156 ) | ( n17017 & n17156 ) ;
  assign n17158 = n17156 ^ n17017 ^ n16806 ;
  assign n17159 = n8086 & ~n14770 ;
  assign n17160 = ( n8088 & ~n14781 ) | ( n8088 & n17159 ) | ( ~n14781 & n17159 ) ;
  assign n17161 = n17159 | n17160 ;
  assign n17162 = ( n8090 & ~n14814 ) | ( n8090 & n17159 ) | ( ~n14814 & n17159 ) ;
  assign n17163 = n17161 | n17162 ;
  assign n17164 = n17124 & ~n17163 ;
  assign n17165 = ( n8089 & n17163 ) | ( n8089 & ~n17164 ) | ( n17163 & ~n17164 ) ;
  assign n17166 = n17165 ^ x2 ^ 1'b0 ;
  assign n17167 = ( n16994 & n17122 ) | ( n16994 & n17166 ) | ( n17122 & n17166 ) ;
  assign n17168 = n7669 & ~n14720 ;
  assign n17169 = ( n7667 & ~n14770 ) | ( n7667 & n17168 ) | ( ~n14770 & n17168 ) ;
  assign n17170 = ( n7674 & ~n14692 ) | ( n7674 & n17168 ) | ( ~n14692 & n17168 ) ;
  assign n17171 = n17168 | n17170 ;
  assign n17172 = n7838 & ~n17057 ;
  assign n17173 = n17169 | n17171 ;
  assign n17174 = n7666 & ~n17057 ;
  assign n17175 = n17173 | n17174 ;
  assign n17176 = n17175 ^ x14 ^ 1'b0 ;
  assign n17177 = ( n16895 & n17010 ) | ( n16895 & n17176 ) | ( n17010 & n17176 ) ;
  assign n17178 = n17176 ^ n17010 ^ n16895 ;
  assign n17179 = n7829 & ~n14720 ;
  assign n17180 = ( n7833 & ~n14692 ) | ( n7833 & n17179 ) | ( ~n14692 & n17179 ) ;
  assign n17181 = n17179 | n17180 ;
  assign n17182 = ( n7834 & ~n14770 ) | ( n7834 & n17179 ) | ( ~n14770 & n17179 ) ;
  assign n17183 = n17181 | n17182 ;
  assign n17184 = n7037 & ~n14770 ;
  assign n17185 = n17172 | n17183 ;
  assign n17186 = ( n7036 & ~n14720 ) | ( n7036 & n17184 ) | ( ~n14720 & n17184 ) ;
  assign n17187 = n17185 ^ x11 ^ 1'b0 ;
  assign n17188 = n17187 ^ n17075 ^ n16834 ;
  assign n17189 = ( n16834 & n17075 ) | ( n16834 & n17187 ) | ( n17075 & n17187 ) ;
  assign n17190 = n7188 & ~n14770 ;
  assign n17191 = ( n7190 & ~n14692 ) | ( n7190 & n17190 ) | ( ~n14692 & n17190 ) ;
  assign n17192 = n17190 | n17191 ;
  assign n17193 = ( n7192 & ~n14720 ) | ( n7192 & n17190 ) | ( ~n14720 & n17190 ) ;
  assign n17194 = n17192 | n17193 ;
  assign n17195 = n7196 & ~n17057 ;
  assign n17196 = n17184 | n17186 ;
  assign n17197 = ( n7052 & ~n14692 ) | ( n7052 & n17184 ) | ( ~n14692 & n17184 ) ;
  assign n17198 = n17194 | n17195 ;
  assign n17199 = n17196 | n17197 ;
  assign n17200 = n17198 ^ x23 ^ 1'b0 ;
  assign n17201 = n7339 & ~n14770 ;
  assign n17202 = ( n7337 & ~n14781 ) | ( n7337 & n17201 ) | ( ~n14781 & n17201 ) ;
  assign n17203 = n17201 | n17202 ;
  assign n17204 = ( n7338 & ~n14720 ) | ( n7338 & n17201 ) | ( ~n14720 & n17201 ) ;
  assign n17205 = n17203 | n17204 ;
  assign n17206 = n7035 & ~n17057 ;
  assign n17207 = n17199 & ~n17206 ;
  assign n17208 = n17207 ^ n17206 ^ x26 ;
  assign n17209 = n17200 ^ n17042 ^ n16884 ;
  assign n17210 = ( ~n16884 & n17042 ) | ( ~n16884 & n17200 ) | ( n17042 & n17200 ) ;
  assign n17211 = n7340 & ~n17118 ;
  assign n17212 = n17205 & ~n17211 ;
  assign n17213 = n17212 ^ n17211 ^ x20 ;
  assign n17214 = n17213 ^ n17065 ^ n16875 ;
  assign n17215 = ( ~n16875 & n17065 ) | ( ~n16875 & n17213 ) | ( n17065 & n17213 ) ;
  assign n17216 = n6918 & ~n17057 ;
  assign n17217 = n6901 & ~n14720 ;
  assign n17218 = ( n6906 & ~n14692 ) | ( n6906 & n17217 ) | ( ~n14692 & n17217 ) ;
  assign n17219 = n7930 & ~n17057 ;
  assign n17220 = n17217 | n17218 ;
  assign n17221 = ( n6907 & ~n14770 ) | ( n6907 & n17217 ) | ( ~n14770 & n17217 ) ;
  assign n17222 = n17220 | n17221 ;
  assign n17223 = n17216 | n17222 ;
  assign n17224 = n7932 & ~n14720 ;
  assign n17225 = ( ~n16753 & n17054 ) | ( ~n16753 & n17208 ) | ( n17054 & n17208 ) ;
  assign n17226 = ( n7943 & ~n14692 ) | ( n7943 & n17224 ) | ( ~n14692 & n17224 ) ;
  assign n17227 = n17208 ^ n17054 ^ n16753 ;
  assign n17228 = ( n7929 & ~n14770 ) | ( n7929 & n17224 ) | ( ~n14770 & n17224 ) ;
  assign n17229 = n17224 | n17226 ;
  assign n17230 = n17228 | n17229 ;
  assign n17231 = n17219 | n17230 ;
  assign n17232 = n17231 ^ x8 ^ 1'b0 ;
  assign n17233 = ( n16864 & n17030 ) | ( n16864 & n17232 ) | ( n17030 & n17232 ) ;
  assign n17234 = n17232 ^ n17030 ^ n16864 ;
  assign n17235 = n8029 & ~n14770 ;
  assign n17236 = ( n8037 & ~n14720 ) | ( n8037 & n17235 ) | ( ~n14720 & n17235 ) ;
  assign n17237 = n17235 | n17236 ;
  assign n17238 = ( n8033 & ~n14781 ) | ( n8033 & n17235 ) | ( ~n14781 & n17235 ) ;
  assign n17239 = n17237 | n17238 ;
  assign n17240 = n8034 & ~n17118 ;
  assign n17241 = n17239 | n17240 ;
  assign n17242 = n17241 ^ x5 ^ 1'b0 ;
  assign n17243 = ( n16924 & n17107 ) | ( n16924 & n17242 ) | ( n17107 & n17242 ) ;
  assign n17244 = n17242 ^ n17107 ^ n16924 ;
  assign n17245 = n7669 & ~n14770 ;
  assign n17246 = ( n7674 & ~n14720 ) | ( n7674 & n17245 ) | ( ~n14720 & n17245 ) ;
  assign n17247 = n17245 | n17246 ;
  assign n17248 = ( n7667 & ~n14781 ) | ( n7667 & n17245 ) | ( ~n14781 & n17245 ) ;
  assign n17249 = n17247 | n17248 ;
  assign n17250 = n7666 & ~n17118 ;
  assign n17251 = n17249 | n17250 ;
  assign n17252 = n17251 ^ x14 ^ 1'b0 ;
  assign n17253 = ( n16904 & n17177 ) | ( n16904 & n17252 ) | ( n17177 & n17252 ) ;
  assign n17254 = n17252 ^ n17177 ^ n16904 ;
  assign n17255 = n7188 & ~n14781 ;
  assign n17256 = ( n7190 & ~n14720 ) | ( n7190 & n17255 ) | ( ~n14720 & n17255 ) ;
  assign n17257 = n17255 | n17256 ;
  assign n17258 = ( n7192 & ~n14770 ) | ( n7192 & n17255 ) | ( ~n14770 & n17255 ) ;
  assign n17259 = n17257 | n17258 ;
  assign n17260 = n7196 & ~n17118 ;
  assign n17261 = n17259 | n17260 ;
  assign n17262 = n17261 ^ x23 ^ 1'b0 ;
  assign n17263 = n17262 ^ n17210 ^ n16955 ;
  assign n17264 = ( ~n16955 & n17210 ) | ( ~n16955 & n17262 ) | ( n17210 & n17262 ) ;
  assign n17265 = n7037 & ~n14781 ;
  assign n17266 = ( n7036 & ~n14770 ) | ( n7036 & n17265 ) | ( ~n14770 & n17265 ) ;
  assign n17267 = n17265 | n17266 ;
  assign n17268 = ( n7052 & ~n14720 ) | ( n7052 & n17265 ) | ( ~n14720 & n17265 ) ;
  assign n17269 = n17267 | n17268 ;
  assign n17270 = n7035 & ~n17118 ;
  assign n17271 = n17269 | n17270 ;
  assign n17272 = n17271 ^ x26 ^ 1'b0 ;
  assign n17273 = ( n16752 & ~n16785 ) | ( n16752 & n17272 ) | ( ~n16785 & n17272 ) ;
  assign n17274 = n17272 ^ n16785 ^ n16752 ;
  assign n17275 = n6791 & ~n14770 ;
  assign n17276 = ( n6788 & ~n14781 ) | ( n6788 & n17275 ) | ( ~n14781 & n17275 ) ;
  assign n17277 = n17275 | n17276 ;
  assign n17278 = ( n6790 & ~n14720 ) | ( n6790 & n17275 ) | ( ~n14720 & n17275 ) ;
  assign n17279 = n17277 | n17278 ;
  assign n17280 = n6789 & ~n17118 ;
  assign n17281 = n17279 | n17280 ;
  assign n17282 = ( x8 & n6513 ) | ( x8 & ~n6648 ) | ( n6513 & ~n6648 ) ;
  assign n17283 = n6648 ^ n6513 ^ x8 ;
  assign n17284 = n17283 ^ n17281 ^ n17145 ;
  assign n17285 = ( ~n17145 & n17281 ) | ( ~n17145 & n17283 ) | ( n17281 & n17283 ) ;
  assign n17286 = n6901 & ~n14770 ;
  assign n17287 = ( n6906 & ~n14720 ) | ( n6906 & n17286 ) | ( ~n14720 & n17286 ) ;
  assign n17288 = n17286 | n17287 ;
  assign n17289 = ( n6907 & ~n14781 ) | ( n6907 & n17286 ) | ( ~n14781 & n17286 ) ;
  assign n17290 = n17288 | n17289 ;
  assign n17291 = n6918 & ~n17118 ;
  assign n17292 = n17290 | n17291 ;
  assign n17293 = n17292 ^ x29 ^ 1'b0 ;
  assign n17294 = n17293 ^ n17110 ^ n16796 ;
  assign n17295 = ( n16796 & n17110 ) | ( n16796 & n17293 ) | ( n17110 & n17293 ) ;
  assign n17296 = n7485 & ~n14770 ;
  assign n17297 = ( n7486 & ~n14781 ) | ( n7486 & n17296 ) | ( ~n14781 & n17296 ) ;
  assign n17298 = n17296 | n17297 ;
  assign n17299 = ( n7493 & ~n14720 ) | ( n7493 & n17296 ) | ( ~n14720 & n17296 ) ;
  assign n17300 = n17298 | n17299 ;
  assign n17301 = n7487 & ~n17118 ;
  assign n17302 = n17300 | n17301 ;
  assign n17303 = n17302 ^ x17 ^ 1'b0 ;
  assign n17304 = ( n16934 & n17157 ) | ( n16934 & n17303 ) | ( n17157 & n17303 ) ;
  assign n17305 = n17303 ^ n17157 ^ n16934 ;
  assign n17306 = n7829 & ~n14770 ;
  assign n17307 = ( n7833 & ~n14720 ) | ( n7833 & n17306 ) | ( ~n14720 & n17306 ) ;
  assign n17308 = n17306 | n17307 ;
  assign n17309 = ( n7834 & ~n14781 ) | ( n7834 & n17306 ) | ( ~n14781 & n17306 ) ;
  assign n17310 = n17308 | n17309 ;
  assign n17311 = n7838 & ~n17118 ;
  assign n17312 = n17310 | n17311 ;
  assign n17313 = n7932 & ~n14770 ;
  assign n17314 = ( n7943 & ~n14720 ) | ( n7943 & n17313 ) | ( ~n14720 & n17313 ) ;
  assign n17315 = n17312 ^ x11 ^ 1'b0 ;
  assign n17316 = n17313 | n17314 ;
  assign n17317 = ( n7929 & ~n14781 ) | ( n7929 & n17313 ) | ( ~n14781 & n17313 ) ;
  assign n17318 = n7930 & ~n17118 ;
  assign n17319 = n17316 | n17317 ;
  assign n17320 = n17315 ^ n17189 ^ n16965 ;
  assign n17321 = ( n16965 & n17189 ) | ( n16965 & n17315 ) | ( n17189 & n17315 ) ;
  assign n17322 = n7339 & ~n14781 ;
  assign n17323 = ( n7337 & ~n14814 ) | ( n7337 & n17322 ) | ( ~n14814 & n17322 ) ;
  assign n17324 = n17322 | n17323 ;
  assign n17325 = ( n7338 & ~n14770 ) | ( n7338 & n17322 ) | ( ~n14770 & n17322 ) ;
  assign n17326 = n17324 | n17325 ;
  assign n17327 = n17318 | n17319 ;
  assign n17328 = n17327 ^ x8 ^ 1'b0 ;
  assign n17329 = n7340 & ~n17124 ;
  assign n17330 = n17326 & ~n17329 ;
  assign n17331 = ( n16944 & n17233 ) | ( n16944 & n17328 ) | ( n17233 & n17328 ) ;
  assign n17332 = n17330 ^ n17329 ^ x20 ;
  assign n17333 = n7669 & ~n14781 ;
  assign n17334 = n17328 ^ n17233 ^ n16944 ;
  assign n17335 = n7666 & ~n17124 ;
  assign n17336 = ( n17043 & n17215 ) | ( n17043 & n17332 ) | ( n17215 & n17332 ) ;
  assign n17337 = n17332 ^ n17215 ^ n17043 ;
  assign n17338 = ( n7667 & ~n14814 ) | ( n7667 & n17333 ) | ( ~n14814 & n17333 ) ;
  assign n17339 = ( n7674 & ~n14770 ) | ( n7674 & n17333 ) | ( ~n14770 & n17333 ) ;
  assign n17340 = n17333 | n17339 ;
  assign n17341 = n17338 | n17340 ;
  assign n17342 = ~n17335 & n17341 ;
  assign n17343 = n17342 ^ n17335 ^ x14 ;
  assign n17344 = n17343 ^ n17253 ^ n17018 ;
  assign n17345 = ( ~n17018 & n17253 ) | ( ~n17018 & n17343 ) | ( n17253 & n17343 ) ;
  assign n17346 = n8029 & ~n14781 ;
  assign n17347 = ( n8033 & ~n14814 ) | ( n8033 & n17346 ) | ( ~n14814 & n17346 ) ;
  assign n17348 = ( n8037 & ~n14770 ) | ( n8037 & n17346 ) | ( ~n14770 & n17346 ) ;
  assign n17349 = n17346 | n17348 ;
  assign n17350 = n17347 | n17349 ;
  assign n17351 = n8034 & ~n17124 ;
  assign n17352 = n17350 | n17351 ;
  assign n17353 = n17352 ^ x5 ^ 1'b0 ;
  assign n17354 = ( n17031 & n17243 ) | ( n17031 & n17353 ) | ( n17243 & n17353 ) ;
  assign n17355 = n17353 ^ n17243 ^ n17031 ;
  assign n17356 = n7037 & ~n14814 ;
  assign n17357 = ( n7036 & ~n14781 ) | ( n7036 & n17356 ) | ( ~n14781 & n17356 ) ;
  assign n17358 = n7035 & ~n17124 ;
  assign n17359 = n17356 | n17357 ;
  assign n17360 = n7196 & ~n17124 ;
  assign n17361 = ( n7052 & ~n14770 ) | ( n7052 & n17356 ) | ( ~n14770 & n17356 ) ;
  assign n17362 = n17359 | n17361 ;
  assign n17363 = n7188 & ~n14814 ;
  assign n17364 = n17358 | n17362 ;
  assign n17365 = ( n7190 & ~n14770 ) | ( n7190 & n17363 ) | ( ~n14770 & n17363 ) ;
  assign n17366 = n17363 | n17365 ;
  assign n17367 = ( n7192 & ~n14781 ) | ( n7192 & n17363 ) | ( ~n14781 & n17363 ) ;
  assign n17368 = n17366 | n17367 ;
  assign n17369 = n7829 & ~n14781 ;
  assign n17370 = n17360 | n17368 ;
  assign n17371 = n17364 ^ x26 ^ 1'b0 ;
  assign n17372 = n17370 ^ x23 ^ 1'b0 ;
  assign n17373 = n17100 ^ x29 ^ 1'b0 ;
  assign n17374 = n17372 ^ n17264 ^ n17053 ;
  assign n17375 = ( ~n17053 & n17264 ) | ( ~n17053 & n17372 ) | ( n17264 & n17372 ) ;
  assign n17376 = n7932 & ~n14781 ;
  assign n17377 = ( n7943 & ~n14770 ) | ( n7943 & n17376 ) | ( ~n14770 & n17376 ) ;
  assign n17378 = n17376 | n17377 ;
  assign n17379 = ( n7929 & ~n14814 ) | ( n7929 & n17376 ) | ( ~n14814 & n17376 ) ;
  assign n17380 = n17378 | n17379 ;
  assign n17381 = n7930 & ~n17124 ;
  assign n17382 = n17380 | n17381 ;
  assign n17383 = n17382 ^ x8 ^ 1'b0 ;
  assign n17384 = ( n17074 & n17331 ) | ( n17074 & n17383 ) | ( n17331 & n17383 ) ;
  assign n17385 = n17383 ^ n17331 ^ n17074 ;
  assign n17386 = ( n16794 & n17371 ) | ( n16794 & n17373 ) | ( n17371 & n17373 ) ;
  assign n17387 = n7485 & ~n14781 ;
  assign n17388 = n17373 ^ n17371 ^ n16794 ;
  assign n17389 = ( n7493 & ~n14770 ) | ( n7493 & n17387 ) | ( ~n14770 & n17387 ) ;
  assign n17390 = ( n7486 & ~n14814 ) | ( n7486 & n17387 ) | ( ~n14814 & n17387 ) ;
  assign n17391 = n17387 | n17390 ;
  assign n17392 = n17389 | n17391 ;
  assign n17393 = n7487 & ~n17124 ;
  assign n17394 = n17392 | n17393 ;
  assign n17395 = ( n7833 & ~n14770 ) | ( n7833 & n17369 ) | ( ~n14770 & n17369 ) ;
  assign n17396 = n6791 & ~n14781 ;
  assign n17397 = n17369 | n17395 ;
  assign n17398 = ( n7834 & ~n14814 ) | ( n7834 & n17369 ) | ( ~n14814 & n17369 ) ;
  assign n17399 = ( n6790 & ~n14770 ) | ( n6790 & n17396 ) | ( ~n14770 & n17396 ) ;
  assign n17400 = n17397 | n17398 ;
  assign n17401 = ( n6788 & ~n14814 ) | ( n6788 & n17396 ) | ( ~n14814 & n17396 ) ;
  assign n17402 = n17396 | n17401 ;
  assign n17403 = n7838 & ~n17124 ;
  assign n17404 = n17399 | n17402 ;
  assign n17405 = n6789 & ~n17124 ;
  assign n17406 = n17404 | n17405 ;
  assign n17407 = n17394 ^ x17 ^ 1'b0 ;
  assign n17408 = ( ~n17040 & n17304 ) | ( ~n17040 & n17407 ) | ( n17304 & n17407 ) ;
  assign n17409 = n17400 | n17403 ;
  assign n17410 = n17407 ^ n17304 ^ n17040 ;
  assign n17411 = n17409 ^ x11 ^ 1'b0 ;
  assign n17412 = n17411 ^ n17321 ^ n17009 ;
  assign n17413 = ( n17009 & n17321 ) | ( n17009 & n17411 ) | ( n17321 & n17411 ) ;
  assign n17414 = n8086 & ~n14781 ;
  assign n17415 = ( n8088 & ~n14814 ) | ( n8088 & n17414 ) | ( ~n14814 & n17414 ) ;
  assign n17416 = n17414 | n17415 ;
  assign n17417 = ( n8090 & n14843 ) | ( n8090 & n17414 ) | ( n14843 & n17414 ) ;
  assign n17418 = ( n14781 & n14814 ) | ( n14781 & n17123 ) | ( n14814 & n17123 ) ;
  assign n17419 = ( n14814 & ~n14843 ) | ( n14814 & n17418 ) | ( ~n14843 & n17418 ) ;
  assign n17420 = n17416 | n17417 ;
  assign n17421 = n17418 ^ n14843 ^ n14814 ;
  assign n17422 = ~n8089 & n17421 ;
  assign n17423 = ( n17420 & n17421 ) | ( n17420 & ~n17422 ) | ( n17421 & ~n17422 ) ;
  assign n17424 = n17423 ^ x2 ^ 1'b0 ;
  assign n17425 = n8086 & ~n14814 ;
  assign n17426 = ( n17108 & n17167 ) | ( n17108 & n17424 ) | ( n17167 & n17424 ) ;
  assign n17427 = ( n8090 & n14888 ) | ( n8090 & n17425 ) | ( n14888 & n17425 ) ;
  assign n17428 = ( n8088 & n14843 ) | ( n8088 & n17425 ) | ( n14843 & n17425 ) ;
  assign n17429 = n17425 | n17428 ;
  assign n17430 = n17427 | n17429 ;
  assign n17431 = n17419 ^ n14888 ^ n14843 ;
  assign n17432 = ~n17430 & n17431 ;
  assign n17433 = ( n8089 & n17430 ) | ( n8089 & ~n17432 ) | ( n17430 & ~n17432 ) ;
  assign n17434 = n8029 & n14843 ;
  assign n17435 = n17433 ^ x2 ^ 1'b0 ;
  assign n17436 = ( n17244 & n17426 ) | ( n17244 & n17435 ) | ( n17426 & n17435 ) ;
  assign n17437 = ( n8033 & n14888 ) | ( n8033 & n17434 ) | ( n14888 & n17434 ) ;
  assign n17438 = ( n8037 & ~n14814 ) | ( n8037 & n17434 ) | ( ~n14814 & n17434 ) ;
  assign n17439 = n17434 | n17438 ;
  assign n17440 = n17437 | n17439 ;
  assign n17441 = n8029 & ~n14814 ;
  assign n17442 = ( n8037 & ~n14781 ) | ( n8037 & n17441 ) | ( ~n14781 & n17441 ) ;
  assign n17443 = n17441 | n17442 ;
  assign n17444 = ( n8033 & n14843 ) | ( n8033 & n17441 ) | ( n14843 & n17441 ) ;
  assign n17445 = n17443 | n17444 ;
  assign n17446 = ( n8034 & n17421 ) | ( n8034 & n17445 ) | ( n17421 & n17445 ) ;
  assign n17447 = n17445 | n17446 ;
  assign n17448 = n17447 ^ x5 ^ 1'b0 ;
  assign n17449 = n17448 ^ n17354 ^ n17234 ;
  assign n17450 = ( n17234 & n17354 ) | ( n17234 & n17448 ) | ( n17354 & n17448 ) ;
  assign n17451 = n8034 & ~n17431 ;
  assign n17452 = n17440 & ~n17451 ;
  assign n17453 = n17452 ^ n17451 ^ x5 ;
  assign n17454 = n8086 & n14843 ;
  assign n17455 = ( n17334 & n17450 ) | ( n17334 & n17453 ) | ( n17450 & n17453 ) ;
  assign n17456 = n17453 ^ n17450 ^ n17334 ;
  assign n17457 = ( n8090 & ~n14907 ) | ( n8090 & n17454 ) | ( ~n14907 & n17454 ) ;
  assign n17458 = ( n14843 & n14888 ) | ( n14843 & ~n17419 ) | ( n14888 & ~n17419 ) ;
  assign n17459 = ( n8088 & n14888 ) | ( n8088 & n17454 ) | ( n14888 & n17454 ) ;
  assign n17460 = n17454 | n17459 ;
  assign n17461 = n17458 ^ n14907 ^ n14888 ;
  assign n17462 = n17457 | n17460 ;
  assign n17463 = n17461 & ~n17462 ;
  assign n17464 = ( n8089 & n17462 ) | ( n8089 & ~n17463 ) | ( n17462 & ~n17463 ) ;
  assign n17465 = n17464 ^ x2 ^ 1'b0 ;
  assign n17466 = n8029 & n14888 ;
  assign n17467 = ( n17355 & n17436 ) | ( n17355 & n17465 ) | ( n17436 & n17465 ) ;
  assign n17468 = ( n8033 & ~n14907 ) | ( n8033 & n17466 ) | ( ~n14907 & n17466 ) ;
  assign n17469 = ( n8037 & n14843 ) | ( n8037 & n17466 ) | ( n14843 & n17466 ) ;
  assign n17470 = n17466 | n17469 ;
  assign n17471 = n17468 | n17470 ;
  assign n17472 = n8034 & ~n17461 ;
  assign n17473 = n17471 & ~n17472 ;
  assign n17474 = n17473 ^ n17472 ^ x5 ;
  assign n17475 = ( n17385 & n17455 ) | ( n17385 & n17474 ) | ( n17455 & n17474 ) ;
  assign n17476 = n17474 ^ n17455 ^ n17385 ;
  assign n17477 = n7339 & ~n14814 ;
  assign n17478 = ( n7337 & n14843 ) | ( n7337 & n17477 ) | ( n14843 & n17477 ) ;
  assign n17479 = n17477 | n17478 ;
  assign n17480 = ( n7338 & ~n14781 ) | ( n7338 & n17477 ) | ( ~n14781 & n17477 ) ;
  assign n17481 = n17479 | n17480 ;
  assign n17482 = ( n7340 & n17421 ) | ( n7340 & n17481 ) | ( n17421 & n17481 ) ;
  assign n17483 = n17481 | n17482 ;
  assign n17484 = n17483 ^ x20 ^ 1'b0 ;
  assign n17485 = ( ~n17209 & n17336 ) | ( ~n17209 & n17484 ) | ( n17336 & n17484 ) ;
  assign n17486 = n17484 ^ n17336 ^ n17209 ;
  assign n17487 = n7037 & n14843 ;
  assign n17488 = ( n7036 & ~n14814 ) | ( n7036 & n17487 ) | ( ~n14814 & n17487 ) ;
  assign n17489 = n17487 | n17488 ;
  assign n17490 = ( n7052 & ~n14781 ) | ( n7052 & n17487 ) | ( ~n14781 & n17487 ) ;
  assign n17491 = n17489 | n17490 ;
  assign n17492 = n7035 & n17421 ;
  assign n17493 = n17491 | n17492 ;
  assign n17494 = n17493 ^ x26 ^ 1'b0 ;
  assign n17495 = n17223 ^ x29 ^ 1'b0 ;
  assign n17496 = ( n16797 & n17494 ) | ( n16797 & n17495 ) | ( n17494 & n17495 ) ;
  assign n17497 = n17495 ^ n17494 ^ n16797 ;
  assign n17498 = n7339 & n14843 ;
  assign n17499 = ( n7337 & n14888 ) | ( n7337 & n17498 ) | ( n14888 & n17498 ) ;
  assign n17500 = n17498 | n17499 ;
  assign n17501 = ( n7338 & ~n14814 ) | ( n7338 & n17498 ) | ( ~n14814 & n17498 ) ;
  assign n17502 = n17500 | n17501 ;
  assign n17503 = n7340 & ~n17431 ;
  assign n17504 = n17502 & ~n17503 ;
  assign n17505 = n17504 ^ n17503 ^ x20 ;
  assign n17506 = ( ~n17263 & n17485 ) | ( ~n17263 & n17505 ) | ( n17485 & n17505 ) ;
  assign n17507 = n17505 ^ n17485 ^ n17263 ;
  assign n17508 = n17282 ^ n6783 ^ 1'b0 ;
  assign n17509 = n7037 & n14888 ;
  assign n17510 = n17508 ^ n17406 ^ 1'b0 ;
  assign n17511 = ( n6783 & ~n17282 ) | ( n6783 & n17406 ) | ( ~n17282 & n17406 ) ;
  assign n17512 = ( n7036 & n14843 ) | ( n7036 & n17509 ) | ( n14843 & n17509 ) ;
  assign n17513 = n17509 | n17512 ;
  assign n17514 = ( n7052 & ~n14814 ) | ( n7052 & n17509 ) | ( ~n14814 & n17509 ) ;
  assign n17515 = n17513 | n17514 ;
  assign n17516 = n7035 & ~n17431 ;
  assign n17517 = n17515 | n17516 ;
  assign n17518 = n17517 ^ x26 ^ 1'b0 ;
  assign n17519 = n17518 ^ n17496 ^ n17294 ;
  assign n17520 = ( n17294 & n17496 ) | ( n17294 & n17518 ) | ( n17496 & n17518 ) ;
  assign n17521 = n7188 & n14888 ;
  assign n17522 = ( n7190 & ~n14814 ) | ( n7190 & n17521 ) | ( ~n14814 & n17521 ) ;
  assign n17523 = n17521 | n17522 ;
  assign n17524 = ( n7192 & n14843 ) | ( n7192 & n17521 ) | ( n14843 & n17521 ) ;
  assign n17525 = n17523 | n17524 ;
  assign n17526 = ( n6649 & n6783 ) | ( n6649 & n17511 ) | ( n6783 & n17511 ) ;
  assign n17527 = n17511 ^ n6783 ^ n6649 ;
  assign n17528 = n6783 ^ n6683 ^ x11 ;
  assign n17529 = ( x11 & n6683 ) | ( x11 & n6783 ) | ( n6683 & n6783 ) ;
  assign n17530 = n7196 & ~n17431 ;
  assign n17531 = n17525 | n17530 ;
  assign n17532 = n17531 ^ x23 ^ 1'b0 ;
  assign n17533 = n17532 ^ n17274 ^ n17225 ;
  assign n17534 = ( n17225 & ~n17274 ) | ( n17225 & n17532 ) | ( ~n17274 & n17532 ) ;
  assign n17535 = n6791 & n14843 ;
  assign n17536 = ( n6788 & n14888 ) | ( n6788 & n17535 ) | ( n14888 & n17535 ) ;
  assign n17537 = n17535 | n17536 ;
  assign n17538 = ( n6790 & ~n14814 ) | ( n6790 & n17535 ) | ( ~n14814 & n17535 ) ;
  assign n17539 = n17537 | n17538 ;
  assign n17540 = n6789 & ~n17431 ;
  assign n17541 = n17539 | n17540 ;
  assign n17542 = ( n17526 & ~n17528 ) | ( n17526 & n17541 ) | ( ~n17528 & n17541 ) ;
  assign n17543 = n17541 ^ n17528 ^ n17526 ;
  assign n17544 = n7485 & ~n14814 ;
  assign n17545 = ( n7486 & n14843 ) | ( n7486 & n17544 ) | ( n14843 & n17544 ) ;
  assign n17546 = n17544 | n17545 ;
  assign n17547 = ( n7493 & ~n14781 ) | ( n7493 & n17544 ) | ( ~n14781 & n17544 ) ;
  assign n17548 = n17546 | n17547 ;
  assign n17549 = n7487 & n17421 ;
  assign n17550 = n17548 | n17549 ;
  assign n17551 = n17550 ^ x17 ^ 1'b0 ;
  assign n17552 = n17551 ^ n17408 ^ n17064 ;
  assign n17553 = ( ~n17064 & n17408 ) | ( ~n17064 & n17551 ) | ( n17408 & n17551 ) ;
  assign n17554 = n7932 & ~n14814 ;
  assign n17555 = ( n7943 & ~n14781 ) | ( n7943 & n17554 ) | ( ~n14781 & n17554 ) ;
  assign n17556 = n17554 | n17555 ;
  assign n17557 = ( n7929 & n14843 ) | ( n7929 & n17554 ) | ( n14843 & n17554 ) ;
  assign n17558 = n17556 | n17557 ;
  assign n17559 = ( n7930 & n17421 ) | ( n7930 & n17558 ) | ( n17421 & n17558 ) ;
  assign n17560 = n17558 | n17559 ;
  assign n17561 = n17560 ^ x8 ^ 1'b0 ;
  assign n17562 = n17561 ^ n17384 ^ n17188 ;
  assign n17563 = ( n17188 & n17384 ) | ( n17188 & n17561 ) | ( n17384 & n17561 ) ;
  assign n17564 = n7829 & ~n14814 ;
  assign n17565 = ( n7833 & ~n14781 ) | ( n7833 & n17564 ) | ( ~n14781 & n17564 ) ;
  assign n17566 = n17564 | n17565 ;
  assign n17567 = ( n7834 & n14843 ) | ( n7834 & n17564 ) | ( n14843 & n17564 ) ;
  assign n17568 = n17566 | n17567 ;
  assign n17569 = ( n7838 & n17421 ) | ( n7838 & n17568 ) | ( n17421 & n17568 ) ;
  assign n17570 = n17568 | n17569 ;
  assign n17571 = n17570 ^ x11 ^ 1'b0 ;
  assign n17572 = n17571 ^ n17413 ^ n17178 ;
  assign n17573 = ( n17178 & n17413 ) | ( n17178 & n17571 ) | ( n17413 & n17571 ) ;
  assign n17574 = n7669 & ~n14814 ;
  assign n17575 = ( n7674 & ~n14781 ) | ( n7674 & n17574 ) | ( ~n14781 & n17574 ) ;
  assign n17576 = n17574 | n17575 ;
  assign n17577 = ( n7667 & n14843 ) | ( n7667 & n17574 ) | ( n14843 & n17574 ) ;
  assign n17578 = n17576 | n17577 ;
  assign n17579 = ( n7666 & n17421 ) | ( n7666 & n17578 ) | ( n17421 & n17578 ) ;
  assign n17580 = n17578 | n17579 ;
  assign n17581 = n17580 ^ x14 ^ 1'b0 ;
  assign n17582 = ( ~n17158 & n17345 ) | ( ~n17158 & n17581 ) | ( n17345 & n17581 ) ;
  assign n17583 = n17581 ^ n17345 ^ n17158 ;
  assign n17584 = n7485 & n14843 ;
  assign n17585 = ( n7486 & n14888 ) | ( n7486 & n17584 ) | ( n14888 & n17584 ) ;
  assign n17586 = n17584 | n17585 ;
  assign n17587 = ( n7493 & ~n14814 ) | ( n7493 & n17584 ) | ( ~n14814 & n17584 ) ;
  assign n17588 = n17586 | n17587 ;
  assign n17589 = n7487 & ~n17431 ;
  assign n17590 = n17588 | n17589 ;
  assign n17591 = n17590 ^ x17 ^ 1'b0 ;
  assign n17592 = n17591 ^ n17553 ^ n17214 ;
  assign n17593 = ( ~n17214 & n17553 ) | ( ~n17214 & n17591 ) | ( n17553 & n17591 ) ;
  assign n17594 = n7932 & n14843 ;
  assign n17595 = ( n7943 & ~n14814 ) | ( n7943 & n17594 ) | ( ~n14814 & n17594 ) ;
  assign n17596 = n17594 | n17595 ;
  assign n17597 = ( n7929 & n14888 ) | ( n7929 & n17594 ) | ( n14888 & n17594 ) ;
  assign n17598 = n17596 | n17597 ;
  assign n17599 = n7930 & ~n17431 ;
  assign n17600 = n17598 & ~n17599 ;
  assign n17601 = n17600 ^ n17599 ^ x8 ;
  assign n17602 = n17601 ^ n17563 ^ n17320 ;
  assign n17603 = ( n17320 & n17563 ) | ( n17320 & n17601 ) | ( n17563 & n17601 ) ;
  assign n17604 = n6901 & n14843 ;
  assign n17605 = ( n6906 & ~n14814 ) | ( n6906 & n17604 ) | ( ~n14814 & n17604 ) ;
  assign n17606 = n17604 | n17605 ;
  assign n17607 = ( n6907 & n14888 ) | ( n6907 & n17604 ) | ( n14888 & n17604 ) ;
  assign n17608 = n17606 | n17607 ;
  assign n17609 = n6918 & ~n17431 ;
  assign n17610 = n17608 | n17609 ;
  assign n17611 = n17610 ^ x29 ^ 1'b0 ;
  assign n17612 = n17611 ^ n17284 ^ n17147 ;
  assign n17613 = ( n17147 & ~n17284 ) | ( n17147 & n17611 ) | ( ~n17284 & n17611 ) ;
  assign n17614 = n7666 & ~n17431 ;
  assign n17615 = n7669 & n14843 ;
  assign n17616 = ( n7667 & n14888 ) | ( n7667 & n17615 ) | ( n14888 & n17615 ) ;
  assign n17617 = ( n7674 & ~n14814 ) | ( n7674 & n17615 ) | ( ~n14814 & n17615 ) ;
  assign n17618 = n17615 | n17617 ;
  assign n17619 = n17616 | n17618 ;
  assign n17620 = ~n17614 & n17619 ;
  assign n17621 = n17620 ^ n17614 ^ x14 ;
  assign n17622 = ( n17305 & n17582 ) | ( n17305 & n17621 ) | ( n17582 & n17621 ) ;
  assign n17623 = n17621 ^ n17582 ^ n17305 ;
  assign n17624 = n7838 & ~n17431 ;
  assign n17625 = n7829 & n14843 ;
  assign n17626 = ( n7834 & n14888 ) | ( n7834 & n17625 ) | ( n14888 & n17625 ) ;
  assign n17627 = ( n7833 & ~n14814 ) | ( n7833 & n17625 ) | ( ~n14814 & n17625 ) ;
  assign n17628 = n17625 | n17627 ;
  assign n17629 = n17626 | n17628 ;
  assign n17630 = ~n17624 & n17629 ;
  assign n17631 = n17630 ^ n17624 ^ x11 ;
  assign n17632 = ( n17254 & n17573 ) | ( n17254 & n17631 ) | ( n17573 & n17631 ) ;
  assign n17633 = n17631 ^ n17573 ^ n17254 ;
  assign n17634 = n7487 & ~n17461 ;
  assign n17635 = n7485 & n14888 ;
  assign n17636 = ( n7493 & n14843 ) | ( n7493 & n17635 ) | ( n14843 & n17635 ) ;
  assign n17637 = ( n7486 & ~n14907 ) | ( n7486 & n17635 ) | ( ~n14907 & n17635 ) ;
  assign n17638 = n17635 | n17637 ;
  assign n17639 = n17636 | n17638 ;
  assign n17640 = n17634 | n17639 ;
  assign n17641 = n17640 ^ x17 ^ 1'b0 ;
  assign n17642 = n17641 ^ n17593 ^ n17337 ;
  assign n17643 = ( n17337 & n17593 ) | ( n17337 & n17641 ) | ( n17593 & n17641 ) ;
  assign n17644 = n7196 & n17421 ;
  assign n17645 = n7188 & n14843 ;
  assign n17646 = ( n7192 & ~n14814 ) | ( n7192 & n17645 ) | ( ~n14814 & n17645 ) ;
  assign n17647 = ( n7190 & ~n14781 ) | ( n7190 & n17645 ) | ( ~n14781 & n17645 ) ;
  assign n17648 = n17645 | n17647 ;
  assign n17649 = n17646 | n17648 ;
  assign n17650 = n17644 | n17649 ;
  assign n17651 = n17650 ^ x23 ^ 1'b0 ;
  assign n17652 = n17651 ^ n17375 ^ n17227 ;
  assign n17653 = ( ~n17227 & n17375 ) | ( ~n17227 & n17651 ) | ( n17375 & n17651 ) ;
  assign n17654 = n7196 & ~n17461 ;
  assign n17655 = n7188 & ~n14907 ;
  assign n17656 = ( n7192 & n14888 ) | ( n7192 & n17655 ) | ( n14888 & n17655 ) ;
  assign n17657 = ( n7190 & n14843 ) | ( n7190 & n17655 ) | ( n14843 & n17655 ) ;
  assign n17658 = n17655 | n17657 ;
  assign n17659 = n17656 | n17658 ;
  assign n17660 = n17654 | n17659 ;
  assign n17661 = n17660 ^ x23 ^ 1'b0 ;
  assign n17662 = n17661 ^ n17388 ^ n17273 ;
  assign n17663 = ( n17273 & n17388 ) | ( n17273 & n17661 ) | ( n17388 & n17661 ) ;
  assign n17664 = n6918 & n17421 ;
  assign n17665 = n6901 & ~n14814 ;
  assign n17666 = ( n6907 & n14843 ) | ( n6907 & n17665 ) | ( n14843 & n17665 ) ;
  assign n17667 = ( n6906 & ~n14781 ) | ( n6906 & n17665 ) | ( ~n14781 & n17665 ) ;
  assign n17668 = n17665 | n17667 ;
  assign n17669 = n17666 | n17668 ;
  assign n17670 = n17664 | n17669 ;
  assign n17671 = n6789 & ~n17421 ;
  assign n17672 = n6791 & ~n14814 ;
  assign n17673 = ( n6790 & ~n14781 ) | ( n6790 & n17672 ) | ( ~n14781 & n17672 ) ;
  assign n17674 = ( n6788 & n14843 ) | ( n6788 & n17672 ) | ( n14843 & n17672 ) ;
  assign n17675 = n17672 | n17674 ;
  assign n17676 = n17673 | n17675 ;
  assign n17677 = ( n6789 & ~n17671 ) | ( n6789 & n17676 ) | ( ~n17671 & n17676 ) ;
  assign n17678 = n7037 & ~n14907 ;
  assign n17679 = ( n7036 & n14888 ) | ( n7036 & n17678 ) | ( n14888 & n17678 ) ;
  assign n17680 = n17678 | n17679 ;
  assign n17681 = ( n7052 & n14843 ) | ( n7052 & n17678 ) | ( n14843 & n17678 ) ;
  assign n17682 = n17680 | n17681 ;
  assign n17683 = n7035 & ~n17461 ;
  assign n17684 = n17682 | n17683 ;
  assign n17685 = n17684 ^ x26 ^ 1'b0 ;
  assign n17686 = n17685 ^ n17295 ^ n17136 ;
  assign n17687 = ( n17136 & n17295 ) | ( n17136 & n17685 ) | ( n17295 & n17685 ) ;
  assign n17688 = n7669 & n14888 ;
  assign n17689 = ( n7674 & n14843 ) | ( n7674 & n17688 ) | ( n14843 & n17688 ) ;
  assign n17690 = n17688 | n17689 ;
  assign n17691 = ( n7667 & ~n14907 ) | ( n7667 & n17688 ) | ( ~n14907 & n17688 ) ;
  assign n17692 = n17690 | n17691 ;
  assign n17693 = n7666 & ~n17461 ;
  assign n17694 = n17692 & ~n17693 ;
  assign n17695 = n17694 ^ n17693 ^ x14 ;
  assign n17696 = n17695 ^ n17622 ^ n17410 ;
  assign n17697 = ( ~n17410 & n17622 ) | ( ~n17410 & n17695 ) | ( n17622 & n17695 ) ;
  assign n17698 = n7339 & n14888 ;
  assign n17699 = ( n7337 & ~n14907 ) | ( n7337 & n17698 ) | ( ~n14907 & n17698 ) ;
  assign n17700 = n17698 | n17699 ;
  assign n17701 = ( n7338 & n14843 ) | ( n7338 & n17698 ) | ( n14843 & n17698 ) ;
  assign n17702 = n17700 | n17701 ;
  assign n17703 = n7340 & ~n17461 ;
  assign n17704 = n17702 & ~n17703 ;
  assign n17705 = n17704 ^ n17703 ^ x20 ;
  assign n17706 = n17705 ^ n17506 ^ n17374 ;
  assign n17707 = ( ~n17374 & n17506 ) | ( ~n17374 & n17705 ) | ( n17506 & n17705 ) ;
  assign n17708 = n6901 & n14888 ;
  assign n17709 = ( n6906 & n14843 ) | ( n6906 & n17708 ) | ( n14843 & n17708 ) ;
  assign n17710 = n17708 | n17709 ;
  assign n17711 = ( n6907 & ~n14907 ) | ( n6907 & n17708 ) | ( ~n14907 & n17708 ) ;
  assign n17712 = n17710 | n17711 ;
  assign n17713 = n6918 & ~n17461 ;
  assign n17714 = n17712 & ~n17713 ;
  assign n17715 = n17714 ^ n17713 ^ x29 ;
  assign n17716 = n17715 ^ n17510 ^ n17285 ;
  assign n17717 = ( n17285 & ~n17510 ) | ( n17285 & n17715 ) | ( ~n17510 & n17715 ) ;
  assign n17718 = n7829 & n14888 ;
  assign n17719 = ( n7833 & n14843 ) | ( n7833 & n17718 ) | ( n14843 & n17718 ) ;
  assign n17720 = n17718 | n17719 ;
  assign n17721 = ( n7834 & ~n14907 ) | ( n7834 & n17718 ) | ( ~n14907 & n17718 ) ;
  assign n17722 = n17720 | n17721 ;
  assign n17723 = n7838 & ~n17461 ;
  assign n17724 = n17722 | n17723 ;
  assign n17725 = n17724 ^ x11 ^ 1'b0 ;
  assign n17726 = n17725 ^ n17632 ^ n17344 ;
  assign n17727 = ( ~n17344 & n17632 ) | ( ~n17344 & n17725 ) | ( n17632 & n17725 ) ;
  assign n17728 = n6791 & n14888 ;
  assign n17729 = ( n6788 & ~n14907 ) | ( n6788 & n17728 ) | ( ~n14907 & n17728 ) ;
  assign n17730 = n17728 | n17729 ;
  assign n17731 = ( n6790 & n14843 ) | ( n6790 & n17728 ) | ( n14843 & n17728 ) ;
  assign n17732 = n17730 | n17731 ;
  assign n17733 = n7930 & ~n17461 ;
  assign n17734 = n6789 & ~n17461 ;
  assign n17735 = n17732 | n17734 ;
  assign n17736 = n7932 & n14888 ;
  assign n17737 = ( n7943 & n14843 ) | ( n7943 & n17736 ) | ( n14843 & n17736 ) ;
  assign n17738 = n17736 | n17737 ;
  assign n17739 = ( n7929 & ~n14907 ) | ( n7929 & n17736 ) | ( ~n14907 & n17736 ) ;
  assign n17740 = n17738 | n17739 ;
  assign n17741 = ~n17733 & n17740 ;
  assign n17742 = n17741 ^ n17733 ^ x8 ;
  assign n17743 = ( n17412 & n17603 ) | ( n17412 & n17742 ) | ( n17603 & n17742 ) ;
  assign n17744 = n17742 ^ n17603 ^ n17412 ;
  assign n17745 = n8086 & n14888 ;
  assign n17746 = ( n8090 & n14969 ) | ( n8090 & n17745 ) | ( n14969 & n17745 ) ;
  assign n17747 = ( n14888 & ~n14907 ) | ( n14888 & n17458 ) | ( ~n14907 & n17458 ) ;
  assign n17748 = ( n8088 & ~n14907 ) | ( n8088 & n17745 ) | ( ~n14907 & n17745 ) ;
  assign n17749 = n17745 | n17748 ;
  assign n17750 = n17746 | n17749 ;
  assign n17751 = n17747 ^ n14969 ^ n14907 ;
  assign n17752 = ~n17750 & n17751 ;
  assign n17753 = ( n8089 & n17750 ) | ( n8089 & ~n17752 ) | ( n17750 & ~n17752 ) ;
  assign n17754 = n8086 & ~n14907 ;
  assign n17755 = n17753 ^ x2 ^ 1'b0 ;
  assign n17756 = ( n17449 & n17467 ) | ( n17449 & n17755 ) | ( n17467 & n17755 ) ;
  assign n17757 = ( n8090 & ~n14970 ) | ( n8090 & n17754 ) | ( ~n14970 & n17754 ) ;
  assign n17758 = ( n8088 & n14969 ) | ( n8088 & n17754 ) | ( n14969 & n17754 ) ;
  assign n17759 = n17754 | n17758 ;
  assign n17760 = n17757 | n17759 ;
  assign n17761 = ( ~n14907 & n14969 ) | ( ~n14907 & n17747 ) | ( n14969 & n17747 ) ;
  assign n17762 = n17761 ^ n14970 ^ n14969 ;
  assign n17763 = ~n17760 & n17762 ;
  assign n17764 = ( n8089 & n17760 ) | ( n8089 & ~n17763 ) | ( n17760 & ~n17763 ) ;
  assign n17765 = n17764 ^ x2 ^ 1'b0 ;
  assign n17766 = ( n17456 & n17756 ) | ( n17456 & n17765 ) | ( n17756 & n17765 ) ;
  assign n17767 = ( n14969 & ~n14970 ) | ( n14969 & n17761 ) | ( ~n14970 & n17761 ) ;
  assign n17768 = n8086 & n14969 ;
  assign n17769 = ( n8088 & ~n14970 ) | ( n8088 & n17768 ) | ( ~n14970 & n17768 ) ;
  assign n17770 = n17768 | n17769 ;
  assign n17771 = ( n8090 & n15001 ) | ( n8090 & n17768 ) | ( n15001 & n17768 ) ;
  assign n17772 = n17770 | n17771 ;
  assign n17773 = n17767 ^ n15001 ^ n14970 ;
  assign n17774 = ~n17772 & n17773 ;
  assign n17775 = ( n8089 & n17772 ) | ( n8089 & ~n17774 ) | ( n17772 & ~n17774 ) ;
  assign n17776 = n17775 ^ x2 ^ 1'b0 ;
  assign n17777 = n6901 & ~n14970 ;
  assign n17778 = ( n17476 & n17766 ) | ( n17476 & n17776 ) | ( n17766 & n17776 ) ;
  assign n17779 = ( n6907 & n15001 ) | ( n6907 & n17777 ) | ( n15001 & n17777 ) ;
  assign n17780 = ( n6906 & n14969 ) | ( n6906 & n17777 ) | ( n14969 & n17777 ) ;
  assign n17781 = n17777 | n17780 ;
  assign n17782 = n17779 | n17781 ;
  assign n17783 = n6918 & ~n17773 ;
  assign n17784 = n17529 ^ n6698 ^ 1'b0 ;
  assign n17785 = n17782 & ~n17783 ;
  assign n17786 = n17785 ^ n17783 ^ x29 ;
  assign n17787 = n17784 ^ n17735 ^ 1'b0 ;
  assign n17788 = ( n17542 & n17786 ) | ( n17542 & n17787 ) | ( n17786 & n17787 ) ;
  assign n17789 = n17787 ^ n17786 ^ n17542 ;
  assign n17790 = n6791 & ~n14907 ;
  assign n17791 = ( n6788 & n14969 ) | ( n6788 & n17790 ) | ( n14969 & n17790 ) ;
  assign n17792 = n17790 | n17791 ;
  assign n17793 = ( n6790 & n14888 ) | ( n6790 & n17790 ) | ( n14888 & n17790 ) ;
  assign n17794 = n17792 | n17793 ;
  assign n17795 = n17670 ^ x29 ^ 1'b0 ;
  assign n17796 = n6789 & ~n17751 ;
  assign n17797 = n17794 | n17796 ;
  assign n17798 = ( n6698 & n17529 ) | ( n6698 & ~n17735 ) | ( n17529 & ~n17735 ) ;
  assign n17799 = n17797 ^ n6698 ^ n6670 ;
  assign n17800 = ( n17788 & ~n17798 ) | ( n17788 & n17799 ) | ( ~n17798 & n17799 ) ;
  assign n17801 = n17799 ^ n17798 ^ n17788 ;
  assign n17802 = n7188 & n14969 ;
  assign n17803 = ( n7190 & n14888 ) | ( n7190 & n17802 ) | ( n14888 & n17802 ) ;
  assign n17804 = n17802 | n17803 ;
  assign n17805 = ( n7192 & ~n14907 ) | ( n7192 & n17802 ) | ( ~n14907 & n17802 ) ;
  assign n17806 = n17804 | n17805 ;
  assign n17807 = n6901 & ~n14907 ;
  assign n17808 = ( n6670 & n6698 ) | ( n6670 & ~n17797 ) | ( n6698 & ~n17797 ) ;
  assign n17809 = ( n6906 & n14888 ) | ( n6906 & n17807 ) | ( n14888 & n17807 ) ;
  assign n17810 = n17807 | n17809 ;
  assign n17811 = ( n6907 & n14969 ) | ( n6907 & n17807 ) | ( n14969 & n17807 ) ;
  assign n17812 = n17810 | n17811 ;
  assign n17813 = n6918 & ~n17751 ;
  assign n17814 = n17812 & ~n17813 ;
  assign n17815 = n17814 ^ n17813 ^ x29 ;
  assign n17816 = n17815 ^ n17677 ^ n17527 ;
  assign n17817 = ( n17527 & n17677 ) | ( n17527 & n17815 ) | ( n17677 & n17815 ) ;
  assign n17818 = n7196 & ~n17751 ;
  assign n17819 = n17806 | n17818 ;
  assign n17820 = n17819 ^ x23 ^ 1'b0 ;
  assign n17821 = ( n17386 & n17497 ) | ( n17386 & n17820 ) | ( n17497 & n17820 ) ;
  assign n17822 = n17820 ^ n17497 ^ n17386 ;
  assign n17823 = n7485 & ~n14907 ;
  assign n17824 = ( n7486 & n14969 ) | ( n7486 & n17823 ) | ( n14969 & n17823 ) ;
  assign n17825 = n17823 | n17824 ;
  assign n17826 = ( n7493 & n14888 ) | ( n7493 & n17823 ) | ( n14888 & n17823 ) ;
  assign n17827 = n17825 | n17826 ;
  assign n17828 = n7487 & ~n17751 ;
  assign n17829 = n17827 | n17828 ;
  assign n17830 = n17829 ^ x17 ^ 1'b0 ;
  assign n17831 = ( ~n17486 & n17643 ) | ( ~n17486 & n17830 ) | ( n17643 & n17830 ) ;
  assign n17832 = n17830 ^ n17643 ^ n17486 ;
  assign n17833 = n7339 & ~n14907 ;
  assign n17834 = ( n7337 & n14969 ) | ( n7337 & n17833 ) | ( n14969 & n17833 ) ;
  assign n17835 = n17833 | n17834 ;
  assign n17836 = ( n7338 & n14888 ) | ( n7338 & n17833 ) | ( n14888 & n17833 ) ;
  assign n17837 = n17835 | n17836 ;
  assign n17838 = n7340 & ~n17751 ;
  assign n17839 = n17837 & ~n17838 ;
  assign n17840 = n17839 ^ n17838 ^ x20 ;
  assign n17841 = n17840 ^ n17707 ^ n17652 ;
  assign n17842 = ( ~n17652 & n17707 ) | ( ~n17652 & n17840 ) | ( n17707 & n17840 ) ;
  assign n17843 = n7932 & ~n14907 ;
  assign n17844 = ( n7943 & n14888 ) | ( n7943 & n17843 ) | ( n14888 & n17843 ) ;
  assign n17845 = n17843 | n17844 ;
  assign n17846 = ( n7929 & n14969 ) | ( n7929 & n17843 ) | ( n14969 & n17843 ) ;
  assign n17847 = n17845 | n17846 ;
  assign n17848 = n7930 & ~n17751 ;
  assign n17849 = n17847 | n17848 ;
  assign n17850 = n17849 ^ x8 ^ 1'b0 ;
  assign n17851 = n17850 ^ n17743 ^ n17572 ;
  assign n17852 = ( n17572 & n17743 ) | ( n17572 & n17850 ) | ( n17743 & n17850 ) ;
  assign n17853 = n7829 & ~n14907 ;
  assign n17854 = ( n7833 & n14888 ) | ( n7833 & n17853 ) | ( n14888 & n17853 ) ;
  assign n17855 = n17853 | n17854 ;
  assign n17856 = ( n7834 & n14969 ) | ( n7834 & n17853 ) | ( n14969 & n17853 ) ;
  assign n17857 = n17855 | n17856 ;
  assign n17858 = n7838 & ~n17751 ;
  assign n17859 = n17857 | n17858 ;
  assign n17860 = n17859 ^ x11 ^ 1'b0 ;
  assign n17861 = ( ~n17583 & n17727 ) | ( ~n17583 & n17860 ) | ( n17727 & n17860 ) ;
  assign n17862 = n17860 ^ n17727 ^ n17583 ;
  assign n17863 = n7669 & ~n14907 ;
  assign n17864 = ( n7674 & n14888 ) | ( n7674 & n17863 ) | ( n14888 & n17863 ) ;
  assign n17865 = n17863 | n17864 ;
  assign n17866 = ( n7667 & n14969 ) | ( n7667 & n17863 ) | ( n14969 & n17863 ) ;
  assign n17867 = n17865 | n17866 ;
  assign n17868 = n7666 & ~n17751 ;
  assign n17869 = n17867 & ~n17868 ;
  assign n17870 = n17869 ^ n17868 ^ x14 ;
  assign n17871 = ( ~n17552 & n17697 ) | ( ~n17552 & n17870 ) | ( n17697 & n17870 ) ;
  assign n17872 = n17870 ^ n17697 ^ n17552 ;
  assign n17873 = n7037 & n14969 ;
  assign n17874 = ( n7036 & ~n14907 ) | ( n7036 & n17873 ) | ( ~n14907 & n17873 ) ;
  assign n17875 = n17873 | n17874 ;
  assign n17876 = ( n7052 & n14888 ) | ( n7052 & n17873 ) | ( n14888 & n17873 ) ;
  assign n17877 = n17875 | n17876 ;
  assign n17878 = n7035 & ~n17751 ;
  assign n17879 = n17877 | n17878 ;
  assign n17880 = n8034 & ~n17751 ;
  assign n17881 = n17879 ^ x26 ^ 1'b0 ;
  assign n17882 = n8029 & ~n14907 ;
  assign n17883 = ( n8037 & n14888 ) | ( n8037 & n17882 ) | ( n14888 & n17882 ) ;
  assign n17884 = n17882 | n17883 ;
  assign n17885 = ( n8033 & n14969 ) | ( n8033 & n17882 ) | ( n14969 & n17882 ) ;
  assign n17886 = n17884 | n17885 ;
  assign n17887 = ( ~n17148 & n17795 ) | ( ~n17148 & n17881 ) | ( n17795 & n17881 ) ;
  assign n17888 = n17881 ^ n17795 ^ n17148 ;
  assign n17889 = n17880 | n17886 ;
  assign n17890 = n17889 ^ x5 ^ 1'b0 ;
  assign n17891 = n17890 ^ n17562 ^ n17475 ;
  assign n17892 = ( n17475 & n17562 ) | ( n17475 & n17890 ) | ( n17562 & n17890 ) ;
  assign n17893 = n7037 & ~n14970 ;
  assign n17894 = ( n7036 & n14969 ) | ( n7036 & n17893 ) | ( n14969 & n17893 ) ;
  assign n17895 = n17893 | n17894 ;
  assign n17896 = ( n7052 & ~n14907 ) | ( n7052 & n17893 ) | ( ~n14907 & n17893 ) ;
  assign n17897 = n17895 | n17896 ;
  assign n17898 = n7035 & ~n17762 ;
  assign n17899 = n17897 | n17898 ;
  assign n17900 = n17899 ^ x26 ^ 1'b0 ;
  assign n17901 = ( ~n17612 & n17887 ) | ( ~n17612 & n17900 ) | ( n17887 & n17900 ) ;
  assign n17902 = n17900 ^ n17887 ^ n17612 ;
  assign n17903 = n7932 & n14969 ;
  assign n17904 = ( n7943 & ~n14907 ) | ( n7943 & n17903 ) | ( ~n14907 & n17903 ) ;
  assign n17905 = n17903 | n17904 ;
  assign n17906 = ( n7929 & ~n14970 ) | ( n7929 & n17903 ) | ( ~n14970 & n17903 ) ;
  assign n17907 = n17905 | n17906 ;
  assign n17908 = n7930 & ~n17762 ;
  assign n17909 = n17907 | n17908 ;
  assign n17910 = n17909 ^ x8 ^ 1'b0 ;
  assign n17911 = n17910 ^ n17852 ^ n17633 ;
  assign n17912 = ( n17633 & n17852 ) | ( n17633 & n17910 ) | ( n17852 & n17910 ) ;
  assign n17913 = n7829 & n14969 ;
  assign n17914 = ( n7833 & ~n14907 ) | ( n7833 & n17913 ) | ( ~n14907 & n17913 ) ;
  assign n17915 = n17913 | n17914 ;
  assign n17916 = ( n7834 & ~n14970 ) | ( n7834 & n17913 ) | ( ~n14970 & n17913 ) ;
  assign n17917 = n17915 | n17916 ;
  assign n17918 = n7838 & ~n17762 ;
  assign n17919 = n17917 | n17918 ;
  assign n17920 = n17919 ^ x11 ^ 1'b0 ;
  assign n17921 = n17920 ^ n17861 ^ n17623 ;
  assign n17922 = ( n17623 & n17861 ) | ( n17623 & n17920 ) | ( n17861 & n17920 ) ;
  assign n17923 = n7188 & ~n14970 ;
  assign n17924 = ( n7190 & ~n14907 ) | ( n7190 & n17923 ) | ( ~n14907 & n17923 ) ;
  assign n17925 = n17923 | n17924 ;
  assign n17926 = ( n7192 & n14969 ) | ( n7192 & n17923 ) | ( n14969 & n17923 ) ;
  assign n17927 = n17925 | n17926 ;
  assign n17928 = n7196 & ~n17762 ;
  assign n17929 = n17927 | n17928 ;
  assign n17930 = n17929 ^ x23 ^ 1'b0 ;
  assign n17931 = n17930 ^ n17821 ^ n17519 ;
  assign n17932 = ( n17519 & n17821 ) | ( n17519 & n17930 ) | ( n17821 & n17930 ) ;
  assign n17933 = n8029 & n14969 ;
  assign n17934 = ( n8037 & ~n14907 ) | ( n8037 & n17933 ) | ( ~n14907 & n17933 ) ;
  assign n17935 = n17933 | n17934 ;
  assign n17936 = ( n8033 & ~n14970 ) | ( n8033 & n17933 ) | ( ~n14970 & n17933 ) ;
  assign n17937 = n17935 | n17936 ;
  assign n17938 = n8034 & ~n17762 ;
  assign n17939 = n17937 | n17938 ;
  assign n17940 = n17939 ^ x5 ^ 1'b0 ;
  assign n17941 = n17940 ^ n17892 ^ n17602 ;
  assign n17942 = ( n17602 & n17892 ) | ( n17602 & n17940 ) | ( n17892 & n17940 ) ;
  assign n17943 = n7339 & n14969 ;
  assign n17944 = ( n7337 & ~n14970 ) | ( n7337 & n17943 ) | ( ~n14970 & n17943 ) ;
  assign n17945 = n17943 | n17944 ;
  assign n17946 = ( n7338 & ~n14907 ) | ( n7338 & n17943 ) | ( ~n14907 & n17943 ) ;
  assign n17947 = n17945 | n17946 ;
  assign n17948 = n7340 & ~n17762 ;
  assign n17949 = n17947 | n17948 ;
  assign n17950 = n17949 ^ x20 ^ 1'b0 ;
  assign n17951 = n17950 ^ n17653 ^ n17533 ;
  assign n17952 = ( ~n17533 & n17653 ) | ( ~n17533 & n17950 ) | ( n17653 & n17950 ) ;
  assign n17953 = n7669 & n14969 ;
  assign n17954 = ( n7674 & ~n14907 ) | ( n7674 & n17953 ) | ( ~n14907 & n17953 ) ;
  assign n17955 = n17953 | n17954 ;
  assign n17956 = ( n7667 & ~n14970 ) | ( n7667 & n17953 ) | ( ~n14970 & n17953 ) ;
  assign n17957 = n17955 | n17956 ;
  assign n17958 = n7666 & ~n17762 ;
  assign n17959 = n17957 & ~n17958 ;
  assign n17960 = n17959 ^ n17958 ^ x14 ;
  assign n17961 = ( ~n17592 & n17871 ) | ( ~n17592 & n17960 ) | ( n17871 & n17960 ) ;
  assign n17962 = n17960 ^ n17871 ^ n17592 ;
  assign n17963 = n7485 & n14969 ;
  assign n17964 = ( n7486 & ~n14970 ) | ( n7486 & n17963 ) | ( ~n14970 & n17963 ) ;
  assign n17965 = n17963 | n17964 ;
  assign n17966 = ( n7493 & ~n14907 ) | ( n7493 & n17963 ) | ( ~n14907 & n17963 ) ;
  assign n17967 = n17965 | n17966 ;
  assign n17968 = n7487 & ~n17762 ;
  assign n17969 = n17967 | n17968 ;
  assign n17970 = n17969 ^ x17 ^ 1'b0 ;
  assign n17971 = n17970 ^ n17831 ^ n17507 ;
  assign n17972 = ( ~n17507 & n17831 ) | ( ~n17507 & n17970 ) | ( n17831 & n17970 ) ;
  assign n17973 = n6901 & n14969 ;
  assign n17974 = ( n6906 & ~n14907 ) | ( n6906 & n17973 ) | ( ~n14907 & n17973 ) ;
  assign n17975 = n17973 | n17974 ;
  assign n17976 = ( n6907 & ~n14970 ) | ( n6907 & n17973 ) | ( ~n14970 & n17973 ) ;
  assign n17977 = n17975 | n17976 ;
  assign n17978 = n6918 & ~n17762 ;
  assign n17979 = n17977 | n17978 ;
  assign n17980 = n6791 & n14969 ;
  assign n17981 = ( n6788 & ~n14970 ) | ( n6788 & n17980 ) | ( ~n14970 & n17980 ) ;
  assign n17982 = ( n6790 & ~n14907 ) | ( n6790 & n17980 ) | ( ~n14907 & n17980 ) ;
  assign n17983 = n17980 | n17981 ;
  assign n17984 = n17982 | n17983 ;
  assign n17985 = n8029 & ~n14970 ;
  assign n17986 = ( n8037 & n14969 ) | ( n8037 & n17985 ) | ( n14969 & n17985 ) ;
  assign n17987 = n17985 | n17986 ;
  assign n17988 = ( n8033 & n15001 ) | ( n8033 & n17985 ) | ( n15001 & n17985 ) ;
  assign n17989 = n17987 | n17988 ;
  assign n17990 = n8034 & ~n17773 ;
  assign n17991 = n17989 | n17990 ;
  assign n17992 = n17991 ^ x5 ^ 1'b0 ;
  assign n17993 = ( n17744 & n17942 ) | ( n17744 & n17992 ) | ( n17942 & n17992 ) ;
  assign n17994 = n6789 & ~n17762 ;
  assign n17995 = n17992 ^ n17942 ^ n17744 ;
  assign n17996 = n7829 & ~n14970 ;
  assign n17997 = ( n7833 & n14969 ) | ( n7833 & n17996 ) | ( n14969 & n17996 ) ;
  assign n17998 = n17996 | n17997 ;
  assign n17999 = ( n7834 & n15001 ) | ( n7834 & n17996 ) | ( n15001 & n17996 ) ;
  assign n18000 = n17998 | n17999 ;
  assign n18001 = n7838 & ~n17773 ;
  assign n18002 = n18000 | n18001 ;
  assign n18003 = n6698 ^ n6697 ^ x14 ;
  assign n18004 = n18002 ^ x11 ^ 1'b0 ;
  assign n18005 = n17984 | n17994 ;
  assign n18006 = ( ~n17808 & n18003 ) | ( ~n17808 & n18005 ) | ( n18003 & n18005 ) ;
  assign n18007 = n18005 ^ n18003 ^ n17808 ;
  assign n18008 = n7188 & n15001 ;
  assign n18009 = n17979 ^ x29 ^ 1'b0 ;
  assign n18010 = n18009 ^ n17817 ^ n17543 ;
  assign n18011 = ( ~n17543 & n17817 ) | ( ~n17543 & n18009 ) | ( n17817 & n18009 ) ;
  assign n18012 = ( n7190 & n14969 ) | ( n7190 & n18008 ) | ( n14969 & n18008 ) ;
  assign n18013 = ( n7192 & ~n14970 ) | ( n7192 & n18008 ) | ( ~n14970 & n18008 ) ;
  assign n18014 = n18008 | n18012 ;
  assign n18015 = n7196 & ~n17773 ;
  assign n18016 = ( x14 & n6697 ) | ( x14 & ~n6698 ) | ( n6697 & ~n6698 ) ;
  assign n18017 = n7932 & ~n14970 ;
  assign n18018 = n18013 | n18014 ;
  assign n18019 = n18015 | n18018 ;
  assign n18020 = n18019 ^ x23 ^ 1'b0 ;
  assign n18021 = n18020 ^ n17686 ^ n17520 ;
  assign n18022 = n7669 & ~n14970 ;
  assign n18023 = ( n17520 & n17686 ) | ( n17520 & n18020 ) | ( n17686 & n18020 ) ;
  assign n18024 = ( n7674 & n14969 ) | ( n7674 & n18022 ) | ( n14969 & n18022 ) ;
  assign n18025 = ( n7943 & n14969 ) | ( n7943 & n18017 ) | ( n14969 & n18017 ) ;
  assign n18026 = n18022 | n18024 ;
  assign n18027 = n18017 | n18025 ;
  assign n18028 = ( n7929 & n15001 ) | ( n7929 & n18017 ) | ( n15001 & n18017 ) ;
  assign n18029 = n18027 | n18028 ;
  assign n18030 = n7930 & ~n17773 ;
  assign n18031 = n18029 & ~n18030 ;
  assign n18032 = n18031 ^ n18030 ^ x8 ;
  assign n18033 = ( n7667 & n15001 ) | ( n7667 & n18022 ) | ( n15001 & n18022 ) ;
  assign n18034 = n18026 | n18033 ;
  assign n18035 = n7666 & ~n17773 ;
  assign n18036 = ( ~n17726 & n17912 ) | ( ~n17726 & n18032 ) | ( n17912 & n18032 ) ;
  assign n18037 = n18034 & ~n18035 ;
  assign n18038 = n18037 ^ n18035 ^ x14 ;
  assign n18039 = n18038 ^ n17961 ^ n17642 ;
  assign n18040 = n18032 ^ n17912 ^ n17726 ;
  assign n18041 = ( ~n17696 & n17922 ) | ( ~n17696 & n18004 ) | ( n17922 & n18004 ) ;
  assign n18042 = n18004 ^ n17922 ^ n17696 ;
  assign n18043 = ( n17642 & n17961 ) | ( n17642 & n18038 ) | ( n17961 & n18038 ) ;
  assign n18044 = n7485 & ~n14970 ;
  assign n18045 = ( n7486 & n15001 ) | ( n7486 & n18044 ) | ( n15001 & n18044 ) ;
  assign n18046 = n18044 | n18045 ;
  assign n18047 = ( n7493 & n14969 ) | ( n7493 & n18044 ) | ( n14969 & n18044 ) ;
  assign n18048 = n18046 | n18047 ;
  assign n18049 = n7487 & ~n17773 ;
  assign n18050 = n18048 | n18049 ;
  assign n18051 = n18050 ^ x17 ^ 1'b0 ;
  assign n18052 = ( ~n17706 & n17972 ) | ( ~n17706 & n18051 ) | ( n17972 & n18051 ) ;
  assign n18053 = n18051 ^ n17972 ^ n17706 ;
  assign n18054 = n7037 & n15001 ;
  assign n18055 = ( n7036 & ~n14970 ) | ( n7036 & n18054 ) | ( ~n14970 & n18054 ) ;
  assign n18056 = n18054 | n18055 ;
  assign n18057 = ( n7052 & n14969 ) | ( n7052 & n18054 ) | ( n14969 & n18054 ) ;
  assign n18058 = n18056 | n18057 ;
  assign n18059 = n7035 & ~n17773 ;
  assign n18060 = n18058 | n18059 ;
  assign n18061 = n18060 ^ x26 ^ 1'b0 ;
  assign n18062 = n18061 ^ n17716 ^ n17613 ;
  assign n18063 = ( n17613 & ~n17716 ) | ( n17613 & n18061 ) | ( ~n17716 & n18061 ) ;
  assign n18064 = n7339 & ~n14970 ;
  assign n18065 = ( n7337 & n15001 ) | ( n7337 & n18064 ) | ( n15001 & n18064 ) ;
  assign n18066 = n18064 | n18065 ;
  assign n18067 = ( n7338 & n14969 ) | ( n7338 & n18064 ) | ( n14969 & n18064 ) ;
  assign n18068 = n18066 | n18067 ;
  assign n18069 = n7340 & ~n17773 ;
  assign n18070 = n18068 | n18069 ;
  assign n18071 = n18070 ^ x20 ^ 1'b0 ;
  assign n18072 = ( n17534 & n17662 ) | ( n17534 & n18071 ) | ( n17662 & n18071 ) ;
  assign n18073 = n18071 ^ n17662 ^ n17534 ;
  assign n18074 = n6791 & ~n14970 ;
  assign n18075 = ( n6788 & n15001 ) | ( n6788 & n18074 ) | ( n15001 & n18074 ) ;
  assign n18076 = ( n6790 & n14969 ) | ( n6790 & n18074 ) | ( n14969 & n18074 ) ;
  assign n18077 = n18074 | n18075 ;
  assign n18078 = n8086 & ~n14970 ;
  assign n18079 = n18076 | n18077 ;
  assign n18080 = ( n8088 & n15001 ) | ( n8088 & n18078 ) | ( n15001 & n18078 ) ;
  assign n18081 = n18078 | n18080 ;
  assign n18082 = ( n8090 & ~n15032 ) | ( n8090 & n18078 ) | ( ~n15032 & n18078 ) ;
  assign n18083 = ( ~n14970 & n15001 ) | ( ~n14970 & n17767 ) | ( n15001 & n17767 ) ;
  assign n18084 = n18081 | n18082 ;
  assign n18085 = n18083 ^ n15032 ^ n15001 ;
  assign n18086 = n6789 & ~n17773 ;
  assign n18087 = n18079 | n18086 ;
  assign n18088 = ~n18084 & n18085 ;
  assign n18089 = ( n8089 & n18084 ) | ( n8089 & ~n18088 ) | ( n18084 & ~n18088 ) ;
  assign n18090 = n18089 ^ x2 ^ 1'b0 ;
  assign n18091 = n8034 & ~n18085 ;
  assign n18092 = ( n17778 & n17891 ) | ( n17778 & n18090 ) | ( n17891 & n18090 ) ;
  assign n18093 = n8029 & n15001 ;
  assign n18094 = ( n8037 & ~n14970 ) | ( n8037 & n18093 ) | ( ~n14970 & n18093 ) ;
  assign n18095 = ( n15001 & ~n15032 ) | ( n15001 & n18083 ) | ( ~n15032 & n18083 ) ;
  assign n18096 = n18093 | n18094 ;
  assign n18097 = ( n8033 & ~n15032 ) | ( n8033 & n18093 ) | ( ~n15032 & n18093 ) ;
  assign n18098 = n18096 | n18097 ;
  assign n18099 = n8086 & n15001 ;
  assign n18100 = ~n18091 & n18098 ;
  assign n18101 = n18100 ^ n18091 ^ x5 ;
  assign n18102 = n18101 ^ n17993 ^ n17851 ;
  assign n18103 = ( n17851 & n17993 ) | ( n17851 & n18101 ) | ( n17993 & n18101 ) ;
  assign n18104 = ( n8088 & ~n15032 ) | ( n8088 & n18099 ) | ( ~n15032 & n18099 ) ;
  assign n18105 = n18099 | n18104 ;
  assign n18106 = ( n8090 & ~n15095 ) | ( n8090 & n18099 ) | ( ~n15095 & n18099 ) ;
  assign n18107 = n18105 | n18106 ;
  assign n18108 = n18095 ^ n15095 ^ n15032 ;
  assign n18109 = ~n8089 & n18108 ;
  assign n18110 = ( n18107 & n18108 ) | ( n18107 & ~n18109 ) | ( n18108 & ~n18109 ) ;
  assign n18111 = n18110 ^ x2 ^ 1'b0 ;
  assign n18112 = ( n17941 & n18092 ) | ( n17941 & n18111 ) | ( n18092 & n18111 ) ;
  assign n18113 = n8029 & ~n15032 ;
  assign n18114 = ( n8037 & n15001 ) | ( n8037 & n18113 ) | ( n15001 & n18113 ) ;
  assign n18115 = n18113 | n18114 ;
  assign n18116 = ( n8033 & ~n15095 ) | ( n8033 & n18113 ) | ( ~n15095 & n18113 ) ;
  assign n18117 = n18115 | n18116 ;
  assign n18118 = ( n8034 & n18108 ) | ( n8034 & n18117 ) | ( n18108 & n18117 ) ;
  assign n18119 = n18117 | n18118 ;
  assign n18120 = n18119 ^ x5 ^ 1'b0 ;
  assign n18121 = n18120 ^ n18103 ^ n17911 ;
  assign n18122 = ( n17911 & n18103 ) | ( n17911 & n18120 ) | ( n18103 & n18120 ) ;
  assign n18123 = n7669 & n15001 ;
  assign n18124 = ( n7674 & ~n14970 ) | ( n7674 & n18123 ) | ( ~n14970 & n18123 ) ;
  assign n18125 = n18123 | n18124 ;
  assign n18126 = ( n7667 & ~n15032 ) | ( n7667 & n18123 ) | ( ~n15032 & n18123 ) ;
  assign n18127 = n18125 | n18126 ;
  assign n18128 = n7666 & ~n18085 ;
  assign n18129 = n18127 & ~n18128 ;
  assign n18130 = n18129 ^ n18128 ^ x14 ;
  assign n18131 = ( ~n17832 & n18043 ) | ( ~n17832 & n18130 ) | ( n18043 & n18130 ) ;
  assign n18132 = n18130 ^ n18043 ^ n17832 ;
  assign n18133 = n7829 & n15001 ;
  assign n18134 = ( n7833 & ~n14970 ) | ( n7833 & n18133 ) | ( ~n14970 & n18133 ) ;
  assign n18135 = n18133 | n18134 ;
  assign n18136 = ( n7834 & ~n15032 ) | ( n7834 & n18133 ) | ( ~n15032 & n18133 ) ;
  assign n18137 = n18135 | n18136 ;
  assign n18138 = n7838 & ~n18085 ;
  assign n18139 = n18137 | n18138 ;
  assign n18140 = n18139 ^ x11 ^ 1'b0 ;
  assign n18141 = n18140 ^ n18041 ^ n17872 ;
  assign n18142 = ( ~n17872 & n18041 ) | ( ~n17872 & n18140 ) | ( n18041 & n18140 ) ;
  assign n18143 = n7829 & ~n15032 ;
  assign n18144 = ( n7833 & n15001 ) | ( n7833 & n18143 ) | ( n15001 & n18143 ) ;
  assign n18145 = ( n15032 & n15095 ) | ( n15032 & ~n18095 ) | ( n15095 & ~n18095 ) ;
  assign n18146 = n18143 | n18144 ;
  assign n18147 = ( n7834 & ~n15095 ) | ( n7834 & n18143 ) | ( ~n15095 & n18143 ) ;
  assign n18148 = n18146 | n18147 ;
  assign n18149 = n7838 & n18108 ;
  assign n18150 = n18148 | n18149 ;
  assign n18151 = n18150 ^ x11 ^ 1'b0 ;
  assign n18152 = ( ~n17962 & n18142 ) | ( ~n17962 & n18151 ) | ( n18142 & n18151 ) ;
  assign n18153 = n18151 ^ n18142 ^ n17962 ;
  assign n18154 = n8029 & ~n15095 ;
  assign n18155 = ( n8037 & ~n15032 ) | ( n8037 & n18154 ) | ( ~n15032 & n18154 ) ;
  assign n18156 = n18154 | n18155 ;
  assign n18157 = ( n8033 & ~n15216 ) | ( n8033 & n18154 ) | ( ~n15216 & n18154 ) ;
  assign n18158 = n18145 ^ n15216 ^ n15095 ;
  assign n18159 = n18156 | n18157 ;
  assign n18160 = n8034 & ~n18158 ;
  assign n18161 = n18159 | n18160 ;
  assign n18162 = n18161 ^ x5 ^ 1'b0 ;
  assign n18163 = ( ~n18040 & n18122 ) | ( ~n18040 & n18162 ) | ( n18122 & n18162 ) ;
  assign n18164 = n18162 ^ n18122 ^ n18040 ;
  assign n18165 = n7932 & n15001 ;
  assign n18166 = ( n7943 & ~n14970 ) | ( n7943 & n18165 ) | ( ~n14970 & n18165 ) ;
  assign n18167 = n18165 | n18166 ;
  assign n18168 = ( n7929 & ~n15032 ) | ( n7929 & n18165 ) | ( ~n15032 & n18165 ) ;
  assign n18169 = n18167 | n18168 ;
  assign n18170 = n7930 & ~n18085 ;
  assign n18171 = n18169 & ~n18170 ;
  assign n18172 = n18171 ^ n18170 ^ x8 ;
  assign n18173 = ( ~n17862 & n18036 ) | ( ~n17862 & n18172 ) | ( n18036 & n18172 ) ;
  assign n18174 = n18172 ^ n18036 ^ n17862 ;
  assign n18175 = n8086 & ~n15032 ;
  assign n18176 = ( n8088 & ~n15095 ) | ( n8088 & n18175 ) | ( ~n15095 & n18175 ) ;
  assign n18177 = n18175 | n18176 ;
  assign n18178 = ( n8090 & ~n15216 ) | ( n8090 & n18175 ) | ( ~n15216 & n18175 ) ;
  assign n18179 = n18177 | n18178 ;
  assign n18180 = n18158 & ~n18179 ;
  assign n18181 = ( n8089 & n18179 ) | ( n8089 & ~n18180 ) | ( n18179 & ~n18180 ) ;
  assign n18182 = n18181 ^ x2 ^ 1'b0 ;
  assign n18183 = ( n17995 & n18112 ) | ( n17995 & n18182 ) | ( n18112 & n18182 ) ;
  assign n18184 = n7829 & ~n15095 ;
  assign n18185 = ( n7833 & ~n15032 ) | ( n7833 & n18184 ) | ( ~n15032 & n18184 ) ;
  assign n18186 = n18184 | n18185 ;
  assign n18187 = n7838 & ~n18158 ;
  assign n18188 = ( n7834 & ~n15216 ) | ( n7834 & n18184 ) | ( ~n15216 & n18184 ) ;
  assign n18189 = n18186 | n18188 ;
  assign n18190 = n18187 | n18189 ;
  assign n18191 = n18190 ^ x11 ^ 1'b0 ;
  assign n18192 = n18191 ^ n18152 ^ n18039 ;
  assign n18193 = ( n18039 & n18152 ) | ( n18039 & n18191 ) | ( n18152 & n18191 ) ;
  assign n18194 = ( n15095 & n15216 ) | ( n15095 & n18145 ) | ( n15216 & n18145 ) ;
  assign n18195 = n8086 & ~n15095 ;
  assign n18196 = ( n8088 & ~n15216 ) | ( n8088 & n18195 ) | ( ~n15216 & n18195 ) ;
  assign n18197 = n18195 | n18196 ;
  assign n18198 = ( n8090 & n15218 ) | ( n8090 & n18195 ) | ( n15218 & n18195 ) ;
  assign n18199 = n18197 | n18198 ;
  assign n18200 = n18194 ^ n15218 ^ n15216 ;
  assign n18201 = ~n8089 & n18200 ;
  assign n18202 = ( n18199 & n18200 ) | ( n18199 & ~n18201 ) | ( n18200 & ~n18201 ) ;
  assign n18203 = n18202 ^ x2 ^ 1'b0 ;
  assign n18204 = n7932 & ~n15095 ;
  assign n18205 = ( n18102 & n18183 ) | ( n18102 & n18203 ) | ( n18183 & n18203 ) ;
  assign n18206 = ( n7943 & ~n15032 ) | ( n7943 & n18204 ) | ( ~n15032 & n18204 ) ;
  assign n18207 = n18204 | n18206 ;
  assign n18208 = ( n7929 & ~n15216 ) | ( n7929 & n18204 ) | ( ~n15216 & n18204 ) ;
  assign n18209 = n7932 & ~n15032 ;
  assign n18210 = n18207 | n18208 ;
  assign n18211 = ( n7943 & n15001 ) | ( n7943 & n18209 ) | ( n15001 & n18209 ) ;
  assign n18212 = n18209 | n18211 ;
  assign n18213 = ( n7929 & ~n15095 ) | ( n7929 & n18209 ) | ( ~n15095 & n18209 ) ;
  assign n18214 = n18212 | n18213 ;
  assign n18215 = ( n7930 & n18108 ) | ( n7930 & n18214 ) | ( n18108 & n18214 ) ;
  assign n18216 = n18214 | n18215 ;
  assign n18217 = n18216 ^ x8 ^ 1'b0 ;
  assign n18218 = n18217 ^ n18173 ^ n17921 ;
  assign n18219 = ( n17921 & n18173 ) | ( n17921 & n18217 ) | ( n18173 & n18217 ) ;
  assign n18220 = n7932 & ~n15216 ;
  assign n18221 = ( n7943 & ~n15095 ) | ( n7943 & n18220 ) | ( ~n15095 & n18220 ) ;
  assign n18222 = n18220 | n18221 ;
  assign n18223 = ( n7929 & n15218 ) | ( n7929 & n18220 ) | ( n15218 & n18220 ) ;
  assign n18224 = ( n15216 & ~n15218 ) | ( n15216 & n18194 ) | ( ~n15218 & n18194 ) ;
  assign n18225 = n18222 | n18223 ;
  assign n18226 = ( n7930 & n18200 ) | ( n7930 & n18225 ) | ( n18200 & n18225 ) ;
  assign n18227 = n18225 | n18226 ;
  assign n18228 = n7930 & ~n18158 ;
  assign n18229 = n18210 & ~n18228 ;
  assign n18230 = n18229 ^ n18228 ^ x8 ;
  assign n18231 = n18230 ^ n18219 ^ n18042 ;
  assign n18232 = n18227 ^ x8 ^ 1'b0 ;
  assign n18233 = ( ~n18042 & n18219 ) | ( ~n18042 & n18230 ) | ( n18219 & n18230 ) ;
  assign n18234 = n8086 & ~n15216 ;
  assign n18235 = ( ~n18141 & n18232 ) | ( ~n18141 & n18233 ) | ( n18232 & n18233 ) ;
  assign n18236 = n18233 ^ n18232 ^ n18141 ;
  assign n18237 = n7829 & ~n15216 ;
  assign n18238 = ( n7833 & ~n15095 ) | ( n7833 & n18237 ) | ( ~n15095 & n18237 ) ;
  assign n18239 = n18237 | n18238 ;
  assign n18240 = ( n7834 & n15218 ) | ( n7834 & n18237 ) | ( n15218 & n18237 ) ;
  assign n18241 = n18239 | n18240 ;
  assign n18242 = n7838 & n18200 ;
  assign n18243 = n18241 | n18242 ;
  assign n18244 = n18243 ^ x11 ^ 1'b0 ;
  assign n18245 = ( n8088 & n15218 ) | ( n8088 & n18234 ) | ( n15218 & n18234 ) ;
  assign n18246 = n18234 | n18245 ;
  assign n18247 = ( n8090 & n15219 ) | ( n8090 & n18234 ) | ( n15219 & n18234 ) ;
  assign n18248 = n18246 | n18247 ;
  assign n18249 = n18244 ^ n18193 ^ n18132 ;
  assign n18250 = ( ~n18132 & n18193 ) | ( ~n18132 & n18244 ) | ( n18193 & n18244 ) ;
  assign n18251 = ( n15218 & n15219 ) | ( n15218 & ~n18224 ) | ( n15219 & ~n18224 ) ;
  assign n18252 = n18224 ^ n15219 ^ n15218 ;
  assign n18253 = ~n18248 & n18252 ;
  assign n18254 = ( n8089 & n18248 ) | ( n8089 & ~n18253 ) | ( n18248 & ~n18253 ) ;
  assign n18255 = n18254 ^ x2 ^ 1'b0 ;
  assign n18256 = ( n18121 & n18205 ) | ( n18121 & n18255 ) | ( n18205 & n18255 ) ;
  assign n18257 = n8029 & ~n15216 ;
  assign n18258 = ( n8033 & n15218 ) | ( n8033 & n18257 ) | ( n15218 & n18257 ) ;
  assign n18259 = ( n8037 & ~n15095 ) | ( n8037 & n18257 ) | ( ~n15095 & n18257 ) ;
  assign n18260 = n18257 | n18259 ;
  assign n18261 = n18258 | n18260 ;
  assign n18262 = n8034 & n18200 ;
  assign n18263 = n18261 | n18262 ;
  assign n18264 = n18263 ^ x5 ^ 1'b0 ;
  assign n18265 = ( n18163 & ~n18174 ) | ( n18163 & n18264 ) | ( ~n18174 & n18264 ) ;
  assign n18266 = n8086 & n15218 ;
  assign n18267 = n18264 ^ n18174 ^ n18163 ;
  assign n18268 = ( n8088 & n15219 ) | ( n8088 & n18266 ) | ( n15219 & n18266 ) ;
  assign n18269 = ( n8090 & n15239 ) | ( n8090 & n18266 ) | ( n15239 & n18266 ) ;
  assign n18270 = n18266 | n18268 ;
  assign n18271 = n18269 | n18270 ;
  assign n18272 = n18251 ^ n15239 ^ n15219 ;
  assign n18273 = ~n8089 & n18272 ;
  assign n18274 = ( n18271 & n18272 ) | ( n18271 & ~n18273 ) | ( n18272 & ~n18273 ) ;
  assign n18275 = n8086 & n15219 ;
  assign n18276 = n18274 ^ x2 ^ 1'b0 ;
  assign n18277 = ( ~n18164 & n18256 ) | ( ~n18164 & n18276 ) | ( n18256 & n18276 ) ;
  assign n18278 = ( n8088 & n15239 ) | ( n8088 & n18275 ) | ( n15239 & n18275 ) ;
  assign n18279 = n18275 | n18278 ;
  assign n18280 = ( n8090 & ~n15248 ) | ( n8090 & n18275 ) | ( ~n15248 & n18275 ) ;
  assign n18281 = n18279 | n18280 ;
  assign n18282 = n7932 & n15218 ;
  assign n18283 = ( n15219 & n15239 ) | ( n15219 & n18251 ) | ( n15239 & n18251 ) ;
  assign n18284 = ( n7943 & ~n15216 ) | ( n7943 & n18282 ) | ( ~n15216 & n18282 ) ;
  assign n18285 = n18282 | n18284 ;
  assign n18286 = ( n7929 & n15219 ) | ( n7929 & n18282 ) | ( n15219 & n18282 ) ;
  assign n18287 = n18285 | n18286 ;
  assign n18288 = n7930 & ~n18252 ;
  assign n18289 = n18287 & ~n18288 ;
  assign n18290 = n18289 ^ n18288 ^ x8 ;
  assign n18291 = ( ~n18153 & n18235 ) | ( ~n18153 & n18290 ) | ( n18235 & n18290 ) ;
  assign n18292 = n18290 ^ n18235 ^ n18153 ;
  assign n18293 = n7932 & n15219 ;
  assign n18294 = ( n7943 & n15218 ) | ( n7943 & n18293 ) | ( n15218 & n18293 ) ;
  assign n18295 = n18293 | n18294 ;
  assign n18296 = ( n7929 & n15239 ) | ( n7929 & n18293 ) | ( n15239 & n18293 ) ;
  assign n18297 = n18295 | n18296 ;
  assign n18298 = ( n7930 & n18272 ) | ( n7930 & n18297 ) | ( n18272 & n18297 ) ;
  assign n18299 = n18297 | n18298 ;
  assign n18300 = n18299 ^ x8 ^ 1'b0 ;
  assign n18301 = n18300 ^ n18291 ^ n18192 ;
  assign n18302 = ( n18192 & n18291 ) | ( n18192 & n18300 ) | ( n18291 & n18300 ) ;
  assign n18303 = n18283 ^ n15248 ^ n15239 ;
  assign n18304 = ~n18281 & n18303 ;
  assign n18305 = ( n8089 & n18281 ) | ( n8089 & ~n18304 ) | ( n18281 & ~n18304 ) ;
  assign n18306 = n18305 ^ x2 ^ 1'b0 ;
  assign n18307 = ( ~n18267 & n18277 ) | ( ~n18267 & n18306 ) | ( n18277 & n18306 ) ;
  assign n18308 = n7932 & n15239 ;
  assign n18309 = ( n7943 & n15219 ) | ( n7943 & n18308 ) | ( n15219 & n18308 ) ;
  assign n18310 = n7930 & ~n18303 ;
  assign n18311 = n18308 | n18309 ;
  assign n18312 = ( n7929 & ~n15248 ) | ( n7929 & n18308 ) | ( ~n15248 & n18308 ) ;
  assign n18313 = n18311 | n18312 ;
  assign n18314 = ~n18310 & n18313 ;
  assign n18315 = n18314 ^ n18310 ^ x8 ;
  assign n18316 = n18315 ^ n18302 ^ n18249 ;
  assign n18317 = ( ~n18249 & n18302 ) | ( ~n18249 & n18315 ) | ( n18302 & n18315 ) ;
  assign n18318 = n7669 & ~n15032 ;
  assign n18319 = ( n7667 & ~n15095 ) | ( n7667 & n18318 ) | ( ~n15095 & n18318 ) ;
  assign n18320 = ( n7674 & n15001 ) | ( n7674 & n18318 ) | ( n15001 & n18318 ) ;
  assign n18321 = n18318 | n18320 ;
  assign n18322 = n18319 | n18321 ;
  assign n18323 = ( n7666 & n18108 ) | ( n7666 & n18322 ) | ( n18108 & n18322 ) ;
  assign n18324 = n18322 | n18323 ;
  assign n18325 = n18324 ^ x14 ^ 1'b0 ;
  assign n18326 = ( ~n17971 & n18131 ) | ( ~n17971 & n18325 ) | ( n18131 & n18325 ) ;
  assign n18327 = n18325 ^ n18131 ^ n17971 ;
  assign n18328 = n7838 & ~n18252 ;
  assign n18329 = n7829 & n15218 ;
  assign n18330 = ( n7833 & ~n15216 ) | ( n7833 & n18329 ) | ( ~n15216 & n18329 ) ;
  assign n18331 = n18329 | n18330 ;
  assign n18332 = ( n7834 & n15219 ) | ( n7834 & n18329 ) | ( n15219 & n18329 ) ;
  assign n18333 = n18331 | n18332 ;
  assign n18334 = n18328 | n18333 ;
  assign n18335 = n18334 ^ x11 ^ 1'b0 ;
  assign n18336 = n18335 ^ n18327 ^ n18250 ;
  assign n18337 = ( n18250 & ~n18327 ) | ( n18250 & n18335 ) | ( ~n18327 & n18335 ) ;
  assign n18338 = n8029 & n15218 ;
  assign n18339 = ( n8037 & ~n15216 ) | ( n8037 & n18338 ) | ( ~n15216 & n18338 ) ;
  assign n18340 = n18338 | n18339 ;
  assign n18341 = ( n8033 & n15219 ) | ( n8033 & n18338 ) | ( n15219 & n18338 ) ;
  assign n18342 = n18340 | n18341 ;
  assign n18343 = n8034 & ~n18252 ;
  assign n18344 = n18342 | n18343 ;
  assign n18345 = n18344 ^ x5 ^ 1'b0 ;
  assign n18346 = n18345 ^ n18265 ^ n18218 ;
  assign n18347 = n8086 & n15239 ;
  assign n18348 = ( n18218 & n18265 ) | ( n18218 & n18345 ) | ( n18265 & n18345 ) ;
  assign n18349 = ( n8088 & ~n15248 ) | ( n8088 & n18347 ) | ( ~n15248 & n18347 ) ;
  assign n18350 = ( n8090 & n15271 ) | ( n8090 & n18347 ) | ( n15271 & n18347 ) ;
  assign n18351 = n18347 | n18349 ;
  assign n18352 = n18350 | n18351 ;
  assign n18353 = ( n15239 & ~n15248 ) | ( n15239 & n18283 ) | ( ~n15248 & n18283 ) ;
  assign n18354 = n18353 ^ n15271 ^ n15248 ;
  assign n18355 = ~n18352 & n18354 ;
  assign n18356 = ( n8089 & n18352 ) | ( n8089 & ~n18355 ) | ( n18352 & ~n18355 ) ;
  assign n18357 = n8029 & n15239 ;
  assign n18358 = n18356 ^ x2 ^ 1'b0 ;
  assign n18359 = ( n18307 & n18346 ) | ( n18307 & n18358 ) | ( n18346 & n18358 ) ;
  assign n18360 = ( n8033 & ~n15248 ) | ( n8033 & n18357 ) | ( ~n15248 & n18357 ) ;
  assign n18361 = ( n8037 & n15219 ) | ( n8037 & n18357 ) | ( n15219 & n18357 ) ;
  assign n18362 = n18357 | n18361 ;
  assign n18363 = n18360 | n18362 ;
  assign n18364 = n7669 & ~n15095 ;
  assign n18365 = ( n7674 & ~n15032 ) | ( n7674 & n18364 ) | ( ~n15032 & n18364 ) ;
  assign n18366 = n18364 | n18365 ;
  assign n18367 = ( n7667 & ~n15216 ) | ( n7667 & n18364 ) | ( ~n15216 & n18364 ) ;
  assign n18368 = n18366 | n18367 ;
  assign n18369 = n7666 & ~n18158 ;
  assign n18370 = n18368 & ~n18369 ;
  assign n18371 = n18370 ^ n18369 ^ x14 ;
  assign n18372 = n8034 & ~n18303 ;
  assign n18373 = n18363 | n18372 ;
  assign n18374 = n18373 ^ x5 ^ 1'b0 ;
  assign n18375 = n18371 ^ n18326 ^ n18053 ;
  assign n18376 = ( ~n18053 & n18326 ) | ( ~n18053 & n18371 ) | ( n18326 & n18371 ) ;
  assign n18377 = n8029 & n15219 ;
  assign n18378 = ( n8037 & n15218 ) | ( n8037 & n18377 ) | ( n15218 & n18377 ) ;
  assign n18379 = n18377 | n18378 ;
  assign n18380 = ( n8033 & n15239 ) | ( n8033 & n18377 ) | ( n15239 & n18377 ) ;
  assign n18381 = n18379 | n18380 ;
  assign n18382 = n8034 & n18272 ;
  assign n18383 = n18381 | n18382 ;
  assign n18384 = n18383 ^ x5 ^ 1'b0 ;
  assign n18385 = n18384 ^ n18348 ^ n18231 ;
  assign n18386 = ( ~n18231 & n18348 ) | ( ~n18231 & n18384 ) | ( n18348 & n18384 ) ;
  assign n18387 = n18386 ^ n18374 ^ n18236 ;
  assign n18388 = ( ~n18236 & n18374 ) | ( ~n18236 & n18386 ) | ( n18374 & n18386 ) ;
  assign n18389 = n8029 & ~n15248 ;
  assign n18390 = ( n8037 & n15239 ) | ( n8037 & n18389 ) | ( n15239 & n18389 ) ;
  assign n18391 = n18389 | n18390 ;
  assign n18392 = ( n8033 & n15271 ) | ( n8033 & n18389 ) | ( n15271 & n18389 ) ;
  assign n18393 = n18391 | n18392 ;
  assign n18394 = n8034 & ~n18354 ;
  assign n18395 = n18393 | n18394 ;
  assign n18396 = n18395 ^ x5 ^ 1'b0 ;
  assign n18397 = n18396 ^ n18388 ^ n18292 ;
  assign n18398 = ( ~n18292 & n18388 ) | ( ~n18292 & n18396 ) | ( n18388 & n18396 ) ;
  assign n18399 = n7932 & ~n15248 ;
  assign n18400 = ( n7943 & n15239 ) | ( n7943 & n18399 ) | ( n15239 & n18399 ) ;
  assign n18401 = n18399 | n18400 ;
  assign n18402 = ( n7929 & n15271 ) | ( n7929 & n18399 ) | ( n15271 & n18399 ) ;
  assign n18403 = n18401 | n18402 ;
  assign n18404 = n7930 & ~n18354 ;
  assign n18405 = n18403 & ~n18404 ;
  assign n18406 = n18405 ^ n18404 ^ x8 ;
  assign n18407 = ( n18317 & ~n18336 ) | ( n18317 & n18406 ) | ( ~n18336 & n18406 ) ;
  assign n18408 = n18406 ^ n18336 ^ n18317 ;
  assign n18409 = n7829 & n15219 ;
  assign n18410 = ( n7833 & n15218 ) | ( n7833 & n18409 ) | ( n15218 & n18409 ) ;
  assign n18411 = n18409 | n18410 ;
  assign n18412 = ( n7834 & n15239 ) | ( n7834 & n18409 ) | ( n15239 & n18409 ) ;
  assign n18413 = n18411 | n18412 ;
  assign n18414 = n7838 & n18272 ;
  assign n18415 = n18413 | n18414 ;
  assign n18416 = n18415 ^ x11 ^ 1'b0 ;
  assign n18417 = n18416 ^ n18375 ^ n18337 ;
  assign n18418 = ( n18337 & ~n18375 ) | ( n18337 & n18416 ) | ( ~n18375 & n18416 ) ;
  assign n18419 = n7485 & n15001 ;
  assign n18420 = ( n7486 & ~n15032 ) | ( n7486 & n18419 ) | ( ~n15032 & n18419 ) ;
  assign n18421 = n18419 | n18420 ;
  assign n18422 = ( n7493 & ~n14970 ) | ( n7493 & n18419 ) | ( ~n14970 & n18419 ) ;
  assign n18423 = n18421 | n18422 ;
  assign n18424 = n7487 & ~n18085 ;
  assign n18425 = n18423 | n18424 ;
  assign n18426 = n18425 ^ x17 ^ 1'b0 ;
  assign n18427 = n18426 ^ n18052 ^ n17841 ;
  assign n18428 = ( ~n17841 & n18052 ) | ( ~n17841 & n18426 ) | ( n18052 & n18426 ) ;
  assign n18429 = n7669 & ~n15216 ;
  assign n18430 = ( n7674 & ~n15095 ) | ( n7674 & n18429 ) | ( ~n15095 & n18429 ) ;
  assign n18431 = n18429 | n18430 ;
  assign n18432 = ( n7667 & n15218 ) | ( n7667 & n18429 ) | ( n15218 & n18429 ) ;
  assign n18433 = n18431 | n18432 ;
  assign n18434 = ( n7666 & n18200 ) | ( n7666 & n18433 ) | ( n18200 & n18433 ) ;
  assign n18435 = n18433 | n18434 ;
  assign n18436 = n18435 ^ x14 ^ 1'b0 ;
  assign n18437 = n18436 ^ n18427 ^ n18376 ;
  assign n18438 = ( n18376 & ~n18427 ) | ( n18376 & n18436 ) | ( ~n18427 & n18436 ) ;
  assign n18439 = n7829 & n15239 ;
  assign n18440 = ( n7833 & n15219 ) | ( n7833 & n18439 ) | ( n15219 & n18439 ) ;
  assign n18441 = n18439 | n18440 ;
  assign n18442 = ( n7834 & ~n15248 ) | ( n7834 & n18439 ) | ( ~n15248 & n18439 ) ;
  assign n18443 = n18441 | n18442 ;
  assign n18444 = n7838 & ~n18303 ;
  assign n18445 = n18443 | n18444 ;
  assign n18446 = n18445 ^ x11 ^ 1'b0 ;
  assign n18447 = n18446 ^ n18437 ^ n18418 ;
  assign n18448 = ( n18418 & ~n18437 ) | ( n18418 & n18446 ) | ( ~n18437 & n18446 ) ;
  assign n18449 = ( ~n15248 & n15271 ) | ( ~n15248 & n18353 ) | ( n15271 & n18353 ) ;
  assign n18450 = n8086 & ~n15248 ;
  assign n18451 = ( n8090 & ~n15275 ) | ( n8090 & n18450 ) | ( ~n15275 & n18450 ) ;
  assign n18452 = n8029 & n15271 ;
  assign n18453 = ( n8088 & n15271 ) | ( n8088 & n18450 ) | ( n15271 & n18450 ) ;
  assign n18454 = n18450 | n18453 ;
  assign n18455 = n18451 | n18454 ;
  assign n18456 = n18449 ^ n15275 ^ n15271 ;
  assign n18457 = ~n18455 & n18456 ;
  assign n18458 = ( n8089 & n18455 ) | ( n8089 & ~n18457 ) | ( n18455 & ~n18457 ) ;
  assign n18459 = n18458 ^ x2 ^ 1'b0 ;
  assign n18460 = ( n18359 & ~n18385 ) | ( n18359 & n18459 ) | ( ~n18385 & n18459 ) ;
  assign n18461 = n18459 ^ n18385 ^ n18359 ;
  assign n18462 = ( n8037 & ~n15248 ) | ( n8037 & n18452 ) | ( ~n15248 & n18452 ) ;
  assign n18463 = ( n8033 & ~n15275 ) | ( n8033 & n18452 ) | ( ~n15275 & n18452 ) ;
  assign n18464 = n18452 | n18462 ;
  assign n18465 = n18463 | n18464 ;
  assign n18466 = n7930 & ~n18456 ;
  assign n18467 = n8034 & ~n18456 ;
  assign n18468 = n18465 | n18467 ;
  assign n18469 = n18468 ^ x5 ^ 1'b0 ;
  assign n18470 = n18469 ^ n18398 ^ n18301 ;
  assign n18471 = ( n18301 & n18398 ) | ( n18301 & n18469 ) | ( n18398 & n18469 ) ;
  assign n18472 = n7932 & n15271 ;
  assign n18473 = ( n15271 & ~n15275 ) | ( n15271 & n18449 ) | ( ~n15275 & n18449 ) ;
  assign n18474 = ( n7943 & ~n15248 ) | ( n7943 & n18472 ) | ( ~n15248 & n18472 ) ;
  assign n18475 = n18472 | n18474 ;
  assign n18476 = ( n7929 & ~n15275 ) | ( n7929 & n18472 ) | ( ~n15275 & n18472 ) ;
  assign n18477 = n18475 | n18476 ;
  assign n18478 = ( ~n15275 & n15312 ) | ( ~n15275 & n18473 ) | ( n15312 & n18473 ) ;
  assign n18479 = ~n18466 & n18477 ;
  assign n18480 = n18473 ^ n15312 ^ n15275 ;
  assign n18481 = n18479 ^ n18466 ^ x8 ;
  assign n18482 = ( n18407 & ~n18417 ) | ( n18407 & n18481 ) | ( ~n18417 & n18481 ) ;
  assign n18483 = n18481 ^ n18417 ^ n18407 ;
  assign n18484 = n8086 & n15271 ;
  assign n18485 = ( n8088 & ~n15275 ) | ( n8088 & n18484 ) | ( ~n15275 & n18484 ) ;
  assign n18486 = n18484 | n18485 ;
  assign n18487 = ( n8090 & n15312 ) | ( n8090 & n18484 ) | ( n15312 & n18484 ) ;
  assign n18488 = n18486 | n18487 ;
  assign n18489 = n18480 & ~n18488 ;
  assign n18490 = ( n8089 & n18488 ) | ( n8089 & ~n18489 ) | ( n18488 & ~n18489 ) ;
  assign n18491 = n18490 ^ x2 ^ 1'b0 ;
  assign n18492 = ( ~n18387 & n18460 ) | ( ~n18387 & n18491 ) | ( n18460 & n18491 ) ;
  assign n18493 = n18491 ^ n18460 ^ n18387 ;
  assign n18494 = n7932 & ~n15275 ;
  assign n18495 = ( n7943 & n15271 ) | ( n7943 & n18494 ) | ( n15271 & n18494 ) ;
  assign n18496 = n18494 | n18495 ;
  assign n18497 = ( n7929 & n15312 ) | ( n7929 & n18494 ) | ( n15312 & n18494 ) ;
  assign n18498 = n18496 | n18497 ;
  assign n18499 = n7930 & ~n18480 ;
  assign n18500 = n18498 & ~n18499 ;
  assign n18501 = n18500 ^ n18499 ^ x8 ;
  assign n18502 = n18501 ^ n18482 ^ n18447 ;
  assign n18503 = ( ~n18447 & n18482 ) | ( ~n18447 & n18501 ) | ( n18482 & n18501 ) ;
  assign n18504 = n8029 & ~n15275 ;
  assign n18505 = ( n8037 & n15271 ) | ( n8037 & n18504 ) | ( n15271 & n18504 ) ;
  assign n18506 = n18504 | n18505 ;
  assign n18507 = ( n8033 & n15312 ) | ( n8033 & n18504 ) | ( n15312 & n18504 ) ;
  assign n18508 = n18506 | n18507 ;
  assign n18509 = n8034 & ~n18480 ;
  assign n18510 = n18508 | n18509 ;
  assign n18511 = n18510 ^ x5 ^ 1'b0 ;
  assign n18512 = ( ~n18316 & n18471 ) | ( ~n18316 & n18511 ) | ( n18471 & n18511 ) ;
  assign n18513 = n18511 ^ n18471 ^ n18316 ;
  assign n18514 = n8029 & n15312 ;
  assign n18515 = ( n8037 & ~n15275 ) | ( n8037 & n18514 ) | ( ~n15275 & n18514 ) ;
  assign n18516 = n18514 | n18515 ;
  assign n18517 = ( n8033 & n15308 ) | ( n8033 & n18514 ) | ( n15308 & n18514 ) ;
  assign n18518 = n18516 | n18517 ;
  assign n18519 = n8086 & ~n15275 ;
  assign n18520 = ( n15308 & n15312 ) | ( n15308 & n18478 ) | ( n15312 & n18478 ) ;
  assign n18521 = ( n8088 & n15312 ) | ( n8088 & n18519 ) | ( n15312 & n18519 ) ;
  assign n18522 = n18519 | n18521 ;
  assign n18523 = ( n8090 & n15308 ) | ( n8090 & n18519 ) | ( n15308 & n18519 ) ;
  assign n18524 = n18522 | n18523 ;
  assign n18525 = n18478 ^ n15312 ^ n15308 ;
  assign n18526 = ~n8089 & n18525 ;
  assign n18527 = ( n18524 & n18525 ) | ( n18524 & ~n18526 ) | ( n18525 & ~n18526 ) ;
  assign n18528 = n18527 ^ x2 ^ 1'b0 ;
  assign n18529 = n18528 ^ n18492 ^ n18397 ;
  assign n18530 = ( ~n18397 & n18492 ) | ( ~n18397 & n18528 ) | ( n18492 & n18528 ) ;
  assign n18531 = n18520 ^ n15319 ^ n15308 ;
  assign n18532 = n8086 & n15312 ;
  assign n18533 = ( n8088 & n15308 ) | ( n8088 & n18532 ) | ( n15308 & n18532 ) ;
  assign n18534 = n18532 | n18533 ;
  assign n18535 = ( n8090 & n15319 ) | ( n8090 & n18532 ) | ( n15319 & n18532 ) ;
  assign n18536 = n18534 | n18535 ;
  assign n18537 = ~n8089 & n18531 ;
  assign n18538 = ( n18531 & n18536 ) | ( n18531 & ~n18537 ) | ( n18536 & ~n18537 ) ;
  assign n18539 = n18538 ^ x2 ^ 1'b0 ;
  assign n18540 = ( n18470 & n18530 ) | ( n18470 & n18539 ) | ( n18530 & n18539 ) ;
  assign n18541 = n18539 ^ n18530 ^ n18470 ;
  assign n18542 = n8086 & n15308 ;
  assign n18543 = ( n15308 & n15319 ) | ( n15308 & n18520 ) | ( n15319 & n18520 ) ;
  assign n18544 = ( n8090 & ~n15320 ) | ( n8090 & n18542 ) | ( ~n15320 & n18542 ) ;
  assign n18545 = n8034 & n18525 ;
  assign n18546 = n18518 | n18545 ;
  assign n18547 = ( n8088 & n15319 ) | ( n8088 & n18542 ) | ( n15319 & n18542 ) ;
  assign n18548 = n18542 | n18547 ;
  assign n18549 = ( n15319 & ~n15320 ) | ( n15319 & n18543 ) | ( ~n15320 & n18543 ) ;
  assign n18550 = n18549 ^ n15322 ^ n15320 ;
  assign n18551 = n18544 | n18548 ;
  assign n18552 = n18543 ^ n15320 ^ n15319 ;
  assign n18553 = ~n18551 & n18552 ;
  assign n18554 = ( n8089 & n18551 ) | ( n8089 & ~n18553 ) | ( n18551 & ~n18553 ) ;
  assign n18555 = n8089 & ~n18550 ;
  assign n18556 = ( n8086 & n15319 ) | ( n8086 & n18555 ) | ( n15319 & n18555 ) ;
  assign n18557 = n18555 | n18556 ;
  assign n18558 = ( n8088 & ~n15320 ) | ( n8088 & n18555 ) | ( ~n15320 & n18555 ) ;
  assign n18559 = n18554 ^ x2 ^ 1'b0 ;
  assign n18560 = n18557 | n18558 ;
  assign n18561 = n18559 ^ n18540 ^ n18513 ;
  assign n18562 = ( ~n18513 & n18540 ) | ( ~n18513 & n18559 ) | ( n18540 & n18559 ) ;
  assign n18563 = n18546 ^ x5 ^ 1'b0 ;
  assign n18564 = ( ~n18408 & n18512 ) | ( ~n18408 & n18563 ) | ( n18512 & n18563 ) ;
  assign n18565 = n18560 ^ x2 ^ 1'b0 ;
  assign n18566 = n18563 ^ n18512 ^ n18408 ;
  assign n18567 = n8034 & ~n18550 ;
  assign n18568 = ( n8029 & ~n15320 ) | ( n8029 & n18567 ) | ( ~n15320 & n18567 ) ;
  assign n18569 = n18567 | n18568 ;
  assign n18570 = ( n8037 & n15319 ) | ( n8037 & n18567 ) | ( n15319 & n18567 ) ;
  assign n18571 = n18569 | n18570 ;
  assign n18572 = ( n18562 & n18565 ) | ( n18562 & ~n18566 ) | ( n18565 & ~n18566 ) ;
  assign n18573 = n18566 ^ n18565 ^ n18562 ;
  assign n18574 = n8029 & n15308 ;
  assign n18575 = ( n8037 & n15312 ) | ( n8037 & n18574 ) | ( n15312 & n18574 ) ;
  assign n18576 = n18574 | n18575 ;
  assign n18577 = ( n8033 & n15319 ) | ( n8033 & n18574 ) | ( n15319 & n18574 ) ;
  assign n18578 = n8029 & n15319 ;
  assign n18579 = n18576 | n18577 ;
  assign n18580 = ( n8037 & n15308 ) | ( n8037 & n18578 ) | ( n15308 & n18578 ) ;
  assign n18581 = n18578 | n18580 ;
  assign n18582 = ( n8033 & ~n15320 ) | ( n8033 & n18578 ) | ( ~n15320 & n18578 ) ;
  assign n18583 = n8034 & n18531 ;
  assign n18584 = n8034 & ~n18552 ;
  assign n18585 = n8086 & ~n15320 ;
  assign n18586 = n18579 | n18583 ;
  assign n18587 = n18586 ^ x5 ^ 1'b0 ;
  assign n18588 = n18587 ^ n18564 ^ n18483 ;
  assign n18589 = ( ~n18483 & n18564 ) | ( ~n18483 & n18587 ) | ( n18564 & n18587 ) ;
  assign n18590 = n18581 | n18582 ;
  assign n18591 = n18585 ^ x2 ^ 1'b0 ;
  assign n18592 = n18591 ^ n18588 ^ n18572 ;
  assign n18593 = ( n18572 & ~n18588 ) | ( n18572 & n18591 ) | ( ~n18588 & n18591 ) ;
  assign n18594 = n18584 | n18590 ;
  assign n18595 = n18594 ^ x5 ^ 1'b0 ;
  assign n18596 = n18595 ^ n18502 ^ x2 ;
  assign n18597 = n18596 ^ n18593 ^ n18589 ;
  assign n18598 = ( x2 & ~n18502 ) | ( x2 & n18595 ) | ( ~n18502 & n18595 ) ;
  assign n18599 = ( n18589 & n18593 ) | ( n18589 & ~n18596 ) | ( n18593 & ~n18596 ) ;
  assign n18600 = n7485 & ~n15032 ;
  assign n18601 = ( n7486 & ~n15095 ) | ( n7486 & n18600 ) | ( ~n15095 & n18600 ) ;
  assign n18602 = n18600 | n18601 ;
  assign n18603 = ( n7493 & n15001 ) | ( n7493 & n18600 ) | ( n15001 & n18600 ) ;
  assign n18604 = n18602 | n18603 ;
  assign n18605 = n7487 & n18108 ;
  assign n18606 = n18604 | n18605 ;
  assign n18607 = n18606 ^ x17 ^ 1'b0 ;
  assign n18608 = n18607 ^ n17951 ^ n17842 ;
  assign n18609 = ( n17842 & ~n17951 ) | ( n17842 & n18607 ) | ( ~n17951 & n18607 ) ;
  assign n18610 = n7669 & n15218 ;
  assign n18611 = ( n7674 & ~n15216 ) | ( n7674 & n18610 ) | ( ~n15216 & n18610 ) ;
  assign n18612 = n18610 | n18611 ;
  assign n18613 = ( n7667 & n15219 ) | ( n7667 & n18610 ) | ( n15219 & n18610 ) ;
  assign n18614 = n18612 | n18613 ;
  assign n18615 = n7666 & ~n18252 ;
  assign n18616 = n18614 | n18615 ;
  assign n18617 = n18616 ^ x14 ^ 1'b0 ;
  assign n18618 = ( n18428 & ~n18608 ) | ( n18428 & n18617 ) | ( ~n18608 & n18617 ) ;
  assign n18619 = n18617 ^ n18608 ^ n18428 ;
  assign n18620 = n7829 & ~n15248 ;
  assign n18621 = ( n7833 & n15239 ) | ( n7833 & n18620 ) | ( n15239 & n18620 ) ;
  assign n18622 = n18620 | n18621 ;
  assign n18623 = ( n7834 & n15271 ) | ( n7834 & n18620 ) | ( n15271 & n18620 ) ;
  assign n18624 = n18622 | n18623 ;
  assign n18625 = n7838 & ~n18354 ;
  assign n18626 = n18624 | n18625 ;
  assign n18627 = n18626 ^ x11 ^ 1'b0 ;
  assign n18628 = ( n18438 & ~n18619 ) | ( n18438 & n18627 ) | ( ~n18619 & n18627 ) ;
  assign n18629 = n18627 ^ n18619 ^ n18438 ;
  assign n18630 = n7485 & ~n15095 ;
  assign n18631 = ( n7486 & ~n15216 ) | ( n7486 & n18630 ) | ( ~n15216 & n18630 ) ;
  assign n18632 = n18630 | n18631 ;
  assign n18633 = ( n7493 & ~n15032 ) | ( n7493 & n18630 ) | ( ~n15032 & n18630 ) ;
  assign n18634 = n18571 ^ x5 ^ 1'b0 ;
  assign n18635 = n18632 | n18633 ;
  assign n18636 = n7487 & ~n18158 ;
  assign n18637 = n18635 | n18636 ;
  assign n18638 = n18637 ^ x17 ^ 1'b0 ;
  assign n18639 = ( n17952 & n18073 ) | ( n17952 & n18638 ) | ( n18073 & n18638 ) ;
  assign n18640 = n18638 ^ n18073 ^ n17952 ;
  assign n18641 = n7932 & n15312 ;
  assign n18642 = ( n7943 & ~n15275 ) | ( n7943 & n18641 ) | ( ~n15275 & n18641 ) ;
  assign n18643 = n18641 | n18642 ;
  assign n18644 = ( n7929 & n15308 ) | ( n7929 & n18641 ) | ( n15308 & n18641 ) ;
  assign n18645 = n18643 | n18644 ;
  assign n18646 = n7930 & n18525 ;
  assign n18647 = n18645 | n18646 ;
  assign n18648 = n18647 ^ x8 ^ 1'b0 ;
  assign n18649 = n18648 ^ n18629 ^ n18448 ;
  assign n18650 = ( n18448 & ~n18629 ) | ( n18448 & n18648 ) | ( ~n18629 & n18648 ) ;
  assign n18651 = n18649 ^ n18634 ^ n18503 ;
  assign n18652 = ( n18503 & n18634 ) | ( n18503 & ~n18649 ) | ( n18634 & ~n18649 ) ;
  assign n18653 = n18651 ^ n18599 ^ n18598 ;
  assign n18654 = ( n18598 & n18599 ) | ( n18598 & ~n18651 ) | ( n18599 & ~n18651 ) ;
  assign n18655 = n7669 & n15219 ;
  assign n18656 = ( n7674 & n15218 ) | ( n7674 & n18655 ) | ( n15218 & n18655 ) ;
  assign n18657 = n18655 | n18656 ;
  assign n18658 = ( n7667 & n15239 ) | ( n7667 & n18655 ) | ( n15239 & n18655 ) ;
  assign n18659 = n18657 | n18658 ;
  assign n18660 = n7666 & n18272 ;
  assign n18661 = n18659 | n18660 ;
  assign n18662 = n18661 ^ x14 ^ 1'b0 ;
  assign n18663 = n18662 ^ n18640 ^ n18609 ;
  assign n18664 = ( n18609 & n18640 ) | ( n18609 & n18662 ) | ( n18640 & n18662 ) ;
  assign n18665 = n7829 & n15271 ;
  assign n18666 = ( n7833 & ~n15248 ) | ( n7833 & n18665 ) | ( ~n15248 & n18665 ) ;
  assign n18667 = n18665 | n18666 ;
  assign n18668 = ( n7834 & ~n15275 ) | ( n7834 & n18665 ) | ( ~n15275 & n18665 ) ;
  assign n18669 = n18667 | n18668 ;
  assign n18670 = n7838 & ~n18456 ;
  assign n18671 = n18669 | n18670 ;
  assign n18672 = n18671 ^ x11 ^ 1'b0 ;
  assign n18673 = n18672 ^ n18663 ^ n18618 ;
  assign n18674 = ( n18618 & n18663 ) | ( n18618 & n18672 ) | ( n18663 & n18672 ) ;
  assign n18675 = n7932 & n15308 ;
  assign n18676 = ( n7943 & n15312 ) | ( n7943 & n18675 ) | ( n15312 & n18675 ) ;
  assign n18677 = n18675 | n18676 ;
  assign n18678 = ( n7929 & n15319 ) | ( n7929 & n18675 ) | ( n15319 & n18675 ) ;
  assign n18679 = n18677 | n18678 ;
  assign n18680 = n7930 & n18531 ;
  assign n18681 = n18679 | n18680 ;
  assign n18682 = n18681 ^ x8 ^ 1'b0 ;
  assign n18683 = ( n18628 & n18673 ) | ( n18628 & n18682 ) | ( n18673 & n18682 ) ;
  assign n18684 = n18682 ^ n18673 ^ n18628 ;
  assign n18685 = n7339 & ~n15095 ;
  assign n18686 = ( n7337 & ~n15216 ) | ( n7337 & n18685 ) | ( ~n15216 & n18685 ) ;
  assign n18687 = n18685 | n18686 ;
  assign n18688 = ( n7338 & ~n15032 ) | ( n7338 & n18685 ) | ( ~n15032 & n18685 ) ;
  assign n18689 = n8037 & ~n15320 ;
  assign n18690 = n18689 ^ x5 ^ 1'b0 ;
  assign n18691 = n18687 | n18688 ;
  assign n18692 = ( n18650 & n18684 ) | ( n18650 & n18690 ) | ( n18684 & n18690 ) ;
  assign n18693 = n18690 ^ n18684 ^ n18650 ;
  assign n18694 = n7932 & ~n15320 ;
  assign n18695 = ( n7943 & n15319 ) | ( n7943 & n18694 ) | ( n15319 & n18694 ) ;
  assign n18696 = n18694 | n18695 ;
  assign n18697 = ( n7930 & ~n18550 ) | ( n7930 & n18694 ) | ( ~n18550 & n18694 ) ;
  assign n18698 = n18696 | n18697 ;
  assign n18699 = n7340 & ~n18158 ;
  assign n18700 = n18691 | n18699 ;
  assign n18701 = n18698 ^ x8 ^ 1'b0 ;
  assign n18702 = ( n18652 & n18654 ) | ( n18652 & n18693 ) | ( n18654 & n18693 ) ;
  assign n18703 = n7930 & ~n18552 ;
  assign n18704 = n18693 ^ n18652 ^ 1'b0 ;
  assign n18705 = n7932 & n15319 ;
  assign n18706 = ( n7929 & ~n15320 ) | ( n7929 & n18705 ) | ( ~n15320 & n18705 ) ;
  assign n18707 = n18700 ^ x20 ^ 1'b0 ;
  assign n18708 = ( n17932 & n18021 ) | ( n17932 & n18707 ) | ( n18021 & n18707 ) ;
  assign n18709 = n18704 ^ n18654 ^ 1'b0 ;
  assign n18710 = ( n7943 & n15308 ) | ( n7943 & n18705 ) | ( n15308 & n18705 ) ;
  assign n18711 = n7943 & ~n15320 ;
  assign n18712 = n18707 ^ n18021 ^ n17932 ;
  assign n18713 = n18705 | n18710 ;
  assign n18714 = n18706 | n18713 ;
  assign n18715 = n18703 | n18714 ;
  assign n18716 = n18715 ^ x8 ^ 1'b0 ;
  assign n18717 = n7339 & n15001 ;
  assign n18718 = ( n7337 & ~n15032 ) | ( n7337 & n18717 ) | ( ~n15032 & n18717 ) ;
  assign n18719 = n18717 | n18718 ;
  assign n18720 = ( n7338 & ~n14970 ) | ( n7338 & n18717 ) | ( ~n14970 & n18717 ) ;
  assign n18721 = n18719 | n18720 ;
  assign n18722 = n7340 & ~n18085 ;
  assign n18723 = n18721 | n18722 ;
  assign n18724 = n18723 ^ x20 ^ 1'b0 ;
  assign n18725 = ( n17663 & n17822 ) | ( n17663 & n18724 ) | ( n17822 & n18724 ) ;
  assign n18726 = n18724 ^ n17822 ^ n17663 ;
  assign n18727 = n7485 & ~n15216 ;
  assign n18728 = ( n7486 & n15218 ) | ( n7486 & n18727 ) | ( n15218 & n18727 ) ;
  assign n18729 = n18727 | n18728 ;
  assign n18730 = ( n7493 & ~n15095 ) | ( n7493 & n18727 ) | ( ~n15095 & n18727 ) ;
  assign n18731 = n18729 | n18730 ;
  assign n18732 = n7487 & n18200 ;
  assign n18733 = n18731 | n18732 ;
  assign n18734 = n18733 ^ x17 ^ 1'b0 ;
  assign n18735 = ( n18072 & n18726 ) | ( n18072 & n18734 ) | ( n18726 & n18734 ) ;
  assign n18736 = n18734 ^ n18726 ^ n18072 ;
  assign n18737 = n7339 & ~n15032 ;
  assign n18738 = ( n7337 & ~n15095 ) | ( n7337 & n18737 ) | ( ~n15095 & n18737 ) ;
  assign n18739 = n18737 | n18738 ;
  assign n18740 = ( n7338 & n15001 ) | ( n7338 & n18737 ) | ( n15001 & n18737 ) ;
  assign n18741 = n18739 | n18740 ;
  assign n18742 = n7340 & n18108 ;
  assign n18743 = n18741 | n18742 ;
  assign n18744 = n18743 ^ x20 ^ 1'b0 ;
  assign n18745 = n18744 ^ n18725 ^ n17931 ;
  assign n18746 = ( n17931 & n18725 ) | ( n17931 & n18744 ) | ( n18725 & n18744 ) ;
  assign n18747 = n7669 & n15239 ;
  assign n18748 = ( n7674 & n15219 ) | ( n7674 & n18747 ) | ( n15219 & n18747 ) ;
  assign n18749 = n18747 | n18748 ;
  assign n18750 = ( n7667 & ~n15248 ) | ( n7667 & n18747 ) | ( ~n15248 & n18747 ) ;
  assign n18751 = n18749 | n18750 ;
  assign n18752 = n7666 & ~n18303 ;
  assign n18753 = n18751 | n18752 ;
  assign n18754 = n18753 ^ x14 ^ 1'b0 ;
  assign n18755 = n18754 ^ n18736 ^ n18639 ;
  assign n18756 = ( n18639 & n18736 ) | ( n18639 & n18754 ) | ( n18736 & n18754 ) ;
  assign n18757 = n7829 & ~n15275 ;
  assign n18758 = ( n7833 & n15271 ) | ( n7833 & n18757 ) | ( n15271 & n18757 ) ;
  assign n18759 = n18757 | n18758 ;
  assign n18760 = ( n7834 & n15312 ) | ( n7834 & n18757 ) | ( n15312 & n18757 ) ;
  assign n18761 = n18759 | n18760 ;
  assign n18762 = n7838 & ~n18480 ;
  assign n18763 = n18761 | n18762 ;
  assign n18764 = n18763 ^ x11 ^ 1'b0 ;
  assign n18765 = ( n18664 & n18755 ) | ( n18664 & n18764 ) | ( n18755 & n18764 ) ;
  assign n18766 = n18764 ^ n18755 ^ n18664 ;
  assign n18767 = n7485 & n15218 ;
  assign n18768 = ( n7486 & n15219 ) | ( n7486 & n18767 ) | ( n15219 & n18767 ) ;
  assign n18769 = n18767 | n18768 ;
  assign n18770 = ( n7493 & ~n15216 ) | ( n7493 & n18767 ) | ( ~n15216 & n18767 ) ;
  assign n18771 = n18769 | n18770 ;
  assign n18772 = n7487 & ~n18252 ;
  assign n18773 = n18771 | n18772 ;
  assign n18774 = n18766 ^ n18716 ^ n18674 ;
  assign n18775 = ( n18674 & n18716 ) | ( n18674 & n18766 ) | ( n18716 & n18766 ) ;
  assign n18776 = n18711 ^ x8 ^ 1'b0 ;
  assign n18777 = ( x5 & n18683 ) | ( x5 & n18774 ) | ( n18683 & n18774 ) ;
  assign n18778 = n7666 & ~n18354 ;
  assign n18779 = n18774 ^ n18683 ^ x5 ;
  assign n18780 = n18773 ^ x17 ^ 1'b0 ;
  assign n18781 = n18779 ^ n18692 ^ 1'b0 ;
  assign n18782 = ( n18692 & n18702 ) | ( n18692 & n18779 ) | ( n18702 & n18779 ) ;
  assign n18783 = n7669 & ~n15248 ;
  assign n18784 = n18781 ^ n18702 ^ 1'b0 ;
  assign n18785 = ( n7674 & n15239 ) | ( n7674 & n18783 ) | ( n15239 & n18783 ) ;
  assign n18786 = n18783 | n18785 ;
  assign n18787 = ( n7667 & n15271 ) | ( n7667 & n18783 ) | ( n15271 & n18783 ) ;
  assign n18788 = n18786 | n18787 ;
  assign n18789 = n18778 | n18788 ;
  assign n18790 = n18789 ^ x14 ^ 1'b0 ;
  assign n18791 = ( n18735 & n18745 ) | ( n18735 & n18780 ) | ( n18745 & n18780 ) ;
  assign n18792 = n18780 ^ n18745 ^ n18735 ;
  assign n18793 = n18792 ^ n18790 ^ n18756 ;
  assign n18794 = ( n18756 & n18790 ) | ( n18756 & n18792 ) | ( n18790 & n18792 ) ;
  assign n18795 = n7485 & n15219 ;
  assign n18796 = ( n7486 & n15239 ) | ( n7486 & n18795 ) | ( n15239 & n18795 ) ;
  assign n18797 = n18795 | n18796 ;
  assign n18798 = ( n7493 & n15218 ) | ( n7493 & n18795 ) | ( n15218 & n18795 ) ;
  assign n18799 = n18797 | n18798 ;
  assign n18800 = n7487 & n18272 ;
  assign n18801 = n18799 | n18800 ;
  assign n18802 = n18801 ^ x17 ^ 1'b0 ;
  assign n18803 = ( n18712 & n18746 ) | ( n18712 & n18802 ) | ( n18746 & n18802 ) ;
  assign n18804 = n18802 ^ n18746 ^ n18712 ;
  assign n18805 = n7669 & n15271 ;
  assign n18806 = ( n7674 & ~n15248 ) | ( n7674 & n18805 ) | ( ~n15248 & n18805 ) ;
  assign n18807 = n18805 | n18806 ;
  assign n18808 = ( n7667 & ~n15275 ) | ( n7667 & n18805 ) | ( ~n15275 & n18805 ) ;
  assign n18809 = n18807 | n18808 ;
  assign n18810 = n7666 & ~n18456 ;
  assign n18811 = n18809 | n18810 ;
  assign n18812 = n18811 ^ x14 ^ 1'b0 ;
  assign n18813 = ( n18791 & n18804 ) | ( n18791 & n18812 ) | ( n18804 & n18812 ) ;
  assign n18814 = n18812 ^ n18804 ^ n18791 ;
  assign n18815 = n7829 & n15312 ;
  assign n18816 = ( n7833 & ~n15275 ) | ( n7833 & n18815 ) | ( ~n15275 & n18815 ) ;
  assign n18817 = n18815 | n18816 ;
  assign n18818 = ( n7834 & n15308 ) | ( n7834 & n18815 ) | ( n15308 & n18815 ) ;
  assign n18819 = n18817 | n18818 ;
  assign n18820 = n7838 & n18525 ;
  assign n18821 = n18819 | n18820 ;
  assign n18822 = n18821 ^ x11 ^ 1'b0 ;
  assign n18823 = ( n18765 & n18793 ) | ( n18765 & n18822 ) | ( n18793 & n18822 ) ;
  assign n18824 = n18822 ^ n18793 ^ n18765 ;
  assign n18825 = n18824 ^ n18775 ^ n18701 ;
  assign n18826 = n18825 ^ n18777 ^ 1'b0 ;
  assign n18827 = ( n18777 & n18782 ) | ( n18777 & n18825 ) | ( n18782 & n18825 ) ;
  assign n18828 = n18826 ^ n18782 ^ 1'b0 ;
  assign n18829 = n7829 & n15319 ;
  assign n18830 = ( n18701 & n18775 ) | ( n18701 & n18824 ) | ( n18775 & n18824 ) ;
  assign n18831 = ( n7833 & n15308 ) | ( n7833 & n18829 ) | ( n15308 & n18829 ) ;
  assign n18832 = n7829 & ~n15320 ;
  assign n18833 = ( n7834 & n15322 ) | ( n7834 & n18832 ) | ( n15322 & n18832 ) ;
  assign n18834 = n18829 | n18831 ;
  assign n18835 = ( n7834 & ~n15320 ) | ( n7834 & n18829 ) | ( ~n15320 & n18829 ) ;
  assign n18836 = n18834 | n18835 ;
  assign n18837 = n7838 & ~n18552 ;
  assign n18838 = n18836 | n18837 ;
  assign n18839 = ( n7833 & n15319 ) | ( n7833 & n18832 ) | ( n15319 & n18832 ) ;
  assign n18840 = n18832 | n18839 ;
  assign n18841 = n7838 & ~n18550 ;
  assign n18842 = n7829 & n15308 ;
  assign n18843 = ( n7834 & n15319 ) | ( n7834 & n18842 ) | ( n15319 & n18842 ) ;
  assign n18844 = n18833 | n18840 ;
  assign n18845 = n18841 | n18844 ;
  assign n18846 = ( n7833 & n15312 ) | ( n7833 & n18842 ) | ( n15312 & n18842 ) ;
  assign n18847 = n18842 | n18846 ;
  assign n18848 = n7838 & n18531 ;
  assign n18849 = n18843 | n18847 ;
  assign n18850 = n18848 | n18849 ;
  assign n18851 = n18850 ^ x11 ^ 1'b0 ;
  assign n18852 = ( n18794 & n18814 ) | ( n18794 & n18851 ) | ( n18814 & n18851 ) ;
  assign n18853 = n18851 ^ n18814 ^ n18794 ;
  assign n18854 = n18853 ^ n18823 ^ n18776 ;
  assign n18855 = n18854 ^ n18830 ^ 1'b0 ;
  assign n18856 = ( n18827 & n18830 ) | ( n18827 & n18854 ) | ( n18830 & n18854 ) ;
  assign n18857 = n18855 ^ n18827 ^ 1'b0 ;
  assign n18858 = ( n18776 & n18823 ) | ( n18776 & n18853 ) | ( n18823 & n18853 ) ;
  assign n18859 = n7188 & ~n15032 ;
  assign n18860 = ( n7190 & ~n14970 ) | ( n7190 & n18859 ) | ( ~n14970 & n18859 ) ;
  assign n18861 = n18859 | n18860 ;
  assign n18862 = ( n7192 & n15001 ) | ( n7192 & n18859 ) | ( n15001 & n18859 ) ;
  assign n18863 = n18861 | n18862 ;
  assign n18864 = n7196 & ~n18085 ;
  assign n18865 = n18863 | n18864 ;
  assign n18866 = n18865 ^ x23 ^ 1'b0 ;
  assign n18867 = ( n17687 & ~n17888 ) | ( n17687 & n18866 ) | ( ~n17888 & n18866 ) ;
  assign n18868 = n18866 ^ n17888 ^ n17687 ;
  assign n18869 = n7188 & ~n15095 ;
  assign n18870 = ( n7190 & n15001 ) | ( n7190 & n18869 ) | ( n15001 & n18869 ) ;
  assign n18871 = n18869 | n18870 ;
  assign n18872 = ( n7192 & ~n15032 ) | ( n7192 & n18869 ) | ( ~n15032 & n18869 ) ;
  assign n18873 = n18871 | n18872 ;
  assign n18874 = n7196 & n18108 ;
  assign n18875 = n18873 | n18874 ;
  assign n18876 = n18875 ^ x23 ^ 1'b0 ;
  assign n18877 = n18876 ^ n18867 ^ n17902 ;
  assign n18878 = ( ~n17902 & n18867 ) | ( ~n17902 & n18876 ) | ( n18867 & n18876 ) ;
  assign n18879 = n7339 & ~n15216 ;
  assign n18880 = ( n7337 & n15218 ) | ( n7337 & n18879 ) | ( n15218 & n18879 ) ;
  assign n18881 = n18879 | n18880 ;
  assign n18882 = ( n7338 & ~n15095 ) | ( n7338 & n18879 ) | ( ~n15095 & n18879 ) ;
  assign n18883 = n18881 | n18882 ;
  assign n18884 = n7340 & n18200 ;
  assign n18885 = n18883 | n18884 ;
  assign n18886 = n18885 ^ x20 ^ 1'b0 ;
  assign n18887 = n18886 ^ n18868 ^ n18023 ;
  assign n18888 = ( n18023 & ~n18868 ) | ( n18023 & n18886 ) | ( ~n18868 & n18886 ) ;
  assign n18889 = n7485 & n15239 ;
  assign n18890 = ( n7486 & ~n15248 ) | ( n7486 & n18889 ) | ( ~n15248 & n18889 ) ;
  assign n18891 = n18889 | n18890 ;
  assign n18892 = ( n7493 & n15219 ) | ( n7493 & n18889 ) | ( n15219 & n18889 ) ;
  assign n18893 = n18891 | n18892 ;
  assign n18894 = n7487 & ~n18303 ;
  assign n18895 = n18893 | n18894 ;
  assign n18896 = n18895 ^ x17 ^ 1'b0 ;
  assign n18897 = n18896 ^ n18887 ^ n18708 ;
  assign n18898 = ( n18708 & ~n18887 ) | ( n18708 & n18896 ) | ( ~n18887 & n18896 ) ;
  assign n18899 = n7669 & ~n15275 ;
  assign n18900 = ( n7674 & n15271 ) | ( n7674 & n18899 ) | ( n15271 & n18899 ) ;
  assign n18901 = n18899 | n18900 ;
  assign n18902 = ( n7667 & n15312 ) | ( n7667 & n18899 ) | ( n15312 & n18899 ) ;
  assign n18903 = n18901 | n18902 ;
  assign n18904 = n7666 & ~n18480 ;
  assign n18905 = n18903 | n18904 ;
  assign n18906 = n18905 ^ x14 ^ 1'b0 ;
  assign n18907 = n18906 ^ n18897 ^ n18803 ;
  assign n18908 = n18838 ^ x11 ^ 1'b0 ;
  assign n18909 = n18845 ^ x11 ^ 1'b0 ;
  assign n18910 = ( n18803 & ~n18897 ) | ( n18803 & n18906 ) | ( ~n18897 & n18906 ) ;
  assign n18911 = n18908 ^ n18907 ^ n18813 ;
  assign n18912 = n7487 & ~n18354 ;
  assign n18913 = ( n18813 & ~n18907 ) | ( n18813 & n18908 ) | ( ~n18907 & n18908 ) ;
  assign n18914 = n7485 & ~n15248 ;
  assign n18915 = ( n7486 & n15271 ) | ( n7486 & n18914 ) | ( n15271 & n18914 ) ;
  assign n18916 = n18914 | n18915 ;
  assign n18917 = ( n7493 & n15239 ) | ( n7493 & n18914 ) | ( n15239 & n18914 ) ;
  assign n18918 = n18916 | n18917 ;
  assign n18919 = n18912 | n18918 ;
  assign n18920 = ( x8 & n18852 ) | ( x8 & ~n18911 ) | ( n18852 & ~n18911 ) ;
  assign n18921 = n18911 ^ n18852 ^ x8 ;
  assign n18922 = n18921 ^ n18858 ^ 1'b0 ;
  assign n18923 = ( n18856 & n18858 ) | ( n18856 & ~n18921 ) | ( n18858 & ~n18921 ) ;
  assign n18924 = n7339 & n15218 ;
  assign n18925 = ( n7338 & ~n15216 ) | ( n7338 & n18924 ) | ( ~n15216 & n18924 ) ;
  assign n18926 = n18922 ^ n18856 ^ 1'b0 ;
  assign n18927 = ( n7337 & n15219 ) | ( n7337 & n18924 ) | ( n15219 & n18924 ) ;
  assign n18928 = n18924 | n18927 ;
  assign n18929 = n7340 & ~n18252 ;
  assign n18930 = n18925 | n18928 ;
  assign n18931 = n18929 | n18930 ;
  assign n18932 = n18931 ^ x20 ^ 1'b0 ;
  assign n18933 = ( ~n18877 & n18888 ) | ( ~n18877 & n18932 ) | ( n18888 & n18932 ) ;
  assign n18934 = n18919 ^ x17 ^ 1'b0 ;
  assign n18935 = n18932 ^ n18888 ^ n18877 ;
  assign n18936 = n18935 ^ n18934 ^ n18898 ;
  assign n18937 = ( n18898 & n18934 ) | ( n18898 & ~n18935 ) | ( n18934 & ~n18935 ) ;
  assign n18938 = n7669 & n15312 ;
  assign n18939 = ( n7674 & ~n15275 ) | ( n7674 & n18938 ) | ( ~n15275 & n18938 ) ;
  assign n18940 = n18938 | n18939 ;
  assign n18941 = ( n7667 & n15308 ) | ( n7667 & n18938 ) | ( n15308 & n18938 ) ;
  assign n18942 = n18940 | n18941 ;
  assign n18943 = n7666 & n18525 ;
  assign n18944 = n18942 | n18943 ;
  assign n18945 = n18944 ^ x14 ^ 1'b0 ;
  assign n18946 = n18945 ^ n18936 ^ n18910 ;
  assign n18947 = ( n18910 & ~n18936 ) | ( n18910 & n18945 ) | ( ~n18936 & n18945 ) ;
  assign n18948 = n7669 & n15319 ;
  assign n18949 = ( n7674 & n15308 ) | ( n7674 & n18948 ) | ( n15308 & n18948 ) ;
  assign n18950 = n18948 | n18949 ;
  assign n18951 = ( n7667 & ~n15320 ) | ( n7667 & n18948 ) | ( ~n15320 & n18948 ) ;
  assign n18952 = n18950 | n18951 ;
  assign n18953 = n7666 & ~n18552 ;
  assign n18954 = n18952 | n18953 ;
  assign n18955 = n18946 ^ n18913 ^ n18909 ;
  assign n18956 = ( n18909 & n18913 ) | ( n18909 & ~n18946 ) | ( n18913 & ~n18946 ) ;
  assign n18957 = n7669 & n15308 ;
  assign n18958 = ( n7674 & n15312 ) | ( n7674 & n18957 ) | ( n15312 & n18957 ) ;
  assign n18959 = n18957 | n18958 ;
  assign n18960 = n7833 & ~n15320 ;
  assign n18961 = ( n7667 & n15319 ) | ( n7667 & n18957 ) | ( n15319 & n18957 ) ;
  assign n18962 = n18955 ^ n18920 ^ 1'b0 ;
  assign n18963 = n18959 | n18961 ;
  assign n18964 = n18962 ^ n18923 ^ 1'b0 ;
  assign n18965 = ( n18920 & n18923 ) | ( n18920 & ~n18955 ) | ( n18923 & ~n18955 ) ;
  assign n18966 = n7485 & n15271 ;
  assign n18967 = ( n7486 & ~n15275 ) | ( n7486 & n18966 ) | ( ~n15275 & n18966 ) ;
  assign n18968 = n18966 | n18967 ;
  assign n18969 = ( n7493 & ~n15248 ) | ( n7493 & n18966 ) | ( ~n15248 & n18966 ) ;
  assign n18970 = n7487 & ~n18456 ;
  assign n18971 = n18968 | n18969 ;
  assign n18972 = n18970 | n18971 ;
  assign n18973 = n7188 & ~n15216 ;
  assign n18974 = ( n7190 & ~n15032 ) | ( n7190 & n18973 ) | ( ~n15032 & n18973 ) ;
  assign n18975 = n18972 ^ x17 ^ 1'b0 ;
  assign n18976 = n18973 | n18974 ;
  assign n18977 = ( n7192 & ~n15095 ) | ( n7192 & n18973 ) | ( ~n15095 & n18973 ) ;
  assign n18978 = n18976 | n18977 ;
  assign n18979 = n7196 & ~n18158 ;
  assign n18980 = n18978 | n18979 ;
  assign n18981 = n18980 ^ x23 ^ 1'b0 ;
  assign n18982 = n18981 ^ n18062 ^ n17901 ;
  assign n18983 = ( n17901 & ~n18062 ) | ( n17901 & n18981 ) | ( ~n18062 & n18981 ) ;
  assign n18984 = n7666 & n18531 ;
  assign n18985 = n7339 & n15219 ;
  assign n18986 = n18963 | n18984 ;
  assign n18987 = n18986 ^ x14 ^ 1'b0 ;
  assign n18988 = n7669 & ~n15320 ;
  assign n18989 = n18960 ^ x11 ^ 1'b0 ;
  assign n18990 = ( n7666 & ~n18550 ) | ( n7666 & n18988 ) | ( ~n18550 & n18988 ) ;
  assign n18991 = ( n7337 & n15239 ) | ( n7337 & n18985 ) | ( n15239 & n18985 ) ;
  assign n18992 = n18985 | n18991 ;
  assign n18993 = ( n7338 & n15218 ) | ( n7338 & n18985 ) | ( n15218 & n18985 ) ;
  assign n18994 = n18992 | n18993 ;
  assign n18995 = n7340 & n18272 ;
  assign n18996 = n18994 | n18995 ;
  assign n18997 = n18996 ^ x20 ^ 1'b0 ;
  assign n18998 = ( n18878 & ~n18982 ) | ( n18878 & n18997 ) | ( ~n18982 & n18997 ) ;
  assign n18999 = n18997 ^ n18982 ^ n18878 ;
  assign n19000 = ( n18933 & n18975 ) | ( n18933 & ~n18999 ) | ( n18975 & ~n18999 ) ;
  assign n19001 = n18999 ^ n18975 ^ n18933 ;
  assign n19002 = ( n18937 & n18987 ) | ( n18937 & ~n19001 ) | ( n18987 & ~n19001 ) ;
  assign n19003 = n19001 ^ n18987 ^ n18937 ;
  assign n19004 = ( n18947 & n18989 ) | ( n18947 & ~n19003 ) | ( n18989 & ~n19003 ) ;
  assign n19005 = n19003 ^ n18989 ^ n18947 ;
  assign n19006 = n19005 ^ n18956 ^ 1'b0 ;
  assign n19007 = n19006 ^ n18965 ^ 1'b0 ;
  assign n19008 = ( n18956 & n18965 ) | ( n18956 & ~n19005 ) | ( n18965 & ~n19005 ) ;
  assign n19009 = ( n7674 & n15319 ) | ( n7674 & n18988 ) | ( n15319 & n18988 ) ;
  assign n19010 = n18988 | n19009 ;
  assign n19011 = n7037 & ~n15032 ;
  assign n19012 = n18990 | n19010 ;
  assign n19013 = ( n7036 & n15001 ) | ( n7036 & n19011 ) | ( n15001 & n19011 ) ;
  assign n19014 = n19011 | n19013 ;
  assign n19015 = ( n7052 & ~n14970 ) | ( n7052 & n19011 ) | ( ~n14970 & n19011 ) ;
  assign n19016 = n19014 | n19015 ;
  assign n19017 = n7035 & ~n18085 ;
  assign n19018 = n19016 | n19017 ;
  assign n19019 = n19018 ^ x26 ^ 1'b0 ;
  assign n19020 = ( n17717 & n17816 ) | ( n17717 & n19019 ) | ( n17816 & n19019 ) ;
  assign n19021 = n19019 ^ n17816 ^ n17717 ;
  assign n19022 = n7188 & n15218 ;
  assign n19023 = ( n7190 & ~n15095 ) | ( n7190 & n19022 ) | ( ~n15095 & n19022 ) ;
  assign n19024 = n18954 ^ x14 ^ 1'b0 ;
  assign n19025 = n19022 | n19023 ;
  assign n19026 = ( n7192 & ~n15216 ) | ( n7192 & n19022 ) | ( ~n15216 & n19022 ) ;
  assign n19027 = n19012 ^ x14 ^ 1'b0 ;
  assign n19028 = n19025 | n19026 ;
  assign n19029 = n7196 & n18200 ;
  assign n19030 = n19028 | n19029 ;
  assign n19031 = n19030 ^ x23 ^ 1'b0 ;
  assign n19032 = ( n18063 & n19021 ) | ( n18063 & n19031 ) | ( n19021 & n19031 ) ;
  assign n19033 = n19031 ^ n19021 ^ n18063 ;
  assign n19034 = n7339 & n15239 ;
  assign n19035 = ( n7337 & ~n15248 ) | ( n7337 & n19034 ) | ( ~n15248 & n19034 ) ;
  assign n19036 = n19034 | n19035 ;
  assign n19037 = ( n7338 & n15219 ) | ( n7338 & n19034 ) | ( n15219 & n19034 ) ;
  assign n19038 = n19036 | n19037 ;
  assign n19039 = n18016 ^ n6650 ^ 1'b0 ;
  assign n19040 = n19039 ^ n18087 ^ 1'b0 ;
  assign n19041 = ( n6650 & ~n18016 ) | ( n6650 & n18087 ) | ( ~n18016 & n18087 ) ;
  assign n19042 = n7340 & ~n18303 ;
  assign n19043 = n19038 | n19042 ;
  assign n19044 = n19043 ^ x20 ^ 1'b0 ;
  assign n19045 = n19044 ^ n19033 ^ n18983 ;
  assign n19046 = ( n18983 & n19033 ) | ( n18983 & n19044 ) | ( n19033 & n19044 ) ;
  assign n19047 = n7485 & ~n15275 ;
  assign n19048 = ( n7486 & n15312 ) | ( n7486 & n19047 ) | ( n15312 & n19047 ) ;
  assign n19049 = n19047 | n19048 ;
  assign n19050 = ( n7493 & n15271 ) | ( n7493 & n19047 ) | ( n15271 & n19047 ) ;
  assign n19051 = n19049 | n19050 ;
  assign n19052 = n7487 & ~n18480 ;
  assign n19053 = n19051 | n19052 ;
  assign n19054 = n19053 ^ x17 ^ 1'b0 ;
  assign n19055 = n19054 ^ n19045 ^ n18998 ;
  assign n19056 = ( n18998 & n19045 ) | ( n18998 & n19054 ) | ( n19045 & n19054 ) ;
  assign n19057 = n19055 ^ n19024 ^ n19000 ;
  assign n19058 = n19057 ^ n19002 ^ x11 ;
  assign n19059 = ( x11 & n19002 ) | ( x11 & n19057 ) | ( n19002 & n19057 ) ;
  assign n19060 = n19058 ^ n19004 ^ 1'b0 ;
  assign n19061 = ( n19004 & n19008 ) | ( n19004 & n19058 ) | ( n19008 & n19058 ) ;
  assign n19062 = n19060 ^ n19008 ^ 1'b0 ;
  assign n19063 = n6901 & ~n15032 ;
  assign n19064 = ( n6906 & n15001 ) | ( n6906 & n19063 ) | ( n15001 & n19063 ) ;
  assign n19065 = n19063 | n19064 ;
  assign n19066 = ( n19000 & n19024 ) | ( n19000 & n19055 ) | ( n19024 & n19055 ) ;
  assign n19067 = ( n6907 & ~n15095 ) | ( n6907 & n19063 ) | ( ~n15095 & n19063 ) ;
  assign n19068 = n6918 & n18108 ;
  assign n19069 = n19065 | n19067 ;
  assign n19070 = n19068 | n19069 ;
  assign n19071 = n19070 ^ x29 ^ 1'b0 ;
  assign n19072 = ( n17800 & ~n18007 ) | ( n17800 & n19071 ) | ( ~n18007 & n19071 ) ;
  assign n19073 = n19071 ^ n18007 ^ n17800 ;
  assign n19074 = n7037 & ~n15095 ;
  assign n19075 = ( n7036 & ~n15032 ) | ( n7036 & n19074 ) | ( ~n15032 & n19074 ) ;
  assign n19076 = n19074 | n19075 ;
  assign n19077 = ( n7052 & n15001 ) | ( n7052 & n19074 ) | ( n15001 & n19074 ) ;
  assign n19078 = n19076 | n19077 ;
  assign n19079 = n7035 & n18108 ;
  assign n19080 = n19078 | n19079 ;
  assign n19081 = n19080 ^ x26 ^ 1'b0 ;
  assign n19082 = ( ~n18010 & n19020 ) | ( ~n18010 & n19081 ) | ( n19020 & n19081 ) ;
  assign n19083 = n19081 ^ n19020 ^ n18010 ;
  assign n19084 = n7188 & n15219 ;
  assign n19085 = ( n7190 & ~n15216 ) | ( n7190 & n19084 ) | ( ~n15216 & n19084 ) ;
  assign n19086 = n19084 | n19085 ;
  assign n19087 = ( n7192 & n15218 ) | ( n7192 & n19084 ) | ( n15218 & n19084 ) ;
  assign n19088 = n19086 | n19087 ;
  assign n19089 = n7196 & ~n18252 ;
  assign n19090 = n19088 | n19089 ;
  assign n19091 = n19090 ^ x23 ^ 1'b0 ;
  assign n19092 = ( n19032 & ~n19083 ) | ( n19032 & n19091 ) | ( ~n19083 & n19091 ) ;
  assign n19093 = n19091 ^ n19083 ^ n19032 ;
  assign n19094 = n7339 & ~n15248 ;
  assign n19095 = ( n7337 & n15271 ) | ( n7337 & n19094 ) | ( n15271 & n19094 ) ;
  assign n19096 = n19094 | n19095 ;
  assign n19097 = ( n7338 & n15239 ) | ( n7338 & n19094 ) | ( n15239 & n19094 ) ;
  assign n19098 = n19096 | n19097 ;
  assign n19099 = n7340 & ~n18354 ;
  assign n19100 = n19098 | n19099 ;
  assign n19101 = n19100 ^ x20 ^ 1'b0 ;
  assign n19102 = ( n19046 & ~n19093 ) | ( n19046 & n19101 ) | ( ~n19093 & n19101 ) ;
  assign n19103 = n19101 ^ n19093 ^ n19046 ;
  assign n19104 = n7485 & n15312 ;
  assign n19105 = ( n7486 & n15308 ) | ( n7486 & n19104 ) | ( n15308 & n19104 ) ;
  assign n19106 = n19104 | n19105 ;
  assign n19107 = ( n7493 & ~n15275 ) | ( n7493 & n19104 ) | ( ~n15275 & n19104 ) ;
  assign n19108 = n19106 | n19107 ;
  assign n19109 = n7487 & n18525 ;
  assign n19110 = n19108 | n19109 ;
  assign n19111 = n19110 ^ x17 ^ 1'b0 ;
  assign n19112 = ( n19056 & ~n19103 ) | ( n19056 & n19111 ) | ( ~n19103 & n19111 ) ;
  assign n19113 = n19111 ^ n19103 ^ n19056 ;
  assign n19114 = n6791 & ~n15032 ;
  assign n19115 = ( n6788 & ~n15095 ) | ( n6788 & n19114 ) | ( ~n15095 & n19114 ) ;
  assign n19116 = n19114 | n19115 ;
  assign n19117 = ( n6790 & n15001 ) | ( n6790 & n19114 ) | ( n15001 & n19114 ) ;
  assign n19118 = n19116 | n19117 ;
  assign n19119 = ( ~x17 & n6785 ) | ( ~x17 & n6825 ) | ( n6785 & n6825 ) ;
  assign n19120 = n6789 & ~n18108 ;
  assign n19121 = ( n6789 & n19118 ) | ( n6789 & ~n19120 ) | ( n19118 & ~n19120 ) ;
  assign n19122 = n19041 ^ n6785 ^ n6650 ;
  assign n19123 = ( n6650 & n6785 ) | ( n6650 & ~n19041 ) | ( n6785 & ~n19041 ) ;
  assign n19124 = ( n19027 & n19066 ) | ( n19027 & ~n19113 ) | ( n19066 & ~n19113 ) ;
  assign n19125 = n6825 ^ n6785 ^ x17 ;
  assign n19126 = n19113 ^ n19066 ^ n19027 ;
  assign n19127 = ( ~n19121 & n19123 ) | ( ~n19121 & n19125 ) | ( n19123 & n19125 ) ;
  assign n19128 = n19126 ^ n19059 ^ 1'b0 ;
  assign n19129 = n19128 ^ n19061 ^ 1'b0 ;
  assign n19130 = ( n19059 & n19061 ) | ( n19059 & ~n19126 ) | ( n19061 & ~n19126 ) ;
  assign n19131 = n19125 ^ n19123 ^ n19121 ;
  assign n19132 = n7037 & ~n15216 ;
  assign n19133 = ( n7036 & ~n15095 ) | ( n7036 & n19132 ) | ( ~n15095 & n19132 ) ;
  assign n19134 = n19132 | n19133 ;
  assign n19135 = ( n7052 & ~n15032 ) | ( n7052 & n19132 ) | ( ~n15032 & n19132 ) ;
  assign n19136 = n19134 | n19135 ;
  assign n19137 = n7035 & ~n18158 ;
  assign n19138 = n19136 | n19137 ;
  assign n19139 = n19138 ^ x26 ^ 1'b0 ;
  assign n19140 = n19139 ^ n18011 ^ n17789 ;
  assign n19141 = ( n17789 & n18011 ) | ( n17789 & n19139 ) | ( n18011 & n19139 ) ;
  assign n19142 = n7188 & n15239 ;
  assign n19143 = ( n7190 & n15218 ) | ( n7190 & n19142 ) | ( n15218 & n19142 ) ;
  assign n19144 = n19142 | n19143 ;
  assign n19145 = ( n7192 & n15219 ) | ( n7192 & n19142 ) | ( n15219 & n19142 ) ;
  assign n19146 = n19144 | n19145 ;
  assign n19147 = n7196 & n18272 ;
  assign n19148 = n19146 | n19147 ;
  assign n19149 = n19148 ^ x23 ^ 1'b0 ;
  assign n19150 = ( n19082 & n19140 ) | ( n19082 & n19149 ) | ( n19140 & n19149 ) ;
  assign n19151 = n19149 ^ n19140 ^ n19082 ;
  assign n19152 = n7339 & n15271 ;
  assign n19153 = ( n7337 & ~n15275 ) | ( n7337 & n19152 ) | ( ~n15275 & n19152 ) ;
  assign n19154 = n19152 | n19153 ;
  assign n19155 = ( n7338 & ~n15248 ) | ( n7338 & n19152 ) | ( ~n15248 & n19152 ) ;
  assign n19156 = n19154 | n19155 ;
  assign n19157 = n7340 & ~n18456 ;
  assign n19158 = n19156 | n19157 ;
  assign n19159 = n19158 ^ x20 ^ 1'b0 ;
  assign n19160 = n19159 ^ n19151 ^ n19092 ;
  assign n19161 = ( n19092 & n19151 ) | ( n19092 & n19159 ) | ( n19151 & n19159 ) ;
  assign n19162 = n7485 & n15308 ;
  assign n19163 = ( n7486 & n15319 ) | ( n7486 & n19162 ) | ( n15319 & n19162 ) ;
  assign n19164 = n19162 | n19163 ;
  assign n19165 = ( n7493 & n15312 ) | ( n7493 & n19162 ) | ( n15312 & n19162 ) ;
  assign n19166 = n19164 | n19165 ;
  assign n19167 = n7487 & n18531 ;
  assign n19168 = n19166 | n19167 ;
  assign n19169 = n19168 ^ x17 ^ 1'b0 ;
  assign n19170 = ( n19102 & n19160 ) | ( n19102 & n19169 ) | ( n19160 & n19169 ) ;
  assign n19171 = n19169 ^ n19160 ^ n19102 ;
  assign n19172 = n7674 & ~n15320 ;
  assign n19173 = n19172 ^ x14 ^ 1'b0 ;
  assign n19174 = ( n19112 & n19171 ) | ( n19112 & n19173 ) | ( n19171 & n19173 ) ;
  assign n19175 = n19173 ^ n19171 ^ n19112 ;
  assign n19176 = n7485 & n15319 ;
  assign n19177 = ( n7486 & ~n15320 ) | ( n7486 & n19176 ) | ( ~n15320 & n19176 ) ;
  assign n19178 = n19176 | n19177 ;
  assign n19179 = ( n7493 & n15308 ) | ( n7493 & n19176 ) | ( n15308 & n19176 ) ;
  assign n19180 = n19178 | n19179 ;
  assign n19181 = n7487 & ~n18550 ;
  assign n19182 = n7487 & ~n18552 ;
  assign n19183 = n19180 | n19182 ;
  assign n19184 = n19175 ^ n19124 ^ 1'b0 ;
  assign n19185 = n19184 ^ n19130 ^ 1'b0 ;
  assign n19186 = ( n19124 & n19130 ) | ( n19124 & n19175 ) | ( n19130 & n19175 ) ;
  assign n19187 = n7485 & n15322 ;
  assign n19188 = ( n7493 & ~n15320 ) | ( n7493 & n19187 ) | ( ~n15320 & n19187 ) ;
  assign n19189 = n7485 & ~n15320 ;
  assign n19190 = ( n7493 & n15319 ) | ( n7493 & n19189 ) | ( n15319 & n19189 ) ;
  assign n19191 = ( n7486 & n15322 ) | ( n7486 & n19189 ) | ( n15322 & n19189 ) ;
  assign n19192 = n19189 | n19191 ;
  assign n19193 = n19190 | n19192 ;
  assign n19194 = n19187 | n19188 ;
  assign n19195 = n19181 | n19193 ;
  assign n19196 = n6791 & n15001 ;
  assign n19197 = ( n6788 & ~n15032 ) | ( n6788 & n19196 ) | ( ~n15032 & n19196 ) ;
  assign n19198 = n19196 | n19197 ;
  assign n19199 = ( n6790 & ~n14970 ) | ( n6790 & n19196 ) | ( ~n14970 & n19196 ) ;
  assign n19200 = n6901 & n15001 ;
  assign n19201 = ( n6906 & ~n14970 ) | ( n6906 & n19200 ) | ( ~n14970 & n19200 ) ;
  assign n19202 = n19198 | n19199 ;
  assign n19203 = n19200 | n19201 ;
  assign n19204 = n6789 & ~n18085 ;
  assign n19205 = ( n6907 & ~n15032 ) | ( n6907 & n19200 ) | ( ~n15032 & n19200 ) ;
  assign n19206 = n19203 | n19205 ;
  assign n19207 = n7037 & n15218 ;
  assign n19208 = n6918 & ~n18085 ;
  assign n19209 = n19206 | n19208 ;
  assign n19210 = ( n7036 & ~n15216 ) | ( n7036 & n19207 ) | ( ~n15216 & n19207 ) ;
  assign n19211 = n19207 | n19210 ;
  assign n19212 = n19202 | n19204 ;
  assign n19213 = ( n7052 & ~n15095 ) | ( n7052 & n19207 ) | ( ~n15095 & n19207 ) ;
  assign n19214 = n19211 | n19213 ;
  assign n19215 = n7035 & n18200 ;
  assign n19216 = n19214 | n19215 ;
  assign n19217 = n19209 ^ x29 ^ 1'b0 ;
  assign n19218 = n19216 ^ x26 ^ 1'b0 ;
  assign n19219 = ( ~n17801 & n19217 ) | ( ~n17801 & n19218 ) | ( n19217 & n19218 ) ;
  assign n19220 = n7339 & ~n15275 ;
  assign n19221 = n7674 & n15322 ;
  assign n19222 = n19221 ^ x14 ^ 1'b0 ;
  assign n19223 = n19218 ^ n19217 ^ n17801 ;
  assign n19224 = n7188 & ~n15248 ;
  assign n19225 = ( n7337 & n15312 ) | ( n7337 & n19220 ) | ( n15312 & n19220 ) ;
  assign n19226 = n19220 | n19225 ;
  assign n19227 = ( n7338 & n15271 ) | ( n7338 & n19220 ) | ( n15271 & n19220 ) ;
  assign n19228 = n19226 | n19227 ;
  assign n19229 = n7340 & ~n18480 ;
  assign n19230 = n19183 ^ x17 ^ 1'b0 ;
  assign n19231 = n19228 | n19229 ;
  assign n19232 = ( n7190 & n15219 ) | ( n7190 & n19224 ) | ( n15219 & n19224 ) ;
  assign n19233 = n19224 | n19232 ;
  assign n19234 = ( n7192 & n15239 ) | ( n7192 & n19224 ) | ( n15239 & n19224 ) ;
  assign n19235 = n19231 ^ x20 ^ 1'b0 ;
  assign n19236 = n19233 | n19234 ;
  assign n19237 = n7196 & ~n18303 ;
  assign n19238 = n19236 | n19237 ;
  assign n19239 = n19238 ^ x23 ^ 1'b0 ;
  assign n19240 = ( n19141 & ~n19223 ) | ( n19141 & n19239 ) | ( ~n19223 & n19239 ) ;
  assign n19241 = n19239 ^ n19223 ^ n19141 ;
  assign n19242 = ( n19150 & n19235 ) | ( n19150 & ~n19241 ) | ( n19235 & ~n19241 ) ;
  assign n19243 = n19241 ^ n19235 ^ n19150 ;
  assign n19244 = n19243 ^ n19230 ^ n19161 ;
  assign n19245 = ( n19170 & n19222 ) | ( n19170 & ~n19244 ) | ( n19222 & ~n19244 ) ;
  assign n19246 = ( n19161 & n19230 ) | ( n19161 & ~n19243 ) | ( n19230 & ~n19243 ) ;
  assign n19247 = n19244 ^ n19222 ^ n19170 ;
  assign n19248 = n19247 ^ n19174 ^ 1'b0 ;
  assign n19249 = ( n19174 & n19186 ) | ( n19174 & ~n19247 ) | ( n19186 & ~n19247 ) ;
  assign n19250 = n19248 ^ n19186 ^ 1'b0 ;
  assign n19251 = n7037 & n15219 ;
  assign n19252 = ( n7036 & n15218 ) | ( n7036 & n19251 ) | ( n15218 & n19251 ) ;
  assign n19253 = n19251 | n19252 ;
  assign n19254 = ( n7052 & ~n15216 ) | ( n7052 & n19251 ) | ( ~n15216 & n19251 ) ;
  assign n19255 = n19253 | n19254 ;
  assign n19256 = n7035 & ~n18252 ;
  assign n19257 = n19255 | n19256 ;
  assign n19258 = n19257 ^ x26 ^ 1'b0 ;
  assign n19259 = ( ~n19073 & n19219 ) | ( ~n19073 & n19258 ) | ( n19219 & n19258 ) ;
  assign n19260 = n19258 ^ n19219 ^ n19073 ;
  assign n19261 = n6791 & ~n15095 ;
  assign n19262 = ( n6788 & ~n15216 ) | ( n6788 & n19261 ) | ( ~n15216 & n19261 ) ;
  assign n19263 = n19261 | n19262 ;
  assign n19264 = ( n6790 & ~n15032 ) | ( n6790 & n19261 ) | ( ~n15032 & n19261 ) ;
  assign n19265 = n19263 | n19264 ;
  assign n19266 = n6901 & ~n15095 ;
  assign n19267 = ( n6906 & ~n15032 ) | ( n6906 & n19266 ) | ( ~n15032 & n19266 ) ;
  assign n19268 = n19266 | n19267 ;
  assign n19269 = ( n6907 & ~n15216 ) | ( n6907 & n19266 ) | ( ~n15216 & n19266 ) ;
  assign n19270 = n19268 | n19269 ;
  assign n19271 = n6789 & ~n18158 ;
  assign n19272 = n6918 & ~n18158 ;
  assign n19273 = n19265 | n19271 ;
  assign n19274 = n19270 & ~n19272 ;
  assign n19275 = n7188 & n15271 ;
  assign n19276 = n19274 ^ n19272 ^ x29 ;
  assign n19277 = ( n7190 & n15239 ) | ( n7190 & n19275 ) | ( n15239 & n19275 ) ;
  assign n19278 = n19275 | n19277 ;
  assign n19279 = ( n7192 & ~n15248 ) | ( n7192 & n19275 ) | ( ~n15248 & n19275 ) ;
  assign n19280 = n19278 | n19279 ;
  assign n19281 = n7196 & ~n18354 ;
  assign n19282 = n19280 | n19281 ;
  assign n19283 = n19282 ^ x23 ^ 1'b0 ;
  assign n19284 = n19283 ^ n19260 ^ n19240 ;
  assign n19285 = ( n19240 & ~n19260 ) | ( n19240 & n19283 ) | ( ~n19260 & n19283 ) ;
  assign n19286 = n7339 & n15312 ;
  assign n19287 = ( n7337 & n15308 ) | ( n7337 & n19286 ) | ( n15308 & n19286 ) ;
  assign n19288 = n19286 | n19287 ;
  assign n19289 = ( n7338 & ~n15275 ) | ( n7338 & n19286 ) | ( ~n15275 & n19286 ) ;
  assign n19290 = n19288 | n19289 ;
  assign n19291 = n7340 & n18525 ;
  assign n19292 = n19290 | n19291 ;
  assign n19293 = n19195 ^ x17 ^ 1'b0 ;
  assign n19294 = n19292 ^ x20 ^ 1'b0 ;
  assign n19295 = n19294 ^ n19284 ^ n19242 ;
  assign n19296 = ( n19242 & ~n19284 ) | ( n19242 & n19294 ) | ( ~n19284 & n19294 ) ;
  assign n19297 = ( n19246 & n19293 ) | ( n19246 & ~n19295 ) | ( n19293 & ~n19295 ) ;
  assign n19298 = n19295 ^ n19293 ^ n19246 ;
  assign n19299 = n19298 ^ n19245 ^ 1'b0 ;
  assign n19300 = ( n19245 & n19249 ) | ( n19245 & ~n19298 ) | ( n19249 & ~n19298 ) ;
  assign n19301 = n19299 ^ n19249 ^ 1'b0 ;
  assign n19302 = n18493 ^ n18461 ^ 1'b0 ;
  assign n19303 = n18461 | n18493 ;
  assign n19304 = ( n18006 & ~n19040 ) | ( n18006 & n19276 ) | ( ~n19040 & n19276 ) ;
  assign n19305 = n19276 ^ n19040 ^ n18006 ;
  assign n19306 = n6901 & ~n15216 ;
  assign n19307 = ( n6906 & ~n15095 ) | ( n6906 & n19306 ) | ( ~n15095 & n19306 ) ;
  assign n19308 = n19306 | n19307 ;
  assign n19309 = ( n6907 & n15218 ) | ( n6907 & n19306 ) | ( n15218 & n19306 ) ;
  assign n19310 = n19308 | n19309 ;
  assign n19311 = n19303 ^ n18529 ^ 1'b0 ;
  assign n19312 = n18529 | n19303 ;
  assign n19313 = ( n6918 & n18200 ) | ( n6918 & n19310 ) | ( n18200 & n19310 ) ;
  assign n19314 = n19310 | n19313 ;
  assign n19315 = n18541 & ~n19312 ;
  assign n19316 = n19314 ^ x29 ^ 1'b0 ;
  assign n19317 = n19312 ^ n18541 ^ 1'b0 ;
  assign n19318 = n19315 ^ n18561 ^ 1'b0 ;
  assign n19319 = ~n18561 & n19315 ;
  assign n19320 = ~n18573 & n19319 ;
  assign n19321 = n19319 ^ n18573 ^ 1'b0 ;
  assign n19322 = n6789 & ~n18200 ;
  assign n19323 = n19316 ^ n19212 ^ n19122 ;
  assign n19324 = ( n19122 & n19212 ) | ( n19122 & n19316 ) | ( n19212 & n19316 ) ;
  assign n19325 = n6791 & ~n15216 ;
  assign n19326 = ( n6790 & ~n15095 ) | ( n6790 & n19325 ) | ( ~n15095 & n19325 ) ;
  assign n19327 = ( n6788 & n15218 ) | ( n6788 & n19325 ) | ( n15218 & n19325 ) ;
  assign n19328 = n19325 | n19327 ;
  assign n19329 = n6918 & ~n18252 ;
  assign n19330 = n6789 & ~n18252 ;
  assign n19331 = n19326 | n19328 ;
  assign n19332 = n6901 & n15218 ;
  assign n19333 = ( n6789 & ~n19322 ) | ( n6789 & n19331 ) | ( ~n19322 & n19331 ) ;
  assign n19334 = ( n6906 & ~n15216 ) | ( n6906 & n19332 ) | ( ~n15216 & n19332 ) ;
  assign n19335 = n19332 | n19334 ;
  assign n19336 = ( n6907 & n15219 ) | ( n6907 & n19332 ) | ( n15219 & n19332 ) ;
  assign n19337 = n19335 | n19336 ;
  assign n19338 = ( n6520 & ~n6705 ) | ( n6520 & n19333 ) | ( ~n6705 & n19333 ) ;
  assign n19339 = n19329 | n19337 ;
  assign n19340 = n6791 & n15218 ;
  assign n19341 = n19333 ^ n6705 ^ n6520 ;
  assign n19342 = ( n6788 & n15219 ) | ( n6788 & n19340 ) | ( n15219 & n19340 ) ;
  assign n19343 = n19340 | n19342 ;
  assign n19344 = ( n6790 & ~n15216 ) | ( n6790 & n19340 ) | ( ~n15216 & n19340 ) ;
  assign n19345 = ( x20 & n6520 ) | ( x20 & n6715 ) | ( n6520 & n6715 ) ;
  assign n19346 = n19339 ^ x29 ^ 1'b0 ;
  assign n19347 = n6715 ^ n6520 ^ x20 ;
  assign n19348 = n19343 | n19344 ;
  assign n19349 = n19346 ^ n19324 ^ n19131 ;
  assign n19350 = n19330 | n19348 ;
  assign n19351 = ( n19338 & ~n19347 ) | ( n19338 & n19350 ) | ( ~n19347 & n19350 ) ;
  assign n19352 = n19350 ^ n19347 ^ n19338 ;
  assign n19353 = n19119 ^ n6520 ^ 1'b0 ;
  assign n19354 = n19353 ^ n19273 ^ 1'b0 ;
  assign n19355 = n6901 & n15219 ;
  assign n19356 = ( n6520 & n19119 ) | ( n6520 & n19273 ) | ( n19119 & n19273 ) ;
  assign n19357 = ( n6906 & n15218 ) | ( n6906 & n19355 ) | ( n15218 & n19355 ) ;
  assign n19358 = ( n6907 & n15239 ) | ( n6907 & n19355 ) | ( n15239 & n19355 ) ;
  assign n19359 = n19355 | n19357 ;
  assign n19360 = ( n19131 & n19324 ) | ( n19131 & n19346 ) | ( n19324 & n19346 ) ;
  assign n19361 = n19358 | n19359 ;
  assign n19362 = ( n6918 & n18272 ) | ( n6918 & n19361 ) | ( n18272 & n19361 ) ;
  assign n19363 = n19361 | n19362 ;
  assign n19364 = n19363 ^ x29 ^ 1'b0 ;
  assign n19365 = ( ~n19127 & n19354 ) | ( ~n19127 & n19364 ) | ( n19354 & n19364 ) ;
  assign n19366 = n19365 ^ n19356 ^ n19341 ;
  assign n19367 = ( ~n19341 & n19356 ) | ( ~n19341 & n19365 ) | ( n19356 & n19365 ) ;
  assign n19368 = n19364 ^ n19354 ^ n19127 ;
  assign n19369 = n7037 & n15239 ;
  assign n19370 = ( n7036 & n15219 ) | ( n7036 & n19369 ) | ( n15219 & n19369 ) ;
  assign n19371 = n19369 | n19370 ;
  assign n19372 = ( n7052 & n15218 ) | ( n7052 & n19369 ) | ( n15218 & n19369 ) ;
  assign n19373 = n19371 | n19372 ;
  assign n19374 = n7035 & n18272 ;
  assign n19375 = n19373 | n19374 ;
  assign n19376 = n19375 ^ x26 ^ 1'b0 ;
  assign n19377 = ( n19072 & ~n19305 ) | ( n19072 & n19376 ) | ( ~n19305 & n19376 ) ;
  assign n19378 = n19376 ^ n19305 ^ n19072 ;
  assign n19379 = n6791 & n15219 ;
  assign n19380 = ( n6788 & n15239 ) | ( n6788 & n19379 ) | ( n15239 & n19379 ) ;
  assign n19381 = n19379 | n19380 ;
  assign n19382 = ( n6790 & n15218 ) | ( n6790 & n19379 ) | ( n15218 & n19379 ) ;
  assign n19383 = n19381 | n19382 ;
  assign n19384 = n7188 & ~n15275 ;
  assign n19385 = ( n7190 & ~n15248 ) | ( n7190 & n19384 ) | ( ~n15248 & n19384 ) ;
  assign n19386 = n6789 & ~n18272 ;
  assign n19387 = n19384 | n19385 ;
  assign n19388 = ( n7192 & n15271 ) | ( n7192 & n19384 ) | ( n15271 & n19384 ) ;
  assign n19389 = n19387 | n19388 ;
  assign n19390 = n7196 & ~n18456 ;
  assign n19391 = n19389 | n19390 ;
  assign n19392 = n19391 ^ x23 ^ 1'b0 ;
  assign n19393 = ( n6789 & n19383 ) | ( n6789 & ~n19386 ) | ( n19383 & ~n19386 ) ;
  assign n19394 = n19345 ^ n6702 ^ 1'b0 ;
  assign n19395 = ( n19259 & ~n19378 ) | ( n19259 & n19392 ) | ( ~n19378 & n19392 ) ;
  assign n19396 = ( n6702 & n19345 ) | ( n6702 & ~n19393 ) | ( n19345 & ~n19393 ) ;
  assign n19397 = n19392 ^ n19378 ^ n19259 ;
  assign n19398 = n7339 & n15308 ;
  assign n19399 = ( n7337 & n15319 ) | ( n7337 & n19398 ) | ( n15319 & n19398 ) ;
  assign n19400 = n19398 | n19399 ;
  assign n19401 = ( n7338 & n15312 ) | ( n7338 & n19398 ) | ( n15312 & n19398 ) ;
  assign n19402 = n19400 | n19401 ;
  assign n19403 = n7340 & n18531 ;
  assign n19404 = n19402 | n19403 ;
  assign n19405 = n19404 ^ x20 ^ 1'b0 ;
  assign n19406 = ( n19285 & ~n19397 ) | ( n19285 & n19405 ) | ( ~n19397 & n19405 ) ;
  assign n19407 = n19405 ^ n19397 ^ n19285 ;
  assign n19408 = n19396 ^ n6702 ^ n6451 ;
  assign n19409 = n6791 & ~n15248 ;
  assign n19410 = n19194 ^ x17 ^ 1'b0 ;
  assign n19411 = ( n6451 & n6702 ) | ( n6451 & ~n19396 ) | ( n6702 & ~n19396 ) ;
  assign n19412 = ( n6788 & n15271 ) | ( n6788 & n19409 ) | ( n15271 & n19409 ) ;
  assign n19413 = n19409 | n19412 ;
  assign n19414 = ( n6790 & n15239 ) | ( n6790 & n19409 ) | ( n15239 & n19409 ) ;
  assign n19415 = n19413 | n19414 ;
  assign n19416 = ( x23 & n6451 ) | ( x23 & n6652 ) | ( n6451 & n6652 ) ;
  assign n19417 = n6652 ^ n6451 ^ x23 ;
  assign n19418 = n6789 & ~n18354 ;
  assign n19419 = n19415 | n19418 ;
  assign n19420 = ( n19411 & ~n19417 ) | ( n19411 & n19419 ) | ( ~n19417 & n19419 ) ;
  assign n19421 = n19394 ^ n19393 ^ 1'b0 ;
  assign n19422 = ( n19296 & ~n19407 ) | ( n19296 & n19410 ) | ( ~n19407 & n19410 ) ;
  assign n19423 = n19410 ^ n19407 ^ n19296 ;
  assign n19424 = ( n19297 & n19300 ) | ( n19297 & ~n19423 ) | ( n19300 & ~n19423 ) ;
  assign n19425 = n19423 ^ n19297 ^ 1'b0 ;
  assign n19426 = n19425 ^ n19300 ^ 1'b0 ;
  assign n19427 = n19419 ^ n19417 ^ n19411 ;
  assign n19428 = n6791 & n15271 ;
  assign n19429 = ( n6788 & ~n15275 ) | ( n6788 & n19428 ) | ( ~n15275 & n19428 ) ;
  assign n19430 = n19428 | n19429 ;
  assign n19431 = ( n6790 & ~n15248 ) | ( n6790 & n19428 ) | ( ~n15248 & n19428 ) ;
  assign n19432 = n19430 | n19431 ;
  assign n19433 = n6789 & ~n18456 ;
  assign n19434 = n19432 | n19433 ;
  assign n19435 = ( n6654 & n19416 ) | ( n6654 & ~n19434 ) | ( n19416 & ~n19434 ) ;
  assign n19436 = n19416 ^ n6654 ^ 1'b0 ;
  assign n19437 = n19436 ^ n19434 ^ 1'b0 ;
  assign n19438 = n19435 ^ n6654 ^ n6290 ;
  assign n19439 = n6726 ^ n6654 ^ x26 ;
  assign n19440 = ( n6290 & n6654 ) | ( n6290 & n19435 ) | ( n6654 & n19435 ) ;
  assign n19441 = n6901 & n15308 ;
  assign n19442 = ( n6906 & n15312 ) | ( n6906 & n19441 ) | ( n15312 & n19441 ) ;
  assign n19443 = n19441 | n19442 ;
  assign n19444 = ( n6907 & n15319 ) | ( n6907 & n19441 ) | ( n15319 & n19441 ) ;
  assign n19445 = n19443 | n19444 ;
  assign n19446 = ( n6918 & n18531 ) | ( n6918 & n19445 ) | ( n18531 & n19445 ) ;
  assign n19447 = n19445 | n19446 ;
  assign n19448 = n19447 ^ x29 ^ 1'b0 ;
  assign n19449 = n19448 ^ n19437 ^ n19420 ;
  assign n19450 = ( n19420 & n19437 ) | ( n19420 & n19448 ) | ( n19437 & n19448 ) ;
  assign n19451 = n6791 & ~n15275 ;
  assign n19452 = ( n6788 & n15312 ) | ( n6788 & n19451 ) | ( n15312 & n19451 ) ;
  assign n19453 = n19451 | n19452 ;
  assign n19454 = ( n6790 & n15271 ) | ( n6790 & n19451 ) | ( n15271 & n19451 ) ;
  assign n19455 = n19453 | n19454 ;
  assign n19456 = n6789 & ~n18480 ;
  assign n19457 = n19455 | n19456 ;
  assign n19458 = n19457 ^ n19450 ^ n19438 ;
  assign n19459 = ( ~n19438 & n19450 ) | ( ~n19438 & n19457 ) | ( n19450 & n19457 ) ;
  assign n19460 = n6791 & n15239 ;
  assign n19461 = n6791 & n15312 ;
  assign n19462 = ( n6788 & ~n15248 ) | ( n6788 & n19460 ) | ( ~n15248 & n19460 ) ;
  assign n19463 = n19460 | n19462 ;
  assign n19464 = ( n6788 & n15308 ) | ( n6788 & n19461 ) | ( n15308 & n19461 ) ;
  assign n19465 = ( n6790 & n15219 ) | ( n6790 & n19460 ) | ( n15219 & n19460 ) ;
  assign n19466 = ( n6790 & ~n15275 ) | ( n6790 & n19461 ) | ( ~n15275 & n19461 ) ;
  assign n19467 = n19461 | n19464 ;
  assign n19468 = n6918 & ~n18550 ;
  assign n19469 = n19466 | n19467 ;
  assign n19470 = ( n6901 & ~n15320 ) | ( n6901 & n19468 ) | ( ~n15320 & n19468 ) ;
  assign n19471 = n19468 | n19470 ;
  assign n19472 = n19463 | n19465 ;
  assign n19473 = n6789 & ~n18525 ;
  assign n19474 = ( n6789 & n19469 ) | ( n6789 & ~n19473 ) | ( n19469 & ~n19473 ) ;
  assign n19475 = ( n6906 & n15319 ) | ( n6906 & n19468 ) | ( n15319 & n19468 ) ;
  assign n19476 = n19471 | n19475 ;
  assign n19477 = n6789 & ~n18303 ;
  assign n19478 = n19476 ^ n19459 ^ x29 ;
  assign n19479 = n19472 | n19477 ;
  assign n19480 = n19478 ^ n19474 ^ n19440 ;
  assign n19481 = n7037 & ~n15248 ;
  assign n19482 = ( n7036 & n15239 ) | ( n7036 & n19481 ) | ( n15239 & n19481 ) ;
  assign n19483 = n19481 | n19482 ;
  assign n19484 = ( n7052 & n15219 ) | ( n7052 & n19481 ) | ( n15219 & n19481 ) ;
  assign n19485 = n19483 | n19484 ;
  assign n19486 = n7035 & ~n18303 ;
  assign n19487 = n19485 | n19486 ;
  assign n19488 = n19487 ^ x26 ^ 1'b0 ;
  assign n19489 = ( n19304 & n19323 ) | ( n19304 & n19488 ) | ( n19323 & n19488 ) ;
  assign n19490 = n19488 ^ n19323 ^ n19304 ;
  assign n19491 = n6901 & ~n15248 ;
  assign n19492 = ( n6906 & n15239 ) | ( n6906 & n19491 ) | ( n15239 & n19491 ) ;
  assign n19493 = n19491 | n19492 ;
  assign n19494 = ( n6907 & n15271 ) | ( n6907 & n19491 ) | ( n15271 & n19491 ) ;
  assign n19495 = n19493 | n19494 ;
  assign n19496 = n6918 & ~n18354 ;
  assign n19497 = n19495 | n19496 ;
  assign n19498 = n19497 ^ x29 ^ 1'b0 ;
  assign n19499 = n19498 ^ n19367 ^ n19352 ;
  assign n19500 = ( ~n19352 & n19367 ) | ( ~n19352 & n19498 ) | ( n19367 & n19498 ) ;
  assign n19501 = n7037 & n15271 ;
  assign n19502 = ( n7036 & ~n15248 ) | ( n7036 & n19501 ) | ( ~n15248 & n19501 ) ;
  assign n19503 = n19501 | n19502 ;
  assign n19504 = n7035 & ~n18354 ;
  assign n19505 = ( n7052 & n15239 ) | ( n7052 & n19501 ) | ( n15239 & n19501 ) ;
  assign n19506 = n19503 | n19505 ;
  assign n19507 = n6901 & n15271 ;
  assign n19508 = n19504 | n19506 ;
  assign n19509 = ( n6906 & ~n15248 ) | ( n6906 & n19507 ) | ( ~n15248 & n19507 ) ;
  assign n19510 = n6901 & n15239 ;
  assign n19511 = n19507 | n19509 ;
  assign n19512 = ( n6907 & ~n15275 ) | ( n6907 & n19507 ) | ( ~n15275 & n19507 ) ;
  assign n19513 = n19511 | n19512 ;
  assign n19514 = ( n6906 & n15219 ) | ( n6906 & n19510 ) | ( n15219 & n19510 ) ;
  assign n19515 = n7037 & ~n15275 ;
  assign n19516 = n19510 | n19514 ;
  assign n19517 = n6918 & ~n18303 ;
  assign n19518 = ( n6907 & ~n15248 ) | ( n6907 & n19510 ) | ( ~n15248 & n19510 ) ;
  assign n19519 = n19516 | n19518 ;
  assign n19520 = ( n7036 & n15271 ) | ( n7036 & n19515 ) | ( n15271 & n19515 ) ;
  assign n19521 = ( n7052 & ~n15248 ) | ( n7052 & n19515 ) | ( ~n15248 & n19515 ) ;
  assign n19522 = n19517 | n19519 ;
  assign n19523 = n19515 | n19520 ;
  assign n19524 = n7035 & ~n18456 ;
  assign n19525 = n19521 | n19523 ;
  assign n19526 = n19524 | n19525 ;
  assign n19527 = n19526 ^ x26 ^ 1'b0 ;
  assign n19528 = n19508 ^ x26 ^ 1'b0 ;
  assign n19529 = ( n19360 & ~n19368 ) | ( n19360 & n19527 ) | ( ~n19368 & n19527 ) ;
  assign n19530 = n19528 ^ n19489 ^ n19349 ;
  assign n19531 = n19527 ^ n19368 ^ n19360 ;
  assign n19532 = n6918 & ~n18456 ;
  assign n19533 = n19513 & ~n19532 ;
  assign n19534 = n19533 ^ n19532 ^ x29 ;
  assign n19535 = ( n19349 & n19489 ) | ( n19349 & n19528 ) | ( n19489 & n19528 ) ;
  assign n19536 = ( n19351 & n19421 ) | ( n19351 & n19534 ) | ( n19421 & n19534 ) ;
  assign n19537 = n19534 ^ n19421 ^ n19351 ;
  assign n19538 = ( ~n19408 & n19479 ) | ( ~n19408 & n19536 ) | ( n19479 & n19536 ) ;
  assign n19539 = n19536 ^ n19479 ^ n19408 ;
  assign n19540 = n7037 & n15312 ;
  assign n19541 = ( n7036 & ~n15275 ) | ( n7036 & n19540 ) | ( ~n15275 & n19540 ) ;
  assign n19542 = n19540 | n19541 ;
  assign n19543 = ( n7052 & n15271 ) | ( n7052 & n19540 ) | ( n15271 & n19540 ) ;
  assign n19544 = n19542 | n19543 ;
  assign n19545 = n7035 & ~n18480 ;
  assign n19546 = n19544 | n19545 ;
  assign n19547 = n19546 ^ x26 ^ 1'b0 ;
  assign n19548 = n19522 ^ x29 ^ 1'b0 ;
  assign n19549 = n19548 ^ n19547 ^ n19366 ;
  assign n19550 = ( ~n19366 & n19547 ) | ( ~n19366 & n19548 ) | ( n19547 & n19548 ) ;
  assign n19551 = n6901 & n15312 ;
  assign n19552 = ( n6906 & ~n15275 ) | ( n6906 & n19551 ) | ( ~n15275 & n19551 ) ;
  assign n19553 = n19551 | n19552 ;
  assign n19554 = ( n6907 & n15308 ) | ( n6907 & n19551 ) | ( n15308 & n19551 ) ;
  assign n19555 = n19553 | n19554 ;
  assign n19556 = n6918 & n18525 ;
  assign n19557 = n19555 | n19556 ;
  assign n19558 = n19557 ^ x29 ^ 1'b0 ;
  assign n19559 = n19558 ^ n19538 ^ n19427 ;
  assign n19560 = ( ~n19427 & n19538 ) | ( ~n19427 & n19558 ) | ( n19538 & n19558 ) ;
  assign n19561 = n6901 & ~n15275 ;
  assign n19562 = ( n6906 & n15271 ) | ( n6906 & n19561 ) | ( n15271 & n19561 ) ;
  assign n19563 = n19561 | n19562 ;
  assign n19564 = ( n6907 & n15312 ) | ( n6907 & n19561 ) | ( n15312 & n19561 ) ;
  assign n19565 = n19563 | n19564 ;
  assign n19566 = n6918 & ~n18480 ;
  assign n19567 = n19565 | n19566 ;
  assign n19568 = n7188 & n15312 ;
  assign n19569 = ( n7190 & n15271 ) | ( n7190 & n19568 ) | ( n15271 & n19568 ) ;
  assign n19570 = n19568 | n19569 ;
  assign n19571 = ( n7192 & ~n15275 ) | ( n7192 & n19568 ) | ( ~n15275 & n19568 ) ;
  assign n19572 = n19570 | n19571 ;
  assign n19573 = n6918 & ~n18552 ;
  assign n19574 = n7196 & ~n18480 ;
  assign n19575 = n19572 | n19574 ;
  assign n19576 = n19575 ^ x23 ^ 1'b0 ;
  assign n19577 = n19576 ^ n19490 ^ n19377 ;
  assign n19578 = ( n19377 & n19490 ) | ( n19377 & n19576 ) | ( n19490 & n19576 ) ;
  assign n19579 = n6901 & n15319 ;
  assign n19580 = ( n6907 & ~n15320 ) | ( n6907 & n19579 ) | ( ~n15320 & n19579 ) ;
  assign n19581 = ( n6906 & n15308 ) | ( n6906 & n19579 ) | ( n15308 & n19579 ) ;
  assign n19582 = n19579 | n19581 ;
  assign n19583 = n19580 | n19582 ;
  assign n19584 = n19573 | n19583 ;
  assign n19585 = n19584 ^ x29 ^ 1'b0 ;
  assign n19586 = n19585 ^ n19458 ^ x26 ;
  assign n19587 = ( x26 & ~n19458 ) | ( x26 & n19585 ) | ( ~n19458 & n19585 ) ;
  assign n19588 = n19587 ^ n19480 ^ n19439 ;
  assign n19589 = n7188 & n15308 ;
  assign n19590 = ( n7190 & ~n15275 ) | ( n7190 & n19589 ) | ( ~n15275 & n19589 ) ;
  assign n19591 = n19589 | n19590 ;
  assign n19592 = ( n7192 & n15312 ) | ( n7192 & n19589 ) | ( n15312 & n19589 ) ;
  assign n19593 = n19591 | n19592 ;
  assign n19594 = n7196 & n18525 ;
  assign n19595 = n19593 | n19594 ;
  assign n19596 = n19595 ^ x23 ^ 1'b0 ;
  assign n19597 = n19596 ^ n19578 ^ n19530 ;
  assign n19598 = ( n19530 & n19578 ) | ( n19530 & n19596 ) | ( n19578 & n19596 ) ;
  assign n19599 = n7037 & n15308 ;
  assign n19600 = ( n7052 & ~n15275 ) | ( n7052 & n19599 ) | ( ~n15275 & n19599 ) ;
  assign n19601 = n7035 & n18525 ;
  assign n19602 = ( n7036 & n15312 ) | ( n7036 & n19599 ) | ( n15312 & n19599 ) ;
  assign n19603 = n19599 | n19602 ;
  assign n19604 = n7037 & n15319 ;
  assign n19605 = n19600 | n19603 ;
  assign n19606 = ( n7036 & n15308 ) | ( n7036 & n19604 ) | ( n15308 & n19604 ) ;
  assign n19607 = n19601 | n19605 ;
  assign n19608 = n19604 | n19606 ;
  assign n19609 = ( n7052 & n15312 ) | ( n7052 & n19604 ) | ( n15312 & n19604 ) ;
  assign n19610 = n19607 ^ x26 ^ 1'b0 ;
  assign n19611 = n7188 & n15319 ;
  assign n19612 = n7188 & ~n15320 ;
  assign n19613 = n19608 | n19609 ;
  assign n19614 = ( n7190 & n15308 ) | ( n7190 & n19612 ) | ( n15308 & n19612 ) ;
  assign n19615 = n19612 | n19614 ;
  assign n19616 = ( n7192 & n15319 ) | ( n7192 & n19612 ) | ( n15319 & n19612 ) ;
  assign n19617 = n19615 | n19616 ;
  assign n19618 = n7196 & ~n18552 ;
  assign n19619 = n19617 | n19618 ;
  assign n19620 = n19619 ^ x23 ^ 1'b0 ;
  assign n19621 = n19620 ^ n19549 ^ n19529 ;
  assign n19622 = ( n19529 & ~n19549 ) | ( n19529 & n19620 ) | ( ~n19549 & n19620 ) ;
  assign n19623 = n7035 & n18531 ;
  assign n19624 = n19613 | n19623 ;
  assign n19625 = n7196 & n18531 ;
  assign n19626 = n7190 & n15319 ;
  assign n19627 = n19624 ^ x26 ^ 1'b0 ;
  assign n19628 = n19627 ^ n19537 ^ n19500 ;
  assign n19629 = ( n19500 & n19537 ) | ( n19500 & n19627 ) | ( n19537 & n19627 ) ;
  assign n19630 = ( n7192 & ~n15320 ) | ( n7192 & n19626 ) | ( ~n15320 & n19626 ) ;
  assign n19631 = n19610 ^ n19550 ^ n19499 ;
  assign n19632 = ( n7196 & ~n18550 ) | ( n7196 & n19626 ) | ( ~n18550 & n19626 ) ;
  assign n19633 = n19626 | n19632 ;
  assign n19634 = n19630 | n19633 ;
  assign n19635 = ( n7192 & n15308 ) | ( n7192 & n19611 ) | ( n15308 & n19611 ) ;
  assign n19636 = n7190 & ~n15320 ;
  assign n19637 = n19636 ^ x23 ^ 1'b0 ;
  assign n19638 = ( n7190 & n15312 ) | ( n7190 & n19611 ) | ( n15312 & n19611 ) ;
  assign n19639 = n19611 | n19638 ;
  assign n19640 = n19635 | n19639 ;
  assign n19641 = n19625 | n19640 ;
  assign n19642 = n19634 ^ x23 ^ 1'b0 ;
  assign n19643 = n19642 ^ n19631 ^ n19622 ;
  assign n19644 = ( n19622 & ~n19631 ) | ( n19622 & n19642 ) | ( ~n19631 & n19642 ) ;
  assign n19645 = ( ~n19499 & n19550 ) | ( ~n19499 & n19610 ) | ( n19550 & n19610 ) ;
  assign n19646 = ( n19628 & n19637 ) | ( n19628 & n19645 ) | ( n19637 & n19645 ) ;
  assign n19647 = n19641 ^ x23 ^ 1'b0 ;
  assign n19648 = n19645 ^ n19637 ^ n19628 ;
  assign n19649 = n19647 ^ n19535 ^ n19531 ;
  assign n19650 = ( ~n19531 & n19535 ) | ( ~n19531 & n19647 ) | ( n19535 & n19647 ) ;
  assign n19651 = n7037 & ~n15320 ;
  assign n19652 = ( n7036 & n15319 ) | ( n7036 & n19651 ) | ( n15319 & n19651 ) ;
  assign n19653 = n19651 | n19652 ;
  assign n19654 = ( n7052 & n15308 ) | ( n7052 & n19651 ) | ( n15308 & n19651 ) ;
  assign n19655 = n19653 | n19654 ;
  assign n19656 = n7037 & n15322 ;
  assign n19657 = n7340 & ~n18552 ;
  assign n19658 = n7035 & ~n18552 ;
  assign n19659 = n19655 | n19658 ;
  assign n19660 = ( n7036 & ~n15320 ) | ( n7036 & n19656 ) | ( ~n15320 & n19656 ) ;
  assign n19661 = n19656 | n19660 ;
  assign n19662 = ( n7052 & n15319 ) | ( n7052 & n19656 ) | ( n15319 & n19656 ) ;
  assign n19663 = n7340 & ~n18550 ;
  assign n19664 = n7035 & ~n18550 ;
  assign n19665 = n7339 & n15319 ;
  assign n19666 = n19661 | n19662 ;
  assign n19667 = ( n7337 & ~n15320 ) | ( n7337 & n19665 ) | ( ~n15320 & n19665 ) ;
  assign n19668 = n7036 & n15322 ;
  assign n19669 = n19665 | n19667 ;
  assign n19670 = n19664 | n19666 ;
  assign n19671 = n19670 ^ x26 ^ 1'b0 ;
  assign n19672 = n7339 & ~n15320 ;
  assign n19673 = ( n7338 & n15319 ) | ( n7338 & n19672 ) | ( n15319 & n19672 ) ;
  assign n19674 = ( n7337 & n15322 ) | ( n7337 & n19672 ) | ( n15322 & n19672 ) ;
  assign n19675 = n19672 | n19674 ;
  assign n19676 = n19673 | n19675 ;
  assign n19677 = n19567 ^ x29 ^ 1'b0 ;
  assign n19678 = n19663 | n19676 ;
  assign n19679 = n19659 ^ x26 ^ 1'b0 ;
  assign n19680 = n19678 ^ x20 ^ 1'b0 ;
  assign n19681 = ( ~n19539 & n19677 ) | ( ~n19539 & n19679 ) | ( n19677 & n19679 ) ;
  assign n19682 = n7339 & n15322 ;
  assign n19683 = ( n7052 & ~n15320 ) | ( n7052 & n19668 ) | ( ~n15320 & n19668 ) ;
  assign n19684 = ( n7338 & n15308 ) | ( n7338 & n19665 ) | ( n15308 & n19665 ) ;
  assign n19685 = n19669 | n19684 ;
  assign n19686 = ( n7338 & ~n15320 ) | ( n7338 & n19682 ) | ( ~n15320 & n19682 ) ;
  assign n19687 = n19679 ^ n19677 ^ n19539 ;
  assign n19688 = n19657 | n19685 ;
  assign n19689 = n19688 ^ x20 ^ 1'b0 ;
  assign n19690 = n19689 ^ n19577 ^ n19395 ;
  assign n19691 = n19682 | n19686 ;
  assign n19692 = n19691 ^ x20 ^ 1'b0 ;
  assign n19693 = n19668 | n19683 ;
  assign n19694 = ( n19598 & ~n19649 ) | ( n19598 & n19692 ) | ( ~n19649 & n19692 ) ;
  assign n19695 = n19692 ^ n19649 ^ n19598 ;
  assign n19696 = ( n19395 & n19577 ) | ( n19395 & n19689 ) | ( n19577 & n19689 ) ;
  assign n19697 = n19696 ^ n19680 ^ n19597 ;
  assign n19698 = ( n19597 & n19680 ) | ( n19597 & n19696 ) | ( n19680 & n19696 ) ;
  assign n19699 = n19681 ^ n19671 ^ n19559 ;
  assign n19700 = ( ~n19559 & n19671 ) | ( ~n19559 & n19681 ) | ( n19671 & n19681 ) ;
  assign n19701 = n19690 ^ n19406 ^ x17 ;
  assign n19702 = ( x17 & n19406 ) | ( x17 & n19690 ) | ( n19406 & n19690 ) ;
  assign n19703 = ( n19422 & n19424 ) | ( n19422 & n19701 ) | ( n19424 & n19701 ) ;
  assign n19704 = n19701 ^ n19422 ^ 1'b0 ;
  assign n19705 = n19650 ^ n19621 ^ x20 ;
  assign n19706 = n19704 ^ n19424 ^ 1'b0 ;
  assign n19707 = n19702 ^ n19697 ^ 1'b0 ;
  assign n19708 = ( n19697 & n19702 ) | ( n19697 & n19703 ) | ( n19702 & n19703 ) ;
  assign n19709 = ( ~n19695 & n19698 ) | ( ~n19695 & n19708 ) | ( n19698 & n19708 ) ;
  assign n19710 = n19707 ^ n19703 ^ 1'b0 ;
  assign n19711 = n19705 ^ n19694 ^ 1'b0 ;
  assign n19712 = ( x20 & ~n19621 ) | ( x20 & n19650 ) | ( ~n19621 & n19650 ) ;
  assign n19713 = ( n19694 & ~n19705 ) | ( n19694 & n19709 ) | ( ~n19705 & n19709 ) ;
  assign n19714 = ( x23 & n19629 ) | ( x23 & ~n19687 ) | ( n19629 & ~n19687 ) ;
  assign n19715 = ( ~n19643 & n19712 ) | ( ~n19643 & n19713 ) | ( n19712 & n19713 ) ;
  assign n19716 = n19698 ^ n19695 ^ 1'b0 ;
  assign n19717 = n19687 ^ n19629 ^ x23 ;
  assign n19718 = ~n18592 & n19320 ;
  assign n19719 = ( n19644 & n19648 ) | ( n19644 & n19715 ) | ( n19648 & n19715 ) ;
  assign n19720 = n19693 ^ x26 ^ 1'b0 ;
  assign n19721 = n19648 ^ n19644 ^ 1'b0 ;
  assign n19722 = n19320 ^ n18592 ^ 1'b0 ;
  assign n19723 = ( n19646 & ~n19717 ) | ( n19646 & n19719 ) | ( ~n19717 & n19719 ) ;
  assign n19724 = ( ~n19699 & n19714 ) | ( ~n19699 & n19723 ) | ( n19714 & n19723 ) ;
  assign n19725 = n19712 ^ n19643 ^ 1'b0 ;
  assign n19726 = n19717 ^ n19646 ^ 1'b0 ;
  assign n19727 = n19726 ^ n19719 ^ 1'b0 ;
  assign n19728 = n19725 ^ n19713 ^ 1'b0 ;
  assign n19729 = ( n19449 & n19560 ) | ( n19449 & n19720 ) | ( n19560 & n19720 ) ;
  assign n19730 = n19720 ^ n19560 ^ n19449 ;
  assign n19731 = n19730 ^ n19700 ^ 1'b0 ;
  assign n19732 = ( n19700 & n19724 ) | ( n19700 & n19730 ) | ( n19724 & n19730 ) ;
  assign n19733 = ( ~n19586 & n19729 ) | ( ~n19586 & n19732 ) | ( n19729 & n19732 ) ;
  assign n19734 = n19718 ^ n18597 ^ 1'b0 ;
  assign n19735 = n19721 ^ n19715 ^ 1'b0 ;
  assign n19736 = n19716 ^ n19708 ^ 1'b0 ;
  assign n19737 = n19729 ^ n19586 ^ 1'b0 ;
  assign n19738 = ~n18597 & n19718 ;
  assign n19739 = n19714 ^ n19699 ^ 1'b0 ;
  assign n19740 = n19739 ^ n19723 ^ 1'b0 ;
  assign n19741 = n19737 ^ n19732 ^ 1'b0 ;
  assign n19742 = n19711 ^ n19709 ^ 1'b0 ;
  assign n19743 = n19731 ^ n19724 ^ 1'b0 ;
  assign n19744 = n19738 ^ n18653 ^ 1'b0 ;
  assign n19745 = ~n18653 & n19738 ;
  assign n19746 = n19745 ^ n18709 ^ 1'b0 ;
  assign n19747 = n18709 & n19745 ;
  assign n19748 = n19747 ^ n18784 ^ 1'b0 ;
  assign n19749 = n18784 & n19747 ;
  assign n19750 = n19749 ^ n18828 ^ 1'b0 ;
  assign n19751 = n18828 & n19749 ;
  assign n19752 = n19751 ^ n18857 ^ 1'b0 ;
  assign n19753 = n18857 & n19751 ;
  assign n19754 = n19753 ^ n18926 ^ 1'b0 ;
  assign n19755 = ~n18926 & n19753 ;
  assign n19756 = n19755 ^ n18964 ^ 1'b0 ;
  assign n19757 = ~n18964 & n19755 ;
  assign n19758 = n19757 ^ n19007 ^ 1'b0 ;
  assign n19759 = ~n19007 & n19757 ;
  assign n19760 = n19759 ^ n19062 ^ 1'b0 ;
  assign n19761 = n19062 & n19759 ;
  assign n19762 = n19761 ^ n19129 ^ 1'b0 ;
  assign n19763 = ~n19129 & n19761 ;
  assign n19764 = n19763 ^ n19185 ^ 1'b0 ;
  assign n19765 = n19185 & n19763 ;
  assign n19766 = n19765 ^ n19250 ^ 1'b0 ;
  assign n19767 = ~n19250 & n19765 ;
  assign n19768 = n19767 ^ n19301 ^ 1'b0 ;
  assign n19769 = ~n19301 & n19767 ;
  assign n19770 = n19769 ^ n19426 ^ 1'b0 ;
  assign n19771 = ~n19426 & n19769 ;
  assign n19772 = n19771 ^ n19706 ^ 1'b0 ;
  assign n19773 = n19706 & n19771 ;
  assign n19774 = n19773 ^ n19710 ^ 1'b0 ;
  assign n19775 = n19710 & n19773 ;
  assign n19776 = n19775 ^ n19736 ^ 1'b0 ;
  assign n19777 = ~n19736 & n19775 ;
  assign n19778 = n19777 ^ n19742 ^ 1'b0 ;
  assign n19779 = ~n19742 & n19777 ;
  assign n19780 = n19779 ^ n19728 ^ 1'b0 ;
  assign n19781 = ~n19728 & n19779 ;
  assign n19782 = n19781 ^ n19735 ^ 1'b0 ;
  assign n19783 = n19735 & n19781 ;
  assign n19784 = n19783 ^ n19727 ^ 1'b0 ;
  assign n19785 = ~n19727 & n19783 ;
  assign n19786 = n19785 ^ n19740 ^ 1'b0 ;
  assign n19787 = ~n19740 & n19785 ;
  assign n19788 = n19787 ^ n19743 ^ 1'b0 ;
  assign n19789 = n19743 & n19787 ;
  assign n19790 = n19789 ^ n19741 ^ 1'b0 ;
  assign n19791 = ~n19741 & n19789 ;
  assign n19792 = n19791 ^ n19733 ^ n19588 ;
  assign y0 = n19302 ;
  assign y1 = n19311 ;
  assign y2 = ~n19317 ;
  assign y3 = ~n19318 ;
  assign y4 = ~n19321 ;
  assign y5 = ~n19722 ;
  assign y6 = ~n19734 ;
  assign y7 = ~n19744 ;
  assign y8 = n19746 ;
  assign y9 = n19748 ;
  assign y10 = n19750 ;
  assign y11 = n19752 ;
  assign y12 = ~n19754 ;
  assign y13 = ~n19756 ;
  assign y14 = ~n19758 ;
  assign y15 = n19760 ;
  assign y16 = ~n19762 ;
  assign y17 = n19764 ;
  assign y18 = ~n19766 ;
  assign y19 = ~n19768 ;
  assign y20 = ~n19770 ;
  assign y21 = n19772 ;
  assign y22 = n19774 ;
  assign y23 = ~n19776 ;
  assign y24 = ~n19778 ;
  assign y25 = ~n19780 ;
  assign y26 = n19782 ;
  assign y27 = ~n19784 ;
  assign y28 = ~n19786 ;
  assign y29 = n19788 ;
  assign y30 = ~n19790 ;
  assign y31 = n19792 ;
endmodule
