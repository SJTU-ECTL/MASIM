module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , y0 , y1 , y2 , y3 , y4 , y5 , y6 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 ;
  wire n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 ;
  assign n12 = x5 & ~x6 ;
  assign n13 = ~x4 & x5 ;
  assign n14 = ~x3 & n12 ;
  assign n15 = ( ~x3 & x7 ) | ( ~x3 & n14 ) | ( x7 & n14 ) ;
  assign n16 = ( x1 & ~x3 ) | ( x1 & n13 ) | ( ~x3 & n13 ) ;
  assign n17 = x4 & ~x6 ;
  assign n18 = ( x0 & x3 ) | ( x0 & n17 ) | ( x3 & n17 ) ;
  assign n19 = ( x1 & x3 ) | ( x1 & n18 ) | ( x3 & n18 ) ;
  assign n20 = n16 & n19 ;
  assign n21 = x3 & ~x4 ;
  assign n22 = ~x1 & n12 ;
  assign n23 = ( x2 & x6 ) | ( x2 & n22 ) | ( x6 & n22 ) ;
  assign n24 = x6 & ~x7 ;
  assign n25 = ( x4 & ~n15 ) | ( x4 & n24 ) | ( ~n15 & n24 ) ;
  assign n26 = ~n15 & n25 ;
  assign n27 = ~x2 & n24 ;
  assign n28 = x5 & x6 ;
  assign n29 = x0 & x1 ;
  assign n30 = x6 ^ x4 ^ 1'b0 ;
  assign n31 = x5 & ~n22 ;
  assign n32 = ( n22 & n23 ) | ( n22 & ~n31 ) | ( n23 & ~n31 ) ;
  assign n33 = n32 ^ n21 ^ x3 ;
  assign n34 = ( n28 & n32 ) | ( n28 & ~n33 ) | ( n32 & ~n33 ) ;
  assign n35 = x7 & n28 ;
  assign n36 = x3 & ~n29 ;
  assign n37 = ( x6 & n30 ) | ( x6 & ~n36 ) | ( n30 & ~n36 ) ;
  assign n38 = x7 & ~n28 ;
  assign n39 = x5 & ~n37 ;
  assign n40 = ( ~n20 & n37 ) | ( ~n20 & n39 ) | ( n37 & n39 ) ;
  assign n41 = x2 & ~n40 ;
  assign n42 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n43 = ( x2 & x3 ) | ( x2 & ~x4 ) | ( x3 & ~x4 ) ;
  assign n44 = ( x3 & x6 ) | ( x3 & n43 ) | ( x6 & n43 ) ;
  assign n45 = n42 & ~n44 ;
  assign n46 = n41 | n45 ;
  assign n47 = x8 & n35 ;
  assign n48 = ( x5 & x7 ) | ( x5 & ~n47 ) | ( x7 & ~n47 ) ;
  assign n49 = ~x7 & n46 ;
  assign n50 = n34 | n49 ;
  assign n51 = ( x3 & n29 ) | ( x3 & n47 ) | ( n29 & n47 ) ;
  assign n52 = ( n47 & ~n48 ) | ( n47 & n51 ) | ( ~n48 & n51 ) ;
  assign n53 = x8 & ~n47 ;
  assign n54 = ( n47 & n52 ) | ( n47 & ~n53 ) | ( n52 & ~n53 ) ;
  assign n55 = x2 & n54 ;
  assign n56 = x1 & x2 ;
  assign n57 = ( x3 & n14 ) | ( x3 & n47 ) | ( n14 & n47 ) ;
  assign n58 = n55 | n57 ;
  assign n59 = n12 & ~n56 ;
  assign n60 = ( ~x9 & n38 ) | ( ~x9 & n59 ) | ( n38 & n59 ) ;
  assign n61 = ( ~x9 & n26 ) | ( ~x9 & n60 ) | ( n26 & n60 ) ;
  assign n62 = ~n60 & n61 ;
  assign n63 = x4 & n58 ;
  assign n64 = x1 & ~x2 ;
  assign n65 = x5 & ~x7 ;
  assign n66 = ( x3 & x4 ) | ( x3 & x7 ) | ( x4 & x7 ) ;
  assign n67 = n64 & ~n65 ;
  assign n68 = ( x3 & ~n64 ) | ( x3 & n67 ) | ( ~n64 & n67 ) ;
  assign n69 = ( n21 & n66 ) | ( n21 & ~n68 ) | ( n66 & ~n68 ) ;
  assign n70 = x4 & x6 ;
  assign n71 = ~x6 & x7 ;
  assign n72 = ( n65 & n70 ) | ( n65 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ( ~x6 & n29 ) | ( ~x6 & n72 ) | ( n29 & n72 ) ;
  assign n74 = ( ~n12 & n72 ) | ( ~n12 & n73 ) | ( n72 & n73 ) ;
  assign n75 = x3 & n71 ;
  assign n76 = n27 | n75 ;
  assign n77 = ( x8 & n71 ) | ( x8 & n72 ) | ( n71 & n72 ) ;
  assign n78 = x2 & x3 ;
  assign n79 = n70 & n78 ;
  assign n80 = n62 & n78 ;
  assign n81 = n74 & n80 ;
  assign n82 = x8 | x9 ;
  assign n83 = n50 & ~n82 ;
  assign n84 = ( x8 & n62 ) | ( x8 & ~n81 ) | ( n62 & ~n81 ) ;
  assign n85 = x6 & ~x9 ;
  assign n86 = ( n17 & n79 ) | ( n17 & n85 ) | ( n79 & n85 ) ;
  assign n87 = ~x4 & n85 ;
  assign n88 = ( ~x3 & n22 ) | ( ~x3 & n87 ) | ( n22 & n87 ) ;
  assign n89 = ( ~x10 & n86 ) | ( ~x10 & n88 ) | ( n86 & n88 ) ;
  assign n90 = x4 & x5 ;
  assign n91 = ( n13 & n79 ) | ( n13 & n90 ) | ( n79 & n90 ) ;
  assign n92 = n14 | n87 ;
  assign n93 = x6 & x7 ;
  assign n94 = n93 ^ n90 ^ 1'b0 ;
  assign n95 = ( n76 & n93 ) | ( n76 & n94 ) | ( n93 & n94 ) ;
  assign n96 = ( ~x9 & n83 ) | ( ~x9 & n95 ) | ( n83 & n95 ) ;
  assign n97 = n77 | n96 ;
  assign n98 = n35 ^ x9 ^ 1'b0 ;
  assign n99 = x5 & x7 ;
  assign n100 = x10 | n84 ;
  assign n101 = n69 ^ x8 ^ 1'b0 ;
  assign n102 = ( n13 & n69 ) | ( n13 & n101 ) | ( n69 & n101 ) ;
  assign n103 = x2 | x7 ;
  assign n104 = n70 & n99 ;
  assign n105 = x3 ^ x2 ^ 1'b0 ;
  assign n106 = n92 & ~n103 ;
  assign n107 = x10 | n89 ;
  assign n108 = ( ~x7 & n106 ) | ( ~x7 & n107 ) | ( n106 & n107 ) ;
  assign n109 = ( x2 & x8 ) | ( x2 & n105 ) | ( x8 & n105 ) ;
  assign n110 = x8 & ~n99 ;
  assign n111 = n104 & n109 ;
  assign n112 = ( ~n35 & n98 ) | ( ~n35 & n111 ) | ( n98 & n111 ) ;
  assign n113 = ( x10 & n100 ) | ( x10 & ~n112 ) | ( n100 & ~n112 ) ;
  assign n114 = ( x5 & x9 ) | ( x5 & ~n93 ) | ( x9 & ~n93 ) ;
  assign n115 = x9 & x10 ;
  assign n116 = x8 | n114 ;
  assign n117 = x8 & ~x10 ;
  assign n118 = ( x9 & n110 ) | ( x9 & n115 ) | ( n110 & n115 ) ;
  assign n119 = ( n93 & ~n116 ) | ( n93 & n117 ) | ( ~n116 & n117 ) ;
  assign n120 = ( n93 & n118 ) | ( n93 & ~n119 ) | ( n118 & ~n119 ) ;
  assign n121 = ~x1 & x4 ;
  assign n122 = x8 & n115 ;
  assign n123 = x10 & n97 ;
  assign n124 = ( n97 & n120 ) | ( n97 & ~n123 ) | ( n120 & ~n123 ) ;
  assign n125 = ( x4 & ~x7 ) | ( x4 & n64 ) | ( ~x7 & n64 ) ;
  assign n126 = n91 ^ n12 ^ x6 ;
  assign n127 = x3 | x8 ;
  assign n128 = ( x4 & ~n64 ) | ( x4 & n127 ) | ( ~n64 & n127 ) ;
  assign n129 = ( x10 & ~n82 ) | ( x10 & n105 ) | ( ~n82 & n105 ) ;
  assign n130 = n125 & ~n128 ;
  assign n131 = x7 & ~n122 ;
  assign n132 = ( ~x7 & x10 ) | ( ~x7 & n129 ) | ( x10 & n129 ) ;
  assign n133 = ( n122 & ~n131 ) | ( n122 & n132 ) | ( ~n131 & n132 ) ;
  assign n134 = ( x2 & x9 ) | ( x2 & ~n56 ) | ( x9 & ~n56 ) ;
  assign n135 = x7 | x8 ;
  assign n136 = ( x9 & n134 ) | ( x9 & ~n135 ) | ( n134 & ~n135 ) ;
  assign n137 = n130 | n136 ;
  assign n138 = x9 | x10 ;
  assign n139 = ( n91 & ~n135 ) | ( n91 & n138 ) | ( ~n135 & n138 ) ;
  assign n140 = ~x6 & n137 ;
  assign n141 = n135 | n139 ;
  assign n142 = n121 ^ x4 ^ x0 ;
  assign n143 = n126 & ~n135 ;
  assign n144 = ( n63 & ~n138 ) | ( n63 & n143 ) | ( ~n138 & n143 ) ;
  assign n145 = x6 & x9 ;
  assign n146 = n145 ^ x5 ^ 1'b0 ;
  assign n147 = ( n140 & n145 ) | ( n140 & n146 ) | ( n145 & n146 ) ;
  assign n148 = x4 | x8 ;
  assign n149 = ( x4 & n142 ) | ( x4 & ~n148 ) | ( n142 & ~n148 ) ;
  assign n150 = x4 & x8 ;
  assign n151 = ( ~x6 & x7 ) | ( ~x6 & n149 ) | ( x7 & n149 ) ;
  assign n152 = ~x7 & n151 ;
  assign n153 = n150 | n152 ;
  assign n154 = ~x5 & n153 ;
  assign n155 = x6 & n133 ;
  assign n156 = n102 | n154 ;
  assign n157 = ~x9 & n156 ;
  assign n158 = ~x6 & x10 ;
  assign n159 = n147 | n157 ;
  assign n160 = ~x7 & n158 ;
  assign n161 = ( n155 & n158 ) | ( n155 & ~n160 ) | ( n158 & ~n160 ) ;
  assign n162 = x10 & n159 ;
  assign n163 = ( n159 & n161 ) | ( n159 & ~n162 ) | ( n161 & ~n162 ) ;
  assign n164 = n108 | n158 ;
  assign n165 = x4 | x9 ;
  assign n166 = n103 & ~n165 ;
  assign n167 = ( x1 & n103 ) | ( x1 & ~n166 ) | ( n103 & ~n166 ) ;
  assign n168 = ~x7 & n167 ;
  assign n169 = ( n82 & n127 ) | ( n82 & n165 ) | ( n127 & n165 ) ;
  assign n170 = ( ~x0 & x4 ) | ( ~x0 & n56 ) | ( x4 & n56 ) ;
  assign n171 = n168 & n170 ;
  assign n172 = ( x0 & ~x2 ) | ( x0 & x4 ) | ( ~x2 & x4 ) ;
  assign n173 = n171 & n172 ;
  assign n174 = n138 | n144 ;
  assign n175 = x8 & ~x9 ;
  assign n176 = n167 & ~n175 ;
  assign n177 = n173 & ~n175 ;
  assign n178 = ( x6 & n176 ) | ( x6 & ~n177 ) | ( n176 & ~n177 ) ;
  assign n179 = x9 ^ x7 ^ 1'b0 ;
  assign n180 = ( x9 & ~n169 ) | ( x9 & n179 ) | ( ~n169 & n179 ) ;
  assign n181 = n178 & ~n180 ;
  assign n182 = ( x2 & x5 ) | ( x2 & ~n150 ) | ( x5 & ~n150 ) ;
  assign n183 = n93 & ~n182 ;
  assign n184 = x10 & n175 ;
  assign n185 = x5 & ~n183 ;
  assign n186 = n93 & n184 ;
  assign n187 = x8 & n164 ;
  assign n188 = ( n164 & n186 ) | ( n164 & ~n187 ) | ( n186 & ~n187 ) ;
  assign n189 = ( ~x3 & x4 ) | ( ~x3 & n82 ) | ( x4 & n82 ) ;
  assign n190 = ( x4 & x7 ) | ( x4 & n56 ) | ( x7 & n56 ) ;
  assign n191 = ( n56 & ~n189 ) | ( n56 & n190 ) | ( ~n189 & n190 ) ;
  assign n192 = x6 | x7 ;
  assign n193 = ( ~x5 & n148 ) | ( ~x5 & n192 ) | ( n148 & n192 ) ;
  assign n194 = ( x3 & x4 ) | ( x3 & ~n192 ) | ( x4 & ~n192 ) ;
  assign n195 = ( n189 & ~n191 ) | ( n189 & n194 ) | ( ~n191 & n194 ) ;
  assign n196 = x5 & ~n185 ;
  assign n197 = ( n185 & n193 ) | ( n185 & ~n196 ) | ( n193 & ~n196 ) ;
  assign n198 = ( x7 & n150 ) | ( x7 & ~n179 ) | ( n150 & ~n179 ) ;
  assign n199 = n198 ^ n82 ^ 1'b0 ;
  assign n200 = ~x6 & n199 ;
  assign n201 = ~x6 & n198 ;
  assign n202 = ( ~x3 & n138 ) | ( ~x3 & n197 ) | ( n138 & n197 ) ;
  assign n203 = n194 & ~n195 ;
  assign n204 = ( x5 & n181 ) | ( x5 & ~n200 ) | ( n181 & ~n200 ) ;
  assign n205 = ( n198 & ~n201 ) | ( n198 & n203 ) | ( ~n201 & n203 ) ;
  assign n206 = x3 | n202 ;
  assign n207 = ( x5 & n200 ) | ( x5 & n205 ) | ( n200 & n205 ) ;
  assign n208 = n204 & n207 ;
  assign n209 = ( x10 & n204 ) | ( x10 & ~n208 ) | ( n204 & ~n208 ) ;
  assign n210 = ~n188 & n209 ;
  assign y0 = n163 ;
  assign y1 = n210 ;
  assign y2 = n124 ;
  assign y3 = n206 ;
  assign y4 = n113 ;
  assign y5 = n174 ;
  assign y6 = n141 ;
endmodule
