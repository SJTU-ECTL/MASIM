module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 ;
  assign n129 = x58 ^ x57 ^ 1'b0 ;
  assign n130 = x57 ^ x56 ^ 1'b0 ;
  assign n131 = x59 ^ x58 ^ 1'b0 ;
  assign n132 = ( n129 & ~n130 ) | ( n129 & n131 ) | ( ~n130 & n131 ) ;
  assign n133 = ~n129 & n132 ;
  assign n134 = n129 & ~n130 ;
  assign n135 = x66 & ~n134 ;
  assign n136 = x65 & n133 ;
  assign n137 = x64 & x65 ;
  assign n138 = x66 & n133 ;
  assign n139 = n137 ^ x66 ^ x65 ;
  assign n140 = n130 & n131 ;
  assign n141 = x69 & ~n134 ;
  assign n142 = n130 & ~n131 ;
  assign n143 = x67 & n133 ;
  assign n144 = x68 & n133 ;
  assign n145 = ( x70 & n142 ) | ( x70 & n144 ) | ( n142 & n144 ) ;
  assign n146 = n144 | n145 ;
  assign n147 = ( x69 & ~n141 ) | ( x69 & n146 ) | ( ~n141 & n146 ) ;
  assign n148 = ( x69 & n142 ) | ( x69 & n143 ) | ( n142 & n143 ) ;
  assign n149 = ( x67 & n136 ) | ( x67 & n142 ) | ( n136 & n142 ) ;
  assign n150 = n139 & n140 ;
  assign n151 = n143 | n148 ;
  assign n152 = x65 & ~n134 ;
  assign n153 = x64 & n133 ;
  assign n154 = ( x68 & n138 ) | ( x68 & n142 ) | ( n138 & n142 ) ;
  assign n155 = n136 | n149 ;
  assign n156 = x68 & ~n134 ;
  assign n157 = ( x68 & n151 ) | ( x68 & ~n156 ) | ( n151 & ~n156 ) ;
  assign n158 = ( x66 & n142 ) | ( x66 & n153 ) | ( n142 & n153 ) ;
  assign n159 = n153 | n158 ;
  assign n160 = ( x65 & x66 ) | ( x65 & n137 ) | ( x66 & n137 ) ;
  assign n161 = n160 ^ x67 ^ x66 ;
  assign n162 = ( x66 & x67 ) | ( x66 & n160 ) | ( x67 & n160 ) ;
  assign n163 = ( x65 & ~n152 ) | ( x65 & n159 ) | ( ~n152 & n159 ) ;
  assign n164 = ( x67 & x68 ) | ( x67 & n162 ) | ( x68 & n162 ) ;
  assign n165 = n150 | n163 ;
  assign n166 = ( x68 & x69 ) | ( x68 & n164 ) | ( x69 & n164 ) ;
  assign n167 = ( x66 & ~n135 ) | ( x66 & n155 ) | ( ~n135 & n155 ) ;
  assign n168 = n166 ^ x70 ^ x69 ;
  assign n169 = n138 | n154 ;
  assign n170 = n140 & n168 ;
  assign n171 = n165 ^ x59 ^ 1'b0 ;
  assign n172 = n164 ^ x69 ^ x68 ;
  assign n173 = n147 | n170 ;
  assign n174 = n173 ^ x59 ^ 1'b0 ;
  assign n175 = n162 ^ x68 ^ x67 ;
  assign n176 = x67 & ~n134 ;
  assign n177 = ( x69 & x70 ) | ( x69 & n166 ) | ( x70 & n166 ) ;
  assign n178 = ( x67 & n169 ) | ( x67 & ~n176 ) | ( n169 & ~n176 ) ;
  assign n179 = x64 & n130 ;
  assign n180 = n140 & n172 ;
  assign n181 = n157 | n180 ;
  assign n182 = n140 & n175 ;
  assign n183 = n178 | n182 ;
  assign n184 = n183 ^ x59 ^ 1'b0 ;
  assign n185 = n140 & n161 ;
  assign n186 = n167 | n185 ;
  assign n187 = n186 ^ x59 ^ 1'b0 ;
  assign n188 = n181 ^ x59 ^ 1'b0 ;
  assign n189 = x60 ^ x59 ^ 1'b0 ;
  assign n190 = x65 ^ x64 ^ 1'b0 ;
  assign n191 = x61 ^ x60 ^ 1'b0 ;
  assign n192 = ~n189 & n191 ;
  assign n193 = x62 ^ x61 ^ 1'b0 ;
  assign n194 = n189 & ~n193 ;
  assign n195 = x64 & n192 ;
  assign n196 = ~x65 & n194 ;
  assign n197 = n189 & n193 ;
  assign n198 = ( n190 & n195 ) | ( n190 & n197 ) | ( n195 & n197 ) ;
  assign n199 = ( ~n189 & n191 ) | ( ~n189 & n193 ) | ( n191 & n193 ) ;
  assign n200 = x64 & n134 ;
  assign n201 = ( n140 & n190 ) | ( n140 & n200 ) | ( n190 & n200 ) ;
  assign n202 = ( n194 & n195 ) | ( n194 & ~n196 ) | ( n195 & ~n196 ) ;
  assign n203 = n198 | n202 ;
  assign n204 = ~x65 & n142 ;
  assign n205 = ( n142 & n200 ) | ( n142 & ~n204 ) | ( n200 & ~n204 ) ;
  assign n206 = x64 & n189 ;
  assign n207 = x59 & ~n179 ;
  assign n208 = ~n191 & n199 ;
  assign n209 = n201 | n205 ;
  assign n210 = x65 & n208 ;
  assign n211 = ( x67 & n194 ) | ( x67 & n210 ) | ( n194 & n210 ) ;
  assign n212 = n210 | n211 ;
  assign n213 = x66 & ~n192 ;
  assign n214 = ( x66 & n212 ) | ( x66 & ~n213 ) | ( n212 & ~n213 ) ;
  assign n215 = n161 & n197 ;
  assign n216 = n214 | n215 ;
  assign n217 = n203 ^ x62 ^ 1'b0 ;
  assign n218 = n209 ^ x59 ^ 1'b0 ;
  assign n219 = x62 & ~n206 ;
  assign n220 = n207 & n218 ;
  assign n221 = n218 ^ n207 ^ 1'b0 ;
  assign n222 = n171 & n220 ;
  assign n223 = n220 ^ n171 ^ 1'b0 ;
  assign n224 = n222 ^ n206 ^ n187 ;
  assign n225 = ( n187 & n206 ) | ( n187 & n222 ) | ( n206 & n222 ) ;
  assign n226 = n217 & n219 ;
  assign n227 = n219 ^ n217 ^ 1'b0 ;
  assign n228 = x64 & n208 ;
  assign n229 = n227 ^ n225 ^ n184 ;
  assign n230 = ( n184 & n225 ) | ( n184 & n227 ) | ( n225 & n227 ) ;
  assign n231 = n139 & n197 ;
  assign n232 = ( x66 & n194 ) | ( x66 & n228 ) | ( n194 & n228 ) ;
  assign n233 = n228 | n232 ;
  assign n234 = x65 & ~n192 ;
  assign n235 = ( x65 & n233 ) | ( x65 & ~n234 ) | ( n233 & ~n234 ) ;
  assign n236 = n231 | n235 ;
  assign n237 = n216 ^ x62 ^ 1'b0 ;
  assign n238 = n236 ^ x62 ^ 1'b0 ;
  assign n239 = n238 ^ n226 ^ 1'b0 ;
  assign n240 = n239 ^ n230 ^ n188 ;
  assign n241 = ( n188 & n230 ) | ( n188 & n239 ) | ( n230 & n239 ) ;
  assign n242 = x63 ^ x62 ^ 1'b0 ;
  assign n243 = x64 & n242 ;
  assign n244 = n226 & n238 ;
  assign n245 = ( n237 & n243 ) | ( n237 & n244 ) | ( n243 & n244 ) ;
  assign n246 = n244 ^ n243 ^ n237 ;
  assign n247 = x66 & n208 ;
  assign n248 = ( x68 & n194 ) | ( x68 & n247 ) | ( n194 & n247 ) ;
  assign n249 = n247 | n248 ;
  assign n250 = x67 & ~n192 ;
  assign n251 = ( x67 & n249 ) | ( x67 & ~n250 ) | ( n249 & ~n250 ) ;
  assign n252 = n175 & n197 ;
  assign n253 = n251 | n252 ;
  assign n254 = n246 ^ n241 ^ n174 ;
  assign n255 = n253 ^ x62 ^ 1'b0 ;
  assign n256 = ( n174 & n241 ) | ( n174 & n246 ) | ( n241 & n246 ) ;
  assign n257 = x56 ^ x55 ^ 1'b0 ;
  assign n258 = x54 ^ x53 ^ 1'b0 ;
  assign n259 = x55 ^ x54 ^ 1'b0 ;
  assign n260 = ~n258 & n259 ;
  assign n261 = x64 & n260 ;
  assign n262 = ( n257 & ~n258 ) | ( n257 & n259 ) | ( ~n258 & n259 ) ;
  assign n263 = ~n259 & n262 ;
  assign n264 = ~n257 & n258 ;
  assign n265 = ~x65 & n264 ;
  assign n266 = x64 & n263 ;
  assign n267 = ( x66 & n264 ) | ( x66 & n266 ) | ( n264 & n266 ) ;
  assign n268 = n266 | n267 ;
  assign n269 = ( n261 & n264 ) | ( n261 & ~n265 ) | ( n264 & ~n265 ) ;
  assign n270 = x65 & ~n260 ;
  assign n271 = ( x65 & n268 ) | ( x65 & ~n270 ) | ( n268 & ~n270 ) ;
  assign n272 = n257 & n258 ;
  assign n273 = x64 & n258 ;
  assign n274 = ( n190 & n261 ) | ( n190 & n272 ) | ( n261 & n272 ) ;
  assign n275 = n139 & n272 ;
  assign n276 = n271 | n275 ;
  assign n277 = n269 | n274 ;
  assign n278 = x56 & ~n273 ;
  assign n279 = n277 ^ x56 ^ 1'b0 ;
  assign n280 = x65 & n263 ;
  assign n281 = ( x67 & n264 ) | ( x67 & n280 ) | ( n264 & n280 ) ;
  assign n282 = n280 | n281 ;
  assign n283 = n278 & n279 ;
  assign n284 = n276 ^ x56 ^ 1'b0 ;
  assign n285 = n279 ^ n278 ^ 1'b0 ;
  assign n286 = n283 & n284 ;
  assign n287 = n284 ^ n283 ^ 1'b0 ;
  assign n288 = x66 & ~n260 ;
  assign n289 = ( x66 & n282 ) | ( x66 & ~n288 ) | ( n282 & ~n288 ) ;
  assign n290 = n161 & n272 ;
  assign n291 = n289 | n290 ;
  assign n292 = n291 ^ x56 ^ 1'b0 ;
  assign n293 = ( n179 & n286 ) | ( n179 & n292 ) | ( n286 & n292 ) ;
  assign n294 = n292 ^ n286 ^ n179 ;
  assign n295 = x66 & n263 ;
  assign n296 = ( x68 & n264 ) | ( x68 & n295 ) | ( n264 & n295 ) ;
  assign n297 = n295 | n296 ;
  assign n298 = x67 & ~n260 ;
  assign n299 = ( x67 & n297 ) | ( x67 & ~n298 ) | ( n297 & ~n298 ) ;
  assign n300 = n175 & n272 ;
  assign n301 = n299 | n300 ;
  assign n302 = n301 ^ x56 ^ 1'b0 ;
  assign n303 = n302 ^ n293 ^ n221 ;
  assign n304 = ( n221 & n293 ) | ( n221 & n302 ) | ( n293 & n302 ) ;
  assign n305 = x67 & n263 ;
  assign n306 = ( x69 & n264 ) | ( x69 & n305 ) | ( n264 & n305 ) ;
  assign n307 = n305 | n306 ;
  assign n308 = x68 & ~n260 ;
  assign n309 = ( x68 & n307 ) | ( x68 & ~n308 ) | ( n307 & ~n308 ) ;
  assign n310 = n172 & n272 ;
  assign n311 = n309 | n310 ;
  assign n312 = n311 ^ x56 ^ 1'b0 ;
  assign n313 = ( n223 & n304 ) | ( n223 & n312 ) | ( n304 & n312 ) ;
  assign n314 = n312 ^ n304 ^ n223 ;
  assign n315 = x68 & n263 ;
  assign n316 = ( x70 & n264 ) | ( x70 & n315 ) | ( n264 & n315 ) ;
  assign n317 = n315 | n316 ;
  assign n318 = x69 & ~n260 ;
  assign n319 = ( x69 & n317 ) | ( x69 & ~n318 ) | ( n317 & ~n318 ) ;
  assign n320 = n168 & n272 ;
  assign n321 = n319 | n320 ;
  assign n322 = n321 ^ x56 ^ 1'b0 ;
  assign n323 = n322 ^ n313 ^ n224 ;
  assign n324 = ( n224 & n313 ) | ( n224 & n322 ) | ( n313 & n322 ) ;
  assign n325 = x62 & x63 ;
  assign n326 = ( x70 & x71 ) | ( x70 & n177 ) | ( x71 & n177 ) ;
  assign n327 = x69 & n133 ;
  assign n328 = n177 ^ x71 ^ x70 ;
  assign n329 = ( x71 & n142 ) | ( x71 & n327 ) | ( n142 & n327 ) ;
  assign n330 = x71 & n263 ;
  assign n331 = ( x73 & n264 ) | ( x73 & n330 ) | ( n264 & n330 ) ;
  assign n332 = x68 & ~n192 ;
  assign n333 = x64 & n325 ;
  assign n334 = x67 & n208 ;
  assign n335 = ( x69 & n194 ) | ( x69 & n334 ) | ( n194 & n334 ) ;
  assign n336 = n334 | n335 ;
  assign n337 = x70 & n133 ;
  assign n338 = ( x68 & ~n332 ) | ( x68 & n336 ) | ( ~n332 & n336 ) ;
  assign n339 = x66 & ~n242 ;
  assign n340 = ( x72 & n142 ) | ( x72 & n337 ) | ( n142 & n337 ) ;
  assign n341 = n337 | n340 ;
  assign n342 = x65 & ~n242 ;
  assign n343 = ( x65 & n333 ) | ( x65 & ~n342 ) | ( n333 & ~n342 ) ;
  assign n344 = n327 | n329 ;
  assign n345 = n172 & n197 ;
  assign n346 = n338 | n345 ;
  assign n347 = ( x71 & x72 ) | ( x71 & n326 ) | ( x72 & n326 ) ;
  assign n348 = ( n245 & n255 ) | ( n245 & n343 ) | ( n255 & n343 ) ;
  assign n349 = n326 ^ x72 ^ x71 ;
  assign n350 = n343 ^ n255 ^ n245 ;
  assign n351 = x71 & ~n134 ;
  assign n352 = n346 ^ x62 ^ 1'b0 ;
  assign n353 = ( x71 & n341 ) | ( x71 & ~n351 ) | ( n341 & ~n351 ) ;
  assign n354 = x65 & n325 ;
  assign n355 = x69 & n263 ;
  assign n356 = n330 | n331 ;
  assign n357 = x72 & ~n260 ;
  assign n358 = ( x72 & n356 ) | ( x72 & ~n357 ) | ( n356 & ~n357 ) ;
  assign n359 = ( x66 & ~n339 ) | ( x66 & n354 ) | ( ~n339 & n354 ) ;
  assign n360 = n359 ^ n352 ^ n348 ;
  assign n361 = n140 & n349 ;
  assign n362 = n353 | n361 ;
  assign n363 = ( n348 & n352 ) | ( n348 & n359 ) | ( n352 & n359 ) ;
  assign n364 = ( x71 & n264 ) | ( x71 & n355 ) | ( n264 & n355 ) ;
  assign n365 = n355 | n364 ;
  assign n366 = x70 & ~n134 ;
  assign n367 = n140 & n328 ;
  assign n368 = ( x72 & x73 ) | ( x72 & n347 ) | ( x73 & n347 ) ;
  assign n369 = ( x70 & n344 ) | ( x70 & ~n366 ) | ( n344 & ~n366 ) ;
  assign n370 = n347 ^ x73 ^ x72 ;
  assign n371 = n272 & n370 ;
  assign n372 = n358 | n371 ;
  assign n373 = x70 & n263 ;
  assign n374 = n367 | n369 ;
  assign n375 = n374 ^ x59 ^ 1'b0 ;
  assign n376 = ( n256 & n350 ) | ( n256 & n375 ) | ( n350 & n375 ) ;
  assign n377 = n375 ^ n350 ^ n256 ;
  assign n378 = x71 & ~n260 ;
  assign n379 = n362 ^ x59 ^ 1'b0 ;
  assign n380 = n372 ^ x56 ^ 1'b0 ;
  assign n381 = ( x72 & n264 ) | ( x72 & n373 ) | ( n264 & n373 ) ;
  assign n382 = n373 | n381 ;
  assign n383 = ( x71 & ~n378 ) | ( x71 & n382 ) | ( ~n378 & n382 ) ;
  assign n384 = n272 & n349 ;
  assign n385 = n272 & n328 ;
  assign n386 = n383 | n384 ;
  assign n387 = ( n360 & n376 ) | ( n360 & n379 ) | ( n376 & n379 ) ;
  assign n388 = n379 ^ n376 ^ n360 ;
  assign n389 = x70 & ~n260 ;
  assign n390 = ( x70 & n365 ) | ( x70 & ~n389 ) | ( n365 & ~n389 ) ;
  assign n391 = n385 | n390 ;
  assign n392 = n391 ^ x56 ^ 1'b0 ;
  assign n393 = ( n229 & n324 ) | ( n229 & n392 ) | ( n324 & n392 ) ;
  assign n394 = n386 ^ x56 ^ 1'b0 ;
  assign n395 = n394 ^ n393 ^ n240 ;
  assign n396 = ( n240 & n393 ) | ( n240 & n394 ) | ( n393 & n394 ) ;
  assign n397 = ( n254 & n380 ) | ( n254 & n396 ) | ( n380 & n396 ) ;
  assign n398 = n392 ^ n324 ^ n229 ;
  assign n399 = n396 ^ n380 ^ n254 ;
  assign n400 = x53 ^ x52 ^ 1'b0 ;
  assign n401 = x51 ^ x50 ^ 1'b0 ;
  assign n402 = n400 & n401 ;
  assign n403 = ~n400 & n401 ;
  assign n404 = x52 ^ x51 ^ 1'b0 ;
  assign n405 = ~x65 & n403 ;
  assign n406 = n139 & n402 ;
  assign n407 = ( n400 & ~n401 ) | ( n400 & n404 ) | ( ~n401 & n404 ) ;
  assign n408 = ~n404 & n407 ;
  assign n409 = x64 & n408 ;
  assign n410 = ~n401 & n404 ;
  assign n411 = x64 & n410 ;
  assign n412 = x64 & n401 ;
  assign n413 = x65 & n408 ;
  assign n414 = ( n403 & ~n405 ) | ( n403 & n411 ) | ( ~n405 & n411 ) ;
  assign n415 = ( n190 & n402 ) | ( n190 & n411 ) | ( n402 & n411 ) ;
  assign n416 = n414 | n415 ;
  assign n417 = n416 ^ x53 ^ 1'b0 ;
  assign n418 = ( x66 & n403 ) | ( x66 & n409 ) | ( n403 & n409 ) ;
  assign n419 = n409 | n418 ;
  assign n420 = x65 & ~n410 ;
  assign n421 = ( x65 & n419 ) | ( x65 & ~n420 ) | ( n419 & ~n420 ) ;
  assign n422 = n406 | n421 ;
  assign n423 = x53 & ~n412 ;
  assign n424 = n417 & n423 ;
  assign n425 = n423 ^ n417 ^ 1'b0 ;
  assign n426 = n422 ^ x53 ^ 1'b0 ;
  assign n427 = n426 ^ n424 ^ 1'b0 ;
  assign n428 = n424 & n426 ;
  assign n429 = ( x67 & n403 ) | ( x67 & n413 ) | ( n403 & n413 ) ;
  assign n430 = n413 | n429 ;
  assign n431 = x66 & ~n410 ;
  assign n432 = ( x66 & n430 ) | ( x66 & ~n431 ) | ( n430 & ~n431 ) ;
  assign n433 = n161 & n402 ;
  assign n434 = n432 | n433 ;
  assign n435 = n434 ^ x53 ^ 1'b0 ;
  assign n436 = ( n273 & n428 ) | ( n273 & n435 ) | ( n428 & n435 ) ;
  assign n437 = n435 ^ n428 ^ n273 ;
  assign n438 = x66 & n408 ;
  assign n439 = ( x68 & n403 ) | ( x68 & n438 ) | ( n403 & n438 ) ;
  assign n440 = n438 | n439 ;
  assign n441 = x67 & ~n410 ;
  assign n442 = ( x67 & n440 ) | ( x67 & ~n441 ) | ( n440 & ~n441 ) ;
  assign n443 = n175 & n402 ;
  assign n444 = n442 | n443 ;
  assign n445 = n444 ^ x53 ^ 1'b0 ;
  assign n446 = ( n285 & n436 ) | ( n285 & n445 ) | ( n436 & n445 ) ;
  assign n447 = n445 ^ n436 ^ n285 ;
  assign n448 = x67 & n408 ;
  assign n449 = ( x69 & n403 ) | ( x69 & n448 ) | ( n403 & n448 ) ;
  assign n450 = n448 | n449 ;
  assign n451 = x68 & ~n410 ;
  assign n452 = ( x68 & n450 ) | ( x68 & ~n451 ) | ( n450 & ~n451 ) ;
  assign n453 = n172 & n402 ;
  assign n454 = n452 | n453 ;
  assign n455 = n454 ^ x53 ^ 1'b0 ;
  assign n456 = n455 ^ n446 ^ n287 ;
  assign n457 = ( n287 & n446 ) | ( n287 & n455 ) | ( n446 & n455 ) ;
  assign n458 = x68 & n408 ;
  assign n459 = ( x70 & n403 ) | ( x70 & n458 ) | ( n403 & n458 ) ;
  assign n460 = n458 | n459 ;
  assign n461 = x69 & ~n410 ;
  assign n462 = ( x69 & n460 ) | ( x69 & ~n461 ) | ( n460 & ~n461 ) ;
  assign n463 = n168 & n402 ;
  assign n464 = n462 | n463 ;
  assign n465 = n464 ^ x53 ^ 1'b0 ;
  assign n466 = ( n294 & n457 ) | ( n294 & n465 ) | ( n457 & n465 ) ;
  assign n467 = n465 ^ n457 ^ n294 ;
  assign n468 = x69 & n408 ;
  assign n469 = ( x71 & n403 ) | ( x71 & n468 ) | ( n403 & n468 ) ;
  assign n470 = n468 | n469 ;
  assign n471 = x70 & ~n410 ;
  assign n472 = ( x70 & n470 ) | ( x70 & ~n471 ) | ( n470 & ~n471 ) ;
  assign n473 = n328 & n402 ;
  assign n474 = n472 | n473 ;
  assign n475 = n474 ^ x53 ^ 1'b0 ;
  assign n476 = ( n303 & n466 ) | ( n303 & n475 ) | ( n466 & n475 ) ;
  assign n477 = n475 ^ n466 ^ n303 ;
  assign n478 = x70 & n408 ;
  assign n479 = x71 & n408 ;
  assign n480 = ( x73 & n403 ) | ( x73 & n479 ) | ( n403 & n479 ) ;
  assign n481 = n479 | n480 ;
  assign n482 = ( x72 & n403 ) | ( x72 & n478 ) | ( n403 & n478 ) ;
  assign n483 = n478 | n482 ;
  assign n484 = x71 & ~n410 ;
  assign n485 = ( x71 & n483 ) | ( x71 & ~n484 ) | ( n483 & ~n484 ) ;
  assign n486 = x72 & ~n410 ;
  assign n487 = ( x72 & n481 ) | ( x72 & ~n486 ) | ( n481 & ~n486 ) ;
  assign n488 = n370 & n402 ;
  assign n489 = n487 | n488 ;
  assign n490 = x72 & n263 ;
  assign n491 = n349 & n402 ;
  assign n492 = n485 | n491 ;
  assign n493 = n492 ^ x53 ^ 1'b0 ;
  assign n494 = ( n314 & n476 ) | ( n314 & n493 ) | ( n476 & n493 ) ;
  assign n495 = n493 ^ n476 ^ n314 ;
  assign n496 = n489 ^ x53 ^ 1'b0 ;
  assign n497 = x72 & n408 ;
  assign n498 = ( x74 & n264 ) | ( x74 & n490 ) | ( n264 & n490 ) ;
  assign n499 = n490 | n498 ;
  assign n500 = ( x74 & n403 ) | ( x74 & n497 ) | ( n403 & n497 ) ;
  assign n501 = n497 | n500 ;
  assign n502 = ( n323 & n494 ) | ( n323 & n496 ) | ( n494 & n496 ) ;
  assign n503 = n496 ^ n494 ^ n323 ;
  assign n504 = n368 ^ x74 ^ x73 ;
  assign n505 = x73 & ~n410 ;
  assign n506 = ( x73 & n501 ) | ( x73 & ~n505 ) | ( n501 & ~n505 ) ;
  assign n507 = x73 & ~n260 ;
  assign n508 = ( x73 & n499 ) | ( x73 & ~n507 ) | ( n499 & ~n507 ) ;
  assign n509 = n272 & n504 ;
  assign n510 = n508 | n509 ;
  assign n511 = n402 & n504 ;
  assign n512 = n510 ^ x56 ^ 1'b0 ;
  assign n513 = n506 | n511 ;
  assign n514 = n513 ^ x53 ^ 1'b0 ;
  assign n515 = n512 ^ n397 ^ n377 ;
  assign n516 = ( n377 & n397 ) | ( n377 & n512 ) | ( n397 & n512 ) ;
  assign n517 = x73 & n408 ;
  assign n518 = ( x75 & n403 ) | ( x75 & n517 ) | ( n403 & n517 ) ;
  assign n519 = n517 | n518 ;
  assign n520 = ( x73 & x74 ) | ( x73 & n368 ) | ( x74 & n368 ) ;
  assign n521 = x74 & ~n410 ;
  assign n522 = ( x74 & n519 ) | ( x74 & ~n521 ) | ( n519 & ~n521 ) ;
  assign n523 = n514 ^ n502 ^ n398 ;
  assign n524 = ( n398 & n502 ) | ( n398 & n514 ) | ( n502 & n514 ) ;
  assign n525 = n520 ^ x75 ^ x74 ;
  assign n526 = n402 & n525 ;
  assign n527 = n522 | n526 ;
  assign n528 = n527 ^ x53 ^ 1'b0 ;
  assign n529 = n528 ^ n524 ^ n395 ;
  assign n530 = ( n395 & n524 ) | ( n395 & n528 ) | ( n524 & n528 ) ;
  assign n531 = x73 & n263 ;
  assign n532 = ( x75 & n264 ) | ( x75 & n531 ) | ( n264 & n531 ) ;
  assign n533 = n531 | n532 ;
  assign n534 = x74 & ~n260 ;
  assign n535 = ( x74 & n533 ) | ( x74 & ~n534 ) | ( n533 & ~n534 ) ;
  assign n536 = n272 & n525 ;
  assign n537 = n535 | n536 ;
  assign n538 = n537 ^ x56 ^ 1'b0 ;
  assign n539 = n538 ^ n516 ^ n388 ;
  assign n540 = ( n388 & n516 ) | ( n388 & n538 ) | ( n516 & n538 ) ;
  assign n541 = x76 & n408 ;
  assign n542 = ( x78 & n403 ) | ( x78 & n541 ) | ( n403 & n541 ) ;
  assign n543 = n541 | n542 ;
  assign n544 = x77 & ~n410 ;
  assign n545 = ( x77 & n543 ) | ( x77 & ~n544 ) | ( n543 & ~n544 ) ;
  assign n546 = ( x74 & x75 ) | ( x74 & n520 ) | ( x75 & n520 ) ;
  assign n547 = x49 ^ x48 ^ 1'b0 ;
  assign n548 = x48 ^ x47 ^ 1'b0 ;
  assign n549 = x50 ^ x49 ^ 1'b0 ;
  assign n550 = n547 & ~n548 ;
  assign n551 = n548 & ~n549 ;
  assign n552 = ~x65 & n551 ;
  assign n553 = n548 & n549 ;
  assign n554 = x64 & n550 ;
  assign n555 = ( n551 & ~n552 ) | ( n551 & n554 ) | ( ~n552 & n554 ) ;
  assign n556 = ( n190 & n553 ) | ( n190 & n554 ) | ( n553 & n554 ) ;
  assign n557 = n139 & n553 ;
  assign n558 = n555 | n556 ;
  assign n559 = x65 & ~n550 ;
  assign n560 = ( n547 & ~n548 ) | ( n547 & n549 ) | ( ~n548 & n549 ) ;
  assign n561 = ~n547 & n560 ;
  assign n562 = x64 & n561 ;
  assign n563 = ( x66 & n551 ) | ( x66 & n562 ) | ( n551 & n562 ) ;
  assign n564 = n562 | n563 ;
  assign n565 = x64 & n548 ;
  assign n566 = ( x65 & ~n559 ) | ( x65 & n564 ) | ( ~n559 & n564 ) ;
  assign n567 = x50 & ~n565 ;
  assign n568 = n557 | n566 ;
  assign n569 = n568 ^ x50 ^ 1'b0 ;
  assign n570 = n558 ^ x50 ^ 1'b0 ;
  assign n571 = n567 & n570 ;
  assign n572 = n571 ^ n569 ^ 1'b0 ;
  assign n573 = n569 & n571 ;
  assign n574 = n570 ^ n567 ^ 1'b0 ;
  assign n575 = x65 & n561 ;
  assign n576 = ( x67 & n551 ) | ( x67 & n575 ) | ( n551 & n575 ) ;
  assign n577 = n575 | n576 ;
  assign n578 = x66 & ~n550 ;
  assign n579 = ( x66 & n577 ) | ( x66 & ~n578 ) | ( n577 & ~n578 ) ;
  assign n580 = n161 & n553 ;
  assign n581 = n579 | n580 ;
  assign n582 = n581 ^ x50 ^ 1'b0 ;
  assign n583 = ( n412 & n573 ) | ( n412 & n582 ) | ( n573 & n582 ) ;
  assign n584 = n582 ^ n573 ^ n412 ;
  assign n585 = x66 & n561 ;
  assign n586 = ( x68 & n551 ) | ( x68 & n585 ) | ( n551 & n585 ) ;
  assign n587 = n585 | n586 ;
  assign n588 = x67 & ~n550 ;
  assign n589 = ( x67 & n587 ) | ( x67 & ~n588 ) | ( n587 & ~n588 ) ;
  assign n590 = n175 & n553 ;
  assign n591 = n589 | n590 ;
  assign n592 = n591 ^ x50 ^ 1'b0 ;
  assign n593 = n592 ^ n583 ^ n425 ;
  assign n594 = ( n425 & n583 ) | ( n425 & n592 ) | ( n583 & n592 ) ;
  assign n595 = x67 & n561 ;
  assign n596 = ( x69 & n551 ) | ( x69 & n595 ) | ( n551 & n595 ) ;
  assign n597 = n595 | n596 ;
  assign n598 = x68 & ~n550 ;
  assign n599 = ( x68 & n597 ) | ( x68 & ~n598 ) | ( n597 & ~n598 ) ;
  assign n600 = n172 & n553 ;
  assign n601 = n599 | n600 ;
  assign n602 = n601 ^ x50 ^ 1'b0 ;
  assign n603 = n602 ^ n594 ^ n427 ;
  assign n604 = ( n427 & n594 ) | ( n427 & n602 ) | ( n594 & n602 ) ;
  assign n605 = x68 & n561 ;
  assign n606 = ( x70 & n551 ) | ( x70 & n605 ) | ( n551 & n605 ) ;
  assign n607 = n605 | n606 ;
  assign n608 = x69 & ~n550 ;
  assign n609 = ( x69 & n607 ) | ( x69 & ~n608 ) | ( n607 & ~n608 ) ;
  assign n610 = n168 & n553 ;
  assign n611 = n609 | n610 ;
  assign n612 = n611 ^ x50 ^ 1'b0 ;
  assign n613 = n612 ^ n604 ^ n437 ;
  assign n614 = ( n437 & n604 ) | ( n437 & n612 ) | ( n604 & n612 ) ;
  assign n615 = x69 & n561 ;
  assign n616 = ( x71 & n551 ) | ( x71 & n615 ) | ( n551 & n615 ) ;
  assign n617 = n615 | n616 ;
  assign n618 = x70 & ~n550 ;
  assign n619 = ( x70 & n617 ) | ( x70 & ~n618 ) | ( n617 & ~n618 ) ;
  assign n620 = n328 & n553 ;
  assign n621 = n619 | n620 ;
  assign n622 = n621 ^ x50 ^ 1'b0 ;
  assign n623 = n622 ^ n614 ^ n447 ;
  assign n624 = ( n447 & n614 ) | ( n447 & n622 ) | ( n614 & n622 ) ;
  assign n625 = x70 & n561 ;
  assign n626 = ( x72 & n551 ) | ( x72 & n625 ) | ( n551 & n625 ) ;
  assign n627 = n625 | n626 ;
  assign n628 = x71 & ~n550 ;
  assign n629 = ( x71 & n627 ) | ( x71 & ~n628 ) | ( n627 & ~n628 ) ;
  assign n630 = n349 & n553 ;
  assign n631 = n629 | n630 ;
  assign n632 = n631 ^ x50 ^ 1'b0 ;
  assign n633 = ( n456 & n624 ) | ( n456 & n632 ) | ( n624 & n632 ) ;
  assign n634 = n632 ^ n624 ^ n456 ;
  assign n635 = x71 & n561 ;
  assign n636 = ( x73 & n551 ) | ( x73 & n635 ) | ( n551 & n635 ) ;
  assign n637 = n635 | n636 ;
  assign n638 = x72 & ~n550 ;
  assign n639 = ( x72 & n637 ) | ( x72 & ~n638 ) | ( n637 & ~n638 ) ;
  assign n640 = n370 & n553 ;
  assign n641 = n639 | n640 ;
  assign n642 = n641 ^ x50 ^ 1'b0 ;
  assign n643 = ( n467 & n633 ) | ( n467 & n642 ) | ( n633 & n642 ) ;
  assign n644 = n642 ^ n633 ^ n467 ;
  assign n645 = x73 & ~n550 ;
  assign n646 = x72 & n561 ;
  assign n647 = ( x74 & n551 ) | ( x74 & n646 ) | ( n551 & n646 ) ;
  assign n648 = n646 | n647 ;
  assign n649 = ( x73 & ~n645 ) | ( x73 & n648 ) | ( ~n645 & n648 ) ;
  assign n650 = n504 & n553 ;
  assign n651 = n649 | n650 ;
  assign n652 = x73 & n561 ;
  assign n653 = ( x75 & n551 ) | ( x75 & n652 ) | ( n551 & n652 ) ;
  assign n654 = n652 | n653 ;
  assign n655 = x74 & ~n550 ;
  assign n656 = ( x74 & n654 ) | ( x74 & ~n655 ) | ( n654 & ~n655 ) ;
  assign n657 = n525 & n553 ;
  assign n658 = n656 | n657 ;
  assign n659 = n651 ^ x50 ^ 1'b0 ;
  assign n660 = ( n477 & n643 ) | ( n477 & n659 ) | ( n643 & n659 ) ;
  assign n661 = n658 ^ x50 ^ 1'b0 ;
  assign n662 = n659 ^ n643 ^ n477 ;
  assign n663 = ( x75 & x76 ) | ( x75 & n546 ) | ( x76 & n546 ) ;
  assign n664 = n546 ^ x76 ^ x75 ;
  assign n665 = n661 ^ n660 ^ n495 ;
  assign n666 = ( n495 & n660 ) | ( n495 & n661 ) | ( n660 & n661 ) ;
  assign n667 = x74 & n561 ;
  assign n668 = ( x76 & n551 ) | ( x76 & n667 ) | ( n551 & n667 ) ;
  assign n669 = n667 | n668 ;
  assign n670 = x75 & ~n550 ;
  assign n671 = ( x75 & n669 ) | ( x75 & ~n670 ) | ( n669 & ~n670 ) ;
  assign n672 = n553 & n664 ;
  assign n673 = n671 | n672 ;
  assign n674 = n673 ^ x50 ^ 1'b0 ;
  assign n675 = n674 ^ n666 ^ n503 ;
  assign n676 = ( n503 & n666 ) | ( n503 & n674 ) | ( n666 & n674 ) ;
  assign n677 = x74 & n408 ;
  assign n678 = ( x76 & n403 ) | ( x76 & n677 ) | ( n403 & n677 ) ;
  assign n679 = n677 | n678 ;
  assign n680 = x75 & ~n410 ;
  assign n681 = ( x75 & n679 ) | ( x75 & ~n680 ) | ( n679 & ~n680 ) ;
  assign n682 = n402 & n664 ;
  assign n683 = n681 | n682 ;
  assign n684 = n683 ^ x53 ^ 1'b0 ;
  assign n685 = n684 ^ n530 ^ n399 ;
  assign n686 = ( n399 & n530 ) | ( n399 & n684 ) | ( n530 & n684 ) ;
  assign n687 = ( x76 & x77 ) | ( x76 & n663 ) | ( x77 & n663 ) ;
  assign n688 = x75 & n561 ;
  assign n689 = ( x77 & n551 ) | ( x77 & n688 ) | ( n551 & n688 ) ;
  assign n690 = n663 ^ x77 ^ x76 ;
  assign n691 = n688 | n689 ;
  assign n692 = x76 & ~n550 ;
  assign n693 = ( x76 & n691 ) | ( x76 & ~n692 ) | ( n691 & ~n692 ) ;
  assign n694 = n553 & n690 ;
  assign n695 = n693 | n694 ;
  assign n696 = n695 ^ x50 ^ 1'b0 ;
  assign n697 = n696 ^ n676 ^ n523 ;
  assign n698 = ( n523 & n676 ) | ( n523 & n696 ) | ( n676 & n696 ) ;
  assign n699 = x75 & n408 ;
  assign n700 = ( x77 & n403 ) | ( x77 & n699 ) | ( n403 & n699 ) ;
  assign n701 = n699 | n700 ;
  assign n702 = x76 & ~n410 ;
  assign n703 = ( x76 & n701 ) | ( x76 & ~n702 ) | ( n701 & ~n702 ) ;
  assign n704 = n402 & n690 ;
  assign n705 = n703 | n704 ;
  assign n706 = n705 ^ x53 ^ 1'b0 ;
  assign n707 = ( n515 & n686 ) | ( n515 & n706 ) | ( n686 & n706 ) ;
  assign n708 = n706 ^ n686 ^ n515 ;
  assign n709 = n687 ^ x78 ^ x77 ;
  assign n710 = n402 & n709 ;
  assign n711 = n545 | n710 ;
  assign n712 = n711 ^ x53 ^ 1'b0 ;
  assign n713 = ( n539 & n707 ) | ( n539 & n712 ) | ( n707 & n712 ) ;
  assign n714 = n712 ^ n707 ^ n539 ;
  assign n715 = ( x77 & x78 ) | ( x77 & n687 ) | ( x78 & n687 ) ;
  assign n716 = x76 & n561 ;
  assign n717 = ( x78 & n551 ) | ( x78 & n716 ) | ( n551 & n716 ) ;
  assign n718 = n716 | n717 ;
  assign n719 = x77 & ~n550 ;
  assign n720 = ( x77 & n718 ) | ( x77 & ~n719 ) | ( n718 & ~n719 ) ;
  assign n721 = n553 & n709 ;
  assign n722 = n720 | n721 ;
  assign n723 = n722 ^ x50 ^ 1'b0 ;
  assign n724 = ( n529 & n698 ) | ( n529 & n723 ) | ( n698 & n723 ) ;
  assign n725 = n723 ^ n698 ^ n529 ;
  assign n726 = x45 ^ x44 ^ 1'b0 ;
  assign n727 = x46 ^ x45 ^ 1'b0 ;
  assign n728 = x47 ^ x46 ^ 1'b0 ;
  assign n729 = ( ~n726 & n727 ) | ( ~n726 & n728 ) | ( n727 & n728 ) ;
  assign n730 = n726 & ~n728 ;
  assign n731 = n726 & n728 ;
  assign n732 = ~n726 & n727 ;
  assign n733 = ~x65 & n730 ;
  assign n734 = x64 & n726 ;
  assign n735 = x47 & ~n734 ;
  assign n736 = x64 & n732 ;
  assign n737 = ( n190 & n731 ) | ( n190 & n736 ) | ( n731 & n736 ) ;
  assign n738 = ( n730 & ~n733 ) | ( n730 & n736 ) | ( ~n733 & n736 ) ;
  assign n739 = n737 | n738 ;
  assign n740 = n739 ^ x47 ^ 1'b0 ;
  assign n741 = n735 & n740 ;
  assign n742 = x65 & ~n732 ;
  assign n743 = n740 ^ n735 ^ 1'b0 ;
  assign n744 = ~n727 & n729 ;
  assign n745 = x64 & n744 ;
  assign n746 = ( x66 & n730 ) | ( x66 & n745 ) | ( n730 & n745 ) ;
  assign n747 = n745 | n746 ;
  assign n748 = x65 & n744 ;
  assign n749 = ( x65 & ~n742 ) | ( x65 & n747 ) | ( ~n742 & n747 ) ;
  assign n750 = n139 & n731 ;
  assign n751 = n749 | n750 ;
  assign n752 = n751 ^ x47 ^ 1'b0 ;
  assign n753 = ( x67 & n730 ) | ( x67 & n748 ) | ( n730 & n748 ) ;
  assign n754 = n748 | n753 ;
  assign n755 = n741 & n752 ;
  assign n756 = n752 ^ n741 ^ 1'b0 ;
  assign n757 = x66 & ~n732 ;
  assign n758 = ( x66 & n754 ) | ( x66 & ~n757 ) | ( n754 & ~n757 ) ;
  assign n759 = n161 & n731 ;
  assign n760 = n758 | n759 ;
  assign n761 = n760 ^ x47 ^ 1'b0 ;
  assign n762 = n761 ^ n755 ^ n565 ;
  assign n763 = ( n565 & n755 ) | ( n565 & n761 ) | ( n755 & n761 ) ;
  assign n764 = x66 & n744 ;
  assign n765 = ( x68 & n730 ) | ( x68 & n764 ) | ( n730 & n764 ) ;
  assign n766 = n764 | n765 ;
  assign n767 = x67 & ~n732 ;
  assign n768 = ( x67 & n766 ) | ( x67 & ~n767 ) | ( n766 & ~n767 ) ;
  assign n769 = n175 & n731 ;
  assign n770 = n768 | n769 ;
  assign n771 = n770 ^ x47 ^ 1'b0 ;
  assign n772 = n771 ^ n763 ^ n574 ;
  assign n773 = ( n574 & n763 ) | ( n574 & n771 ) | ( n763 & n771 ) ;
  assign n774 = x67 & n744 ;
  assign n775 = ( x69 & n730 ) | ( x69 & n774 ) | ( n730 & n774 ) ;
  assign n776 = n774 | n775 ;
  assign n777 = x68 & ~n732 ;
  assign n778 = ( x68 & n776 ) | ( x68 & ~n777 ) | ( n776 & ~n777 ) ;
  assign n779 = n172 & n731 ;
  assign n780 = n778 | n779 ;
  assign n781 = n780 ^ x47 ^ 1'b0 ;
  assign n782 = n781 ^ n773 ^ n572 ;
  assign n783 = ( n572 & n773 ) | ( n572 & n781 ) | ( n773 & n781 ) ;
  assign n784 = x68 & n744 ;
  assign n785 = ( x70 & n730 ) | ( x70 & n784 ) | ( n730 & n784 ) ;
  assign n786 = n784 | n785 ;
  assign n787 = x69 & ~n732 ;
  assign n788 = ( x69 & n786 ) | ( x69 & ~n787 ) | ( n786 & ~n787 ) ;
  assign n789 = n168 & n731 ;
  assign n790 = n788 | n789 ;
  assign n791 = n790 ^ x47 ^ 1'b0 ;
  assign n792 = n791 ^ n783 ^ n584 ;
  assign n793 = ( n584 & n783 ) | ( n584 & n791 ) | ( n783 & n791 ) ;
  assign n794 = x69 & n744 ;
  assign n795 = ( x71 & n730 ) | ( x71 & n794 ) | ( n730 & n794 ) ;
  assign n796 = n794 | n795 ;
  assign n797 = x70 & ~n732 ;
  assign n798 = ( x70 & n796 ) | ( x70 & ~n797 ) | ( n796 & ~n797 ) ;
  assign n799 = n328 & n731 ;
  assign n800 = n798 | n799 ;
  assign n801 = n800 ^ x47 ^ 1'b0 ;
  assign n802 = n801 ^ n793 ^ n593 ;
  assign n803 = ( n593 & n793 ) | ( n593 & n801 ) | ( n793 & n801 ) ;
  assign n804 = x70 & n744 ;
  assign n805 = ( x72 & n730 ) | ( x72 & n804 ) | ( n730 & n804 ) ;
  assign n806 = n804 | n805 ;
  assign n807 = x71 & ~n732 ;
  assign n808 = ( x71 & n806 ) | ( x71 & ~n807 ) | ( n806 & ~n807 ) ;
  assign n809 = n349 & n731 ;
  assign n810 = n808 | n809 ;
  assign n811 = n810 ^ x47 ^ 1'b0 ;
  assign n812 = n811 ^ n803 ^ n603 ;
  assign n813 = ( n603 & n803 ) | ( n603 & n811 ) | ( n803 & n811 ) ;
  assign n814 = x71 & n744 ;
  assign n815 = ( x73 & n730 ) | ( x73 & n814 ) | ( n730 & n814 ) ;
  assign n816 = n814 | n815 ;
  assign n817 = x72 & ~n732 ;
  assign n818 = ( x72 & n816 ) | ( x72 & ~n817 ) | ( n816 & ~n817 ) ;
  assign n819 = n370 & n731 ;
  assign n820 = n818 | n819 ;
  assign n821 = n820 ^ x47 ^ 1'b0 ;
  assign n822 = ( n613 & n813 ) | ( n613 & n821 ) | ( n813 & n821 ) ;
  assign n823 = n821 ^ n813 ^ n613 ;
  assign n824 = x72 & n744 ;
  assign n825 = ( x74 & n730 ) | ( x74 & n824 ) | ( n730 & n824 ) ;
  assign n826 = n824 | n825 ;
  assign n827 = x73 & ~n732 ;
  assign n828 = ( x73 & n826 ) | ( x73 & ~n827 ) | ( n826 & ~n827 ) ;
  assign n829 = n504 & n731 ;
  assign n830 = n828 | n829 ;
  assign n831 = n830 ^ x47 ^ 1'b0 ;
  assign n832 = n831 ^ n822 ^ n623 ;
  assign n833 = ( n623 & n822 ) | ( n623 & n831 ) | ( n822 & n831 ) ;
  assign n834 = x73 & n744 ;
  assign n835 = ( x75 & n730 ) | ( x75 & n834 ) | ( n730 & n834 ) ;
  assign n836 = n834 | n835 ;
  assign n837 = x74 & ~n732 ;
  assign n838 = ( x74 & n836 ) | ( x74 & ~n837 ) | ( n836 & ~n837 ) ;
  assign n839 = n525 & n731 ;
  assign n840 = n838 | n839 ;
  assign n841 = n840 ^ x47 ^ 1'b0 ;
  assign n842 = n841 ^ n833 ^ n634 ;
  assign n843 = ( n634 & n833 ) | ( n634 & n841 ) | ( n833 & n841 ) ;
  assign n844 = x74 & n744 ;
  assign n845 = ( x76 & n730 ) | ( x76 & n844 ) | ( n730 & n844 ) ;
  assign n846 = n844 | n845 ;
  assign n847 = x75 & ~n732 ;
  assign n848 = ( x75 & n846 ) | ( x75 & ~n847 ) | ( n846 & ~n847 ) ;
  assign n849 = n664 & n731 ;
  assign n850 = n848 | n849 ;
  assign n851 = n850 ^ x47 ^ 1'b0 ;
  assign n852 = n851 ^ n843 ^ n644 ;
  assign n853 = ( n644 & n843 ) | ( n644 & n851 ) | ( n843 & n851 ) ;
  assign n854 = x75 & n744 ;
  assign n855 = ( x77 & n730 ) | ( x77 & n854 ) | ( n730 & n854 ) ;
  assign n856 = n854 | n855 ;
  assign n857 = x76 & ~n732 ;
  assign n858 = ( x76 & n856 ) | ( x76 & ~n857 ) | ( n856 & ~n857 ) ;
  assign n859 = n690 & n731 ;
  assign n860 = n858 | n859 ;
  assign n861 = n860 ^ x47 ^ 1'b0 ;
  assign n862 = ( n662 & n853 ) | ( n662 & n861 ) | ( n853 & n861 ) ;
  assign n863 = n861 ^ n853 ^ n662 ;
  assign n864 = x76 & n744 ;
  assign n865 = ( x78 & n730 ) | ( x78 & n864 ) | ( n730 & n864 ) ;
  assign n866 = n864 | n865 ;
  assign n867 = x77 & ~n732 ;
  assign n868 = ( x77 & n866 ) | ( x77 & ~n867 ) | ( n866 & ~n867 ) ;
  assign n869 = n709 & n731 ;
  assign n870 = n868 | n869 ;
  assign n871 = n870 ^ x47 ^ 1'b0 ;
  assign n872 = n871 ^ n862 ^ n665 ;
  assign n873 = ( n665 & n862 ) | ( n665 & n871 ) | ( n862 & n871 ) ;
  assign n874 = x43 ^ x42 ^ 1'b0 ;
  assign n875 = x42 ^ x41 ^ 1'b0 ;
  assign n876 = x44 ^ x43 ^ 1'b0 ;
  assign n877 = n874 & ~n875 ;
  assign n878 = n875 & ~n876 ;
  assign n879 = ~x65 & n878 ;
  assign n880 = n875 & n876 ;
  assign n881 = x64 & n877 ;
  assign n882 = ( n878 & ~n879 ) | ( n878 & n881 ) | ( ~n879 & n881 ) ;
  assign n883 = ( n190 & n880 ) | ( n190 & n881 ) | ( n880 & n881 ) ;
  assign n884 = n139 & n880 ;
  assign n885 = n882 | n883 ;
  assign n886 = x65 & ~n877 ;
  assign n887 = ( n874 & ~n875 ) | ( n874 & n876 ) | ( ~n875 & n876 ) ;
  assign n888 = ~n874 & n887 ;
  assign n889 = x64 & n888 ;
  assign n890 = ( x66 & n878 ) | ( x66 & n889 ) | ( n878 & n889 ) ;
  assign n891 = n889 | n890 ;
  assign n892 = x64 & n875 ;
  assign n893 = ( x65 & ~n886 ) | ( x65 & n891 ) | ( ~n886 & n891 ) ;
  assign n894 = x44 & ~n892 ;
  assign n895 = n884 | n893 ;
  assign n896 = n895 ^ x44 ^ 1'b0 ;
  assign n897 = n885 ^ x44 ^ 1'b0 ;
  assign n898 = n894 & n897 ;
  assign n899 = n898 ^ n896 ^ 1'b0 ;
  assign n900 = n896 & n898 ;
  assign n901 = n897 ^ n894 ^ 1'b0 ;
  assign n902 = x65 & n888 ;
  assign n903 = ( x67 & n878 ) | ( x67 & n902 ) | ( n878 & n902 ) ;
  assign n904 = n902 | n903 ;
  assign n905 = x66 & ~n877 ;
  assign n906 = ( x66 & n904 ) | ( x66 & ~n905 ) | ( n904 & ~n905 ) ;
  assign n907 = n161 & n880 ;
  assign n908 = n906 | n907 ;
  assign n909 = n908 ^ x44 ^ 1'b0 ;
  assign n910 = ( n734 & n900 ) | ( n734 & n909 ) | ( n900 & n909 ) ;
  assign n911 = n909 ^ n900 ^ n734 ;
  assign n912 = x66 & n888 ;
  assign n913 = ( x68 & n878 ) | ( x68 & n912 ) | ( n878 & n912 ) ;
  assign n914 = n912 | n913 ;
  assign n915 = x67 & ~n877 ;
  assign n916 = ( x67 & n914 ) | ( x67 & ~n915 ) | ( n914 & ~n915 ) ;
  assign n917 = n175 & n880 ;
  assign n918 = n916 | n917 ;
  assign n919 = n918 ^ x44 ^ 1'b0 ;
  assign n920 = n919 ^ n910 ^ n743 ;
  assign n921 = ( n743 & n910 ) | ( n743 & n919 ) | ( n910 & n919 ) ;
  assign n922 = x67 & n888 ;
  assign n923 = ( x69 & n878 ) | ( x69 & n922 ) | ( n878 & n922 ) ;
  assign n924 = n922 | n923 ;
  assign n925 = x68 & ~n877 ;
  assign n926 = ( x68 & n924 ) | ( x68 & ~n925 ) | ( n924 & ~n925 ) ;
  assign n927 = n172 & n880 ;
  assign n928 = n926 | n927 ;
  assign n929 = n928 ^ x44 ^ 1'b0 ;
  assign n930 = n929 ^ n921 ^ n756 ;
  assign n931 = ( n756 & n921 ) | ( n756 & n929 ) | ( n921 & n929 ) ;
  assign n932 = x68 & n888 ;
  assign n933 = ( x70 & n878 ) | ( x70 & n932 ) | ( n878 & n932 ) ;
  assign n934 = n932 | n933 ;
  assign n935 = x69 & ~n877 ;
  assign n936 = ( x69 & n934 ) | ( x69 & ~n935 ) | ( n934 & ~n935 ) ;
  assign n937 = n168 & n880 ;
  assign n938 = n936 | n937 ;
  assign n939 = n938 ^ x44 ^ 1'b0 ;
  assign n940 = ( n762 & n931 ) | ( n762 & n939 ) | ( n931 & n939 ) ;
  assign n941 = n939 ^ n931 ^ n762 ;
  assign n942 = x69 & n888 ;
  assign n943 = ( x71 & n878 ) | ( x71 & n942 ) | ( n878 & n942 ) ;
  assign n944 = n942 | n943 ;
  assign n945 = x70 & ~n877 ;
  assign n946 = ( x70 & n944 ) | ( x70 & ~n945 ) | ( n944 & ~n945 ) ;
  assign n947 = n328 & n880 ;
  assign n948 = n946 | n947 ;
  assign n949 = n948 ^ x44 ^ 1'b0 ;
  assign n950 = n949 ^ n940 ^ n772 ;
  assign n951 = ( n772 & n940 ) | ( n772 & n949 ) | ( n940 & n949 ) ;
  assign n952 = x70 & n888 ;
  assign n953 = ( x72 & n878 ) | ( x72 & n952 ) | ( n878 & n952 ) ;
  assign n954 = n952 | n953 ;
  assign n955 = x71 & ~n877 ;
  assign n956 = ( x71 & n954 ) | ( x71 & ~n955 ) | ( n954 & ~n955 ) ;
  assign n957 = n349 & n880 ;
  assign n958 = n956 | n957 ;
  assign n959 = n958 ^ x44 ^ 1'b0 ;
  assign n960 = n959 ^ n951 ^ n782 ;
  assign n961 = ( n782 & n951 ) | ( n782 & n959 ) | ( n951 & n959 ) ;
  assign n962 = x71 & n888 ;
  assign n963 = ( x73 & n878 ) | ( x73 & n962 ) | ( n878 & n962 ) ;
  assign n964 = n962 | n963 ;
  assign n965 = x72 & ~n877 ;
  assign n966 = ( x72 & n964 ) | ( x72 & ~n965 ) | ( n964 & ~n965 ) ;
  assign n967 = n370 & n880 ;
  assign n968 = n966 | n967 ;
  assign n969 = n968 ^ x44 ^ 1'b0 ;
  assign n970 = n969 ^ n961 ^ n792 ;
  assign n971 = ( n792 & n961 ) | ( n792 & n969 ) | ( n961 & n969 ) ;
  assign n972 = x72 & n888 ;
  assign n973 = ( x74 & n878 ) | ( x74 & n972 ) | ( n878 & n972 ) ;
  assign n974 = n972 | n973 ;
  assign n975 = x73 & ~n877 ;
  assign n976 = ( x73 & n974 ) | ( x73 & ~n975 ) | ( n974 & ~n975 ) ;
  assign n977 = n504 & n880 ;
  assign n978 = n976 | n977 ;
  assign n979 = n978 ^ x44 ^ 1'b0 ;
  assign n980 = n979 ^ n971 ^ n802 ;
  assign n981 = ( n802 & n971 ) | ( n802 & n979 ) | ( n971 & n979 ) ;
  assign n982 = x73 & n888 ;
  assign n983 = ( x75 & n878 ) | ( x75 & n982 ) | ( n878 & n982 ) ;
  assign n984 = n982 | n983 ;
  assign n985 = x74 & ~n877 ;
  assign n986 = ( x74 & n984 ) | ( x74 & ~n985 ) | ( n984 & ~n985 ) ;
  assign n987 = n525 & n880 ;
  assign n988 = n986 | n987 ;
  assign n989 = n988 ^ x44 ^ 1'b0 ;
  assign n990 = ( n812 & n981 ) | ( n812 & n989 ) | ( n981 & n989 ) ;
  assign n991 = n989 ^ n981 ^ n812 ;
  assign n992 = x74 & n888 ;
  assign n993 = ( x76 & n878 ) | ( x76 & n992 ) | ( n878 & n992 ) ;
  assign n994 = n992 | n993 ;
  assign n995 = x75 & ~n877 ;
  assign n996 = ( x75 & n994 ) | ( x75 & ~n995 ) | ( n994 & ~n995 ) ;
  assign n997 = n664 & n880 ;
  assign n998 = n996 | n997 ;
  assign n999 = n998 ^ x44 ^ 1'b0 ;
  assign n1000 = n999 ^ n990 ^ n823 ;
  assign n1001 = ( n823 & n990 ) | ( n823 & n999 ) | ( n990 & n999 ) ;
  assign n1002 = x75 & n888 ;
  assign n1003 = ( x77 & n878 ) | ( x77 & n1002 ) | ( n878 & n1002 ) ;
  assign n1004 = n1002 | n1003 ;
  assign n1005 = x76 & ~n877 ;
  assign n1006 = ( x76 & n1004 ) | ( x76 & ~n1005 ) | ( n1004 & ~n1005 ) ;
  assign n1007 = n690 & n880 ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = n1008 ^ x44 ^ 1'b0 ;
  assign n1010 = ( n832 & n1001 ) | ( n832 & n1009 ) | ( n1001 & n1009 ) ;
  assign n1011 = n1009 ^ n1001 ^ n832 ;
  assign n1012 = x77 & n744 ;
  assign n1013 = ( x79 & n730 ) | ( x79 & n1012 ) | ( n730 & n1012 ) ;
  assign n1014 = n1012 | n1013 ;
  assign n1015 = n715 ^ x79 ^ x78 ;
  assign n1016 = x78 & ~n732 ;
  assign n1017 = ( x78 & n1014 ) | ( x78 & ~n1016 ) | ( n1014 & ~n1016 ) ;
  assign n1018 = n731 & n1015 ;
  assign n1019 = n1017 | n1018 ;
  assign n1020 = n1019 ^ x47 ^ 1'b0 ;
  assign n1021 = ( n675 & n873 ) | ( n675 & n1020 ) | ( n873 & n1020 ) ;
  assign n1022 = n1020 ^ n873 ^ n675 ;
  assign n1023 = x76 & n888 ;
  assign n1024 = ( x78 & n878 ) | ( x78 & n1023 ) | ( n878 & n1023 ) ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = x77 & ~n877 ;
  assign n1027 = ( x77 & n1025 ) | ( x77 & ~n1026 ) | ( n1025 & ~n1026 ) ;
  assign n1028 = n709 & n880 ;
  assign n1029 = n1027 | n1028 ;
  assign n1030 = n1029 ^ x44 ^ 1'b0 ;
  assign n1031 = ( n842 & n1010 ) | ( n842 & n1030 ) | ( n1010 & n1030 ) ;
  assign n1032 = n1030 ^ n1010 ^ n842 ;
  assign n1033 = x77 & n888 ;
  assign n1034 = ( x79 & n878 ) | ( x79 & n1033 ) | ( n878 & n1033 ) ;
  assign n1035 = n1033 | n1034 ;
  assign n1036 = x78 & ~n877 ;
  assign n1037 = ( x78 & n1035 ) | ( x78 & ~n1036 ) | ( n1035 & ~n1036 ) ;
  assign n1038 = n880 & n1015 ;
  assign n1039 = n1037 | n1038 ;
  assign n1040 = n1039 ^ x44 ^ 1'b0 ;
  assign n1041 = ( n852 & n1031 ) | ( n852 & n1040 ) | ( n1031 & n1040 ) ;
  assign n1042 = n1040 ^ n1031 ^ n852 ;
  assign n1043 = x77 & n561 ;
  assign n1044 = ( x79 & n551 ) | ( x79 & n1043 ) | ( n551 & n1043 ) ;
  assign n1045 = ( x78 & x79 ) | ( x78 & n715 ) | ( x79 & n715 ) ;
  assign n1046 = n1043 | n1044 ;
  assign n1047 = x78 & ~n550 ;
  assign n1048 = ( x78 & n1046 ) | ( x78 & ~n1047 ) | ( n1046 & ~n1047 ) ;
  assign n1049 = n553 & n1015 ;
  assign n1050 = n1048 | n1049 ;
  assign n1051 = n1050 ^ x50 ^ 1'b0 ;
  assign n1052 = ( n685 & n724 ) | ( n685 & n1051 ) | ( n724 & n1051 ) ;
  assign n1053 = n1051 ^ n724 ^ n685 ;
  assign n1054 = x41 ^ x40 ^ 1'b0 ;
  assign n1055 = x39 ^ x38 ^ 1'b0 ;
  assign n1056 = x40 ^ x39 ^ 1'b0 ;
  assign n1057 = ( n1054 & ~n1055 ) | ( n1054 & n1056 ) | ( ~n1055 & n1056 ) ;
  assign n1058 = ~n1056 & n1057 ;
  assign n1059 = x64 & n1058 ;
  assign n1060 = ~n1055 & n1056 ;
  assign n1061 = x65 & ~n1060 ;
  assign n1062 = x64 & n1060 ;
  assign n1063 = n1054 & n1055 ;
  assign n1064 = ( n190 & n1062 ) | ( n190 & n1063 ) | ( n1062 & n1063 ) ;
  assign n1065 = ~n1054 & n1055 ;
  assign n1066 = ~x65 & n1065 ;
  assign n1067 = ( n1062 & n1065 ) | ( n1062 & ~n1066 ) | ( n1065 & ~n1066 ) ;
  assign n1068 = n1064 | n1067 ;
  assign n1069 = ( x66 & n1059 ) | ( x66 & n1065 ) | ( n1059 & n1065 ) ;
  assign n1070 = n139 & n1063 ;
  assign n1071 = n1059 | n1069 ;
  assign n1072 = ( x65 & ~n1061 ) | ( x65 & n1071 ) | ( ~n1061 & n1071 ) ;
  assign n1073 = x66 & ~n1060 ;
  assign n1074 = x65 & n1058 ;
  assign n1075 = n1070 | n1072 ;
  assign n1076 = ( x67 & n1065 ) | ( x67 & n1074 ) | ( n1065 & n1074 ) ;
  assign n1077 = n1074 | n1076 ;
  assign n1078 = n161 & n1063 ;
  assign n1079 = n1075 ^ x41 ^ 1'b0 ;
  assign n1080 = ( x66 & ~n1073 ) | ( x66 & n1077 ) | ( ~n1073 & n1077 ) ;
  assign n1081 = n1078 | n1080 ;
  assign n1082 = n1081 ^ x41 ^ 1'b0 ;
  assign n1083 = x64 & n1055 ;
  assign n1084 = n1068 ^ x41 ^ 1'b0 ;
  assign n1085 = x41 & ~n1083 ;
  assign n1086 = n1085 ^ n1084 ^ 1'b0 ;
  assign n1087 = n1084 & n1085 ;
  assign n1088 = n1087 ^ n1079 ^ 1'b0 ;
  assign n1089 = n1079 & n1087 ;
  assign n1090 = n1089 ^ n1082 ^ n892 ;
  assign n1091 = ( n892 & n1082 ) | ( n892 & n1089 ) | ( n1082 & n1089 ) ;
  assign n1092 = x66 & n1058 ;
  assign n1093 = ( x68 & n1065 ) | ( x68 & n1092 ) | ( n1065 & n1092 ) ;
  assign n1094 = n1092 | n1093 ;
  assign n1095 = x67 & ~n1060 ;
  assign n1096 = ( x67 & n1094 ) | ( x67 & ~n1095 ) | ( n1094 & ~n1095 ) ;
  assign n1097 = n175 & n1063 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = n1098 ^ x41 ^ 1'b0 ;
  assign n1100 = n1099 ^ n1091 ^ n901 ;
  assign n1101 = ( n901 & n1091 ) | ( n901 & n1099 ) | ( n1091 & n1099 ) ;
  assign n1102 = x67 & n1058 ;
  assign n1103 = ( x69 & n1065 ) | ( x69 & n1102 ) | ( n1065 & n1102 ) ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = x68 & ~n1060 ;
  assign n1106 = ( x68 & n1104 ) | ( x68 & ~n1105 ) | ( n1104 & ~n1105 ) ;
  assign n1107 = n172 & n1063 ;
  assign n1108 = n1106 | n1107 ;
  assign n1109 = n1108 ^ x41 ^ 1'b0 ;
  assign n1110 = ( n899 & n1101 ) | ( n899 & n1109 ) | ( n1101 & n1109 ) ;
  assign n1111 = n1109 ^ n1101 ^ n899 ;
  assign n1112 = x68 & n1058 ;
  assign n1113 = ( x70 & n1065 ) | ( x70 & n1112 ) | ( n1065 & n1112 ) ;
  assign n1114 = n1112 | n1113 ;
  assign n1115 = x69 & ~n1060 ;
  assign n1116 = ( x69 & n1114 ) | ( x69 & ~n1115 ) | ( n1114 & ~n1115 ) ;
  assign n1117 = n168 & n1063 ;
  assign n1118 = n1116 | n1117 ;
  assign n1119 = n1118 ^ x41 ^ 1'b0 ;
  assign n1120 = ( n911 & n1110 ) | ( n911 & n1119 ) | ( n1110 & n1119 ) ;
  assign n1121 = n1119 ^ n1110 ^ n911 ;
  assign n1122 = x69 & n1058 ;
  assign n1123 = ( x71 & n1065 ) | ( x71 & n1122 ) | ( n1065 & n1122 ) ;
  assign n1124 = n1122 | n1123 ;
  assign n1125 = x70 & ~n1060 ;
  assign n1126 = ( x70 & n1124 ) | ( x70 & ~n1125 ) | ( n1124 & ~n1125 ) ;
  assign n1127 = n328 & n1063 ;
  assign n1128 = n1126 | n1127 ;
  assign n1129 = n1128 ^ x41 ^ 1'b0 ;
  assign n1130 = n1129 ^ n1120 ^ n920 ;
  assign n1131 = ( n920 & n1120 ) | ( n920 & n1129 ) | ( n1120 & n1129 ) ;
  assign n1132 = x70 & n1058 ;
  assign n1133 = ( x72 & n1065 ) | ( x72 & n1132 ) | ( n1065 & n1132 ) ;
  assign n1134 = n1132 | n1133 ;
  assign n1135 = x71 & ~n1060 ;
  assign n1136 = ( x71 & n1134 ) | ( x71 & ~n1135 ) | ( n1134 & ~n1135 ) ;
  assign n1137 = n349 & n1063 ;
  assign n1138 = n1136 | n1137 ;
  assign n1139 = n1138 ^ x41 ^ 1'b0 ;
  assign n1140 = ( n930 & n1131 ) | ( n930 & n1139 ) | ( n1131 & n1139 ) ;
  assign n1141 = n1139 ^ n1131 ^ n930 ;
  assign n1142 = x71 & n1058 ;
  assign n1143 = ( x73 & n1065 ) | ( x73 & n1142 ) | ( n1065 & n1142 ) ;
  assign n1144 = n1142 | n1143 ;
  assign n1145 = x72 & ~n1060 ;
  assign n1146 = ( x72 & n1144 ) | ( x72 & ~n1145 ) | ( n1144 & ~n1145 ) ;
  assign n1147 = n370 & n1063 ;
  assign n1148 = n1146 | n1147 ;
  assign n1149 = n1148 ^ x41 ^ 1'b0 ;
  assign n1150 = ( n941 & n1140 ) | ( n941 & n1149 ) | ( n1140 & n1149 ) ;
  assign n1151 = n1149 ^ n1140 ^ n941 ;
  assign n1152 = x72 & n1058 ;
  assign n1153 = ( x74 & n1065 ) | ( x74 & n1152 ) | ( n1065 & n1152 ) ;
  assign n1154 = n1152 | n1153 ;
  assign n1155 = x73 & ~n1060 ;
  assign n1156 = ( x73 & n1154 ) | ( x73 & ~n1155 ) | ( n1154 & ~n1155 ) ;
  assign n1157 = n504 & n1063 ;
  assign n1158 = n1156 | n1157 ;
  assign n1159 = n1158 ^ x41 ^ 1'b0 ;
  assign n1160 = n1159 ^ n1150 ^ n950 ;
  assign n1161 = ( n950 & n1150 ) | ( n950 & n1159 ) | ( n1150 & n1159 ) ;
  assign n1162 = x73 & n1058 ;
  assign n1163 = ( x75 & n1065 ) | ( x75 & n1162 ) | ( n1065 & n1162 ) ;
  assign n1164 = n1162 | n1163 ;
  assign n1165 = x74 & ~n1060 ;
  assign n1166 = ( x74 & n1164 ) | ( x74 & ~n1165 ) | ( n1164 & ~n1165 ) ;
  assign n1167 = n525 & n1063 ;
  assign n1168 = n1166 | n1167 ;
  assign n1169 = n1168 ^ x41 ^ 1'b0 ;
  assign n1170 = n1169 ^ n1161 ^ n960 ;
  assign n1171 = ( n960 & n1161 ) | ( n960 & n1169 ) | ( n1161 & n1169 ) ;
  assign n1172 = x74 & n1058 ;
  assign n1173 = ( x76 & n1065 ) | ( x76 & n1172 ) | ( n1065 & n1172 ) ;
  assign n1174 = n1172 | n1173 ;
  assign n1175 = x75 & ~n1060 ;
  assign n1176 = ( x75 & n1174 ) | ( x75 & ~n1175 ) | ( n1174 & ~n1175 ) ;
  assign n1177 = n664 & n1063 ;
  assign n1178 = n1176 | n1177 ;
  assign n1179 = n1178 ^ x41 ^ 1'b0 ;
  assign n1180 = n1179 ^ n1171 ^ n970 ;
  assign n1181 = ( n970 & n1171 ) | ( n970 & n1179 ) | ( n1171 & n1179 ) ;
  assign n1182 = x75 & n1058 ;
  assign n1183 = ( x77 & n1065 ) | ( x77 & n1182 ) | ( n1065 & n1182 ) ;
  assign n1184 = n1182 | n1183 ;
  assign n1185 = x76 & ~n1060 ;
  assign n1186 = ( x76 & n1184 ) | ( x76 & ~n1185 ) | ( n1184 & ~n1185 ) ;
  assign n1187 = n690 & n1063 ;
  assign n1188 = n1186 | n1187 ;
  assign n1189 = n1188 ^ x41 ^ 1'b0 ;
  assign n1190 = n1189 ^ n1181 ^ n980 ;
  assign n1191 = ( n980 & n1181 ) | ( n980 & n1189 ) | ( n1181 & n1189 ) ;
  assign n1192 = x76 & n1058 ;
  assign n1193 = ( x78 & n1065 ) | ( x78 & n1192 ) | ( n1065 & n1192 ) ;
  assign n1194 = n1192 | n1193 ;
  assign n1195 = x77 & ~n1060 ;
  assign n1196 = ( x77 & n1194 ) | ( x77 & ~n1195 ) | ( n1194 & ~n1195 ) ;
  assign n1197 = n709 & n1063 ;
  assign n1198 = n1196 | n1197 ;
  assign n1199 = n1198 ^ x41 ^ 1'b0 ;
  assign n1200 = ( n991 & n1191 ) | ( n991 & n1199 ) | ( n1191 & n1199 ) ;
  assign n1201 = n1199 ^ n1191 ^ n991 ;
  assign n1202 = x77 & n1058 ;
  assign n1203 = ( x79 & n1065 ) | ( x79 & n1202 ) | ( n1065 & n1202 ) ;
  assign n1204 = n1202 | n1203 ;
  assign n1205 = x78 & ~n1060 ;
  assign n1206 = ( x78 & n1204 ) | ( x78 & ~n1205 ) | ( n1204 & ~n1205 ) ;
  assign n1207 = n1015 & n1063 ;
  assign n1208 = n1206 | n1207 ;
  assign n1209 = n1208 ^ x41 ^ 1'b0 ;
  assign n1210 = ( n1000 & n1200 ) | ( n1000 & n1209 ) | ( n1200 & n1209 ) ;
  assign n1211 = n1209 ^ n1200 ^ n1000 ;
  assign n1212 = x79 & ~n732 ;
  assign n1213 = x78 & n744 ;
  assign n1214 = ( x80 & n730 ) | ( x80 & n1213 ) | ( n730 & n1213 ) ;
  assign n1215 = n1213 | n1214 ;
  assign n1216 = n1045 ^ x80 ^ x79 ;
  assign n1217 = ( x79 & ~n1212 ) | ( x79 & n1215 ) | ( ~n1212 & n1215 ) ;
  assign n1218 = n731 & n1216 ;
  assign n1219 = n1217 | n1218 ;
  assign n1220 = n1219 ^ x47 ^ 1'b0 ;
  assign n1221 = ( n697 & n1021 ) | ( n697 & n1220 ) | ( n1021 & n1220 ) ;
  assign n1222 = n1220 ^ n1021 ^ n697 ;
  assign n1223 = x78 & n561 ;
  assign n1224 = ( x80 & n551 ) | ( x80 & n1223 ) | ( n551 & n1223 ) ;
  assign n1225 = ( x79 & x80 ) | ( x79 & n1045 ) | ( x80 & n1045 ) ;
  assign n1226 = n1223 | n1224 ;
  assign n1227 = x79 & ~n550 ;
  assign n1228 = ( x79 & n1226 ) | ( x79 & ~n1227 ) | ( n1226 & ~n1227 ) ;
  assign n1229 = n553 & n1216 ;
  assign n1230 = n1228 | n1229 ;
  assign n1231 = n1230 ^ x50 ^ 1'b0 ;
  assign n1232 = ( n708 & n1052 ) | ( n708 & n1231 ) | ( n1052 & n1231 ) ;
  assign n1233 = n1231 ^ n1052 ^ n708 ;
  assign n1234 = x78 & n1058 ;
  assign n1235 = ( x80 & n1065 ) | ( x80 & n1234 ) | ( n1065 & n1234 ) ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = x79 & ~n1060 ;
  assign n1238 = ( x79 & n1236 ) | ( x79 & ~n1237 ) | ( n1236 & ~n1237 ) ;
  assign n1239 = n1063 & n1216 ;
  assign n1240 = n1238 | n1239 ;
  assign n1241 = n1240 ^ x41 ^ 1'b0 ;
  assign n1242 = ( n1011 & n1210 ) | ( n1011 & n1241 ) | ( n1210 & n1241 ) ;
  assign n1243 = n1241 ^ n1210 ^ n1011 ;
  assign n1244 = x78 & n888 ;
  assign n1245 = ( x80 & n878 ) | ( x80 & n1244 ) | ( n878 & n1244 ) ;
  assign n1246 = n1244 | n1245 ;
  assign n1247 = x79 & ~n877 ;
  assign n1248 = ( x79 & n1246 ) | ( x79 & ~n1247 ) | ( n1246 & ~n1247 ) ;
  assign n1249 = n880 & n1216 ;
  assign n1250 = n1248 | n1249 ;
  assign n1251 = n1250 ^ x44 ^ 1'b0 ;
  assign n1252 = n1251 ^ n1041 ^ n863 ;
  assign n1253 = ( n863 & n1041 ) | ( n863 & n1251 ) | ( n1041 & n1251 ) ;
  assign n1254 = x80 & ~n732 ;
  assign n1255 = x79 & n744 ;
  assign n1256 = ( x81 & n730 ) | ( x81 & n1255 ) | ( n730 & n1255 ) ;
  assign n1257 = n1255 | n1256 ;
  assign n1258 = n1225 ^ x81 ^ x80 ;
  assign n1259 = ( x80 & ~n1254 ) | ( x80 & n1257 ) | ( ~n1254 & n1257 ) ;
  assign n1260 = n731 & n1258 ;
  assign n1261 = n1259 | n1260 ;
  assign n1262 = n1261 ^ x47 ^ 1'b0 ;
  assign n1263 = ( n725 & n1221 ) | ( n725 & n1262 ) | ( n1221 & n1262 ) ;
  assign n1264 = n1262 ^ n1221 ^ n725 ;
  assign n1265 = x79 & n561 ;
  assign n1266 = ( x81 & n551 ) | ( x81 & n1265 ) | ( n551 & n1265 ) ;
  assign n1267 = ( x80 & x81 ) | ( x80 & n1225 ) | ( x81 & n1225 ) ;
  assign n1268 = n1265 | n1266 ;
  assign n1269 = x80 & ~n550 ;
  assign n1270 = ( x80 & n1268 ) | ( x80 & ~n1269 ) | ( n1268 & ~n1269 ) ;
  assign n1271 = n553 & n1258 ;
  assign n1272 = n1270 | n1271 ;
  assign n1273 = n1272 ^ x50 ^ 1'b0 ;
  assign n1274 = ( n714 & n1232 ) | ( n714 & n1273 ) | ( n1232 & n1273 ) ;
  assign n1275 = n1273 ^ n1232 ^ n714 ;
  assign n1276 = x79 & n1058 ;
  assign n1277 = ( x81 & n1065 ) | ( x81 & n1276 ) | ( n1065 & n1276 ) ;
  assign n1278 = n1276 | n1277 ;
  assign n1279 = x80 & ~n1060 ;
  assign n1280 = ( x80 & n1278 ) | ( x80 & ~n1279 ) | ( n1278 & ~n1279 ) ;
  assign n1281 = n1063 & n1258 ;
  assign n1282 = n1280 | n1281 ;
  assign n1283 = n1282 ^ x41 ^ 1'b0 ;
  assign n1284 = ( n1032 & n1242 ) | ( n1032 & n1283 ) | ( n1242 & n1283 ) ;
  assign n1285 = n1283 ^ n1242 ^ n1032 ;
  assign n1286 = x79 & n888 ;
  assign n1287 = ( x81 & n878 ) | ( x81 & n1286 ) | ( n878 & n1286 ) ;
  assign n1288 = n1286 | n1287 ;
  assign n1289 = x80 & ~n877 ;
  assign n1290 = ( x80 & n1288 ) | ( x80 & ~n1289 ) | ( n1288 & ~n1289 ) ;
  assign n1291 = n880 & n1258 ;
  assign n1292 = n1290 | n1291 ;
  assign n1293 = n1292 ^ x44 ^ 1'b0 ;
  assign n1294 = n1293 ^ n1253 ^ n872 ;
  assign n1295 = ( n872 & n1253 ) | ( n872 & n1293 ) | ( n1253 & n1293 ) ;
  assign n1296 = x81 & ~n1060 ;
  assign n1297 = x80 & n1058 ;
  assign n1298 = ( x82 & n1065 ) | ( x82 & n1297 ) | ( n1065 & n1297 ) ;
  assign n1299 = n1297 | n1298 ;
  assign n1300 = ( x81 & ~n1296 ) | ( x81 & n1299 ) | ( ~n1296 & n1299 ) ;
  assign n1301 = n1267 ^ x82 ^ x81 ;
  assign n1302 = n1063 & n1301 ;
  assign n1303 = n1300 | n1302 ;
  assign n1304 = x80 & n888 ;
  assign n1305 = n1303 ^ x41 ^ 1'b0 ;
  assign n1306 = ( x81 & x82 ) | ( x81 & n1267 ) | ( x82 & n1267 ) ;
  assign n1307 = ( n1042 & n1284 ) | ( n1042 & n1305 ) | ( n1284 & n1305 ) ;
  assign n1308 = n1305 ^ n1284 ^ n1042 ;
  assign n1309 = x81 & ~n877 ;
  assign n1310 = ( x82 & n878 ) | ( x82 & n1304 ) | ( n878 & n1304 ) ;
  assign n1311 = n1304 | n1310 ;
  assign n1312 = ( x81 & ~n1309 ) | ( x81 & n1311 ) | ( ~n1309 & n1311 ) ;
  assign n1313 = ( x82 & x83 ) | ( x82 & n1306 ) | ( x83 & n1306 ) ;
  assign n1314 = n880 & n1301 ;
  assign n1315 = n1312 | n1314 ;
  assign n1316 = n1315 ^ x44 ^ 1'b0 ;
  assign n1317 = n1316 ^ n1295 ^ n1022 ;
  assign n1318 = ( n1022 & n1295 ) | ( n1022 & n1316 ) | ( n1295 & n1316 ) ;
  assign n1319 = x80 & n744 ;
  assign n1320 = ( x82 & n730 ) | ( x82 & n1319 ) | ( n730 & n1319 ) ;
  assign n1321 = n1319 | n1320 ;
  assign n1322 = x81 & ~n732 ;
  assign n1323 = ( x81 & n1321 ) | ( x81 & ~n1322 ) | ( n1321 & ~n1322 ) ;
  assign n1324 = n731 & n1301 ;
  assign n1325 = n1323 | n1324 ;
  assign n1326 = n1325 ^ x47 ^ 1'b0 ;
  assign n1327 = n1326 ^ n1263 ^ n1053 ;
  assign n1328 = ( n1053 & n1263 ) | ( n1053 & n1326 ) | ( n1263 & n1326 ) ;
  assign n1329 = n1306 ^ x83 ^ x82 ;
  assign n1330 = x81 & n888 ;
  assign n1331 = ( x83 & n878 ) | ( x83 & n1330 ) | ( n878 & n1330 ) ;
  assign n1332 = n1330 | n1331 ;
  assign n1333 = x82 & ~n877 ;
  assign n1334 = ( x82 & n1332 ) | ( x82 & ~n1333 ) | ( n1332 & ~n1333 ) ;
  assign n1335 = n880 & n1329 ;
  assign n1336 = n1334 | n1335 ;
  assign n1337 = n1336 ^ x44 ^ 1'b0 ;
  assign n1338 = ( n1222 & n1318 ) | ( n1222 & n1337 ) | ( n1318 & n1337 ) ;
  assign n1339 = n1337 ^ n1318 ^ n1222 ;
  assign n1340 = x82 & n744 ;
  assign n1341 = x83 & ~n732 ;
  assign n1342 = ( x84 & n730 ) | ( x84 & n1340 ) | ( n730 & n1340 ) ;
  assign n1343 = n1340 | n1342 ;
  assign n1344 = ( x83 & ~n1341 ) | ( x83 & n1343 ) | ( ~n1341 & n1343 ) ;
  assign n1345 = x81 & n744 ;
  assign n1346 = ( x83 & n730 ) | ( x83 & n1345 ) | ( n730 & n1345 ) ;
  assign n1347 = n1345 | n1346 ;
  assign n1348 = x82 & ~n732 ;
  assign n1349 = ( x82 & n1347 ) | ( x82 & ~n1348 ) | ( n1347 & ~n1348 ) ;
  assign n1350 = n731 & n1329 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = n1351 ^ x47 ^ 1'b0 ;
  assign n1353 = n1352 ^ n1328 ^ n1233 ;
  assign n1354 = ( n1233 & n1328 ) | ( n1233 & n1352 ) | ( n1328 & n1352 ) ;
  assign n1355 = n1313 ^ x84 ^ x83 ;
  assign n1356 = ( x83 & x84 ) | ( x83 & n1313 ) | ( x84 & n1313 ) ;
  assign n1357 = n731 & n1355 ;
  assign n1358 = n1344 | n1357 ;
  assign n1359 = n1358 ^ x47 ^ 1'b0 ;
  assign n1360 = ( n1275 & n1354 ) | ( n1275 & n1359 ) | ( n1354 & n1359 ) ;
  assign n1361 = n1359 ^ n1354 ^ n1275 ;
  assign n1362 = x82 & n888 ;
  assign n1363 = ( x84 & n878 ) | ( x84 & n1362 ) | ( n878 & n1362 ) ;
  assign n1364 = n1362 | n1363 ;
  assign n1365 = x83 & ~n877 ;
  assign n1366 = ( x83 & n1364 ) | ( x83 & ~n1365 ) | ( n1364 & ~n1365 ) ;
  assign n1367 = n880 & n1355 ;
  assign n1368 = n1366 | n1367 ;
  assign n1369 = n1368 ^ x44 ^ 1'b0 ;
  assign n1370 = n1369 ^ n1338 ^ n1264 ;
  assign n1371 = ( n1264 & n1338 ) | ( n1264 & n1369 ) | ( n1338 & n1369 ) ;
  assign n1372 = x81 & n1058 ;
  assign n1373 = ( x83 & n1065 ) | ( x83 & n1372 ) | ( n1065 & n1372 ) ;
  assign n1374 = n1372 | n1373 ;
  assign n1375 = x82 & ~n1060 ;
  assign n1376 = ( x82 & n1374 ) | ( x82 & ~n1375 ) | ( n1374 & ~n1375 ) ;
  assign n1377 = n1063 & n1329 ;
  assign n1378 = n1376 | n1377 ;
  assign n1379 = n1378 ^ x41 ^ 1'b0 ;
  assign n1380 = ( n1252 & n1307 ) | ( n1252 & n1379 ) | ( n1307 & n1379 ) ;
  assign n1381 = n1379 ^ n1307 ^ n1252 ;
  assign n1382 = x82 & n1058 ;
  assign n1383 = ( x84 & n1065 ) | ( x84 & n1382 ) | ( n1065 & n1382 ) ;
  assign n1384 = n1382 | n1383 ;
  assign n1385 = x83 & ~n1060 ;
  assign n1386 = ( x83 & n1384 ) | ( x83 & ~n1385 ) | ( n1384 & ~n1385 ) ;
  assign n1387 = n1063 & n1355 ;
  assign n1388 = n1386 | n1387 ;
  assign n1389 = n1388 ^ x41 ^ 1'b0 ;
  assign n1390 = n1389 ^ n1380 ^ n1294 ;
  assign n1391 = ( n1294 & n1380 ) | ( n1294 & n1389 ) | ( n1380 & n1389 ) ;
  assign n1392 = n1356 ^ x85 ^ x84 ;
  assign n1393 = n880 & n1392 ;
  assign n1394 = x83 & n888 ;
  assign n1395 = ( x85 & n878 ) | ( x85 & n1394 ) | ( n878 & n1394 ) ;
  assign n1396 = n1394 | n1395 ;
  assign n1397 = x84 & ~n877 ;
  assign n1398 = ( x84 & n1396 ) | ( x84 & ~n1397 ) | ( n1396 & ~n1397 ) ;
  assign n1399 = n1393 | n1398 ;
  assign n1400 = n1399 ^ x44 ^ 1'b0 ;
  assign n1401 = n1400 ^ n1371 ^ n1327 ;
  assign n1402 = ( n1327 & n1371 ) | ( n1327 & n1400 ) | ( n1371 & n1400 ) ;
  assign n1403 = x83 & n1058 ;
  assign n1404 = ( x85 & n1065 ) | ( x85 & n1403 ) | ( n1065 & n1403 ) ;
  assign n1405 = n1403 | n1404 ;
  assign n1406 = n1063 & n1392 ;
  assign n1407 = x84 & ~n1060 ;
  assign n1408 = ( x84 & n1405 ) | ( x84 & ~n1407 ) | ( n1405 & ~n1407 ) ;
  assign n1409 = n1406 | n1408 ;
  assign n1410 = x84 & n888 ;
  assign n1411 = ( x86 & n878 ) | ( x86 & n1410 ) | ( n878 & n1410 ) ;
  assign n1412 = n1410 | n1411 ;
  assign n1413 = n1409 ^ x41 ^ 1'b0 ;
  assign n1414 = ( n1317 & n1391 ) | ( n1317 & n1413 ) | ( n1391 & n1413 ) ;
  assign n1415 = n1413 ^ n1391 ^ n1317 ;
  assign n1416 = x85 & ~n877 ;
  assign n1417 = ( x85 & n1412 ) | ( x85 & ~n1416 ) | ( n1412 & ~n1416 ) ;
  assign n1418 = ( x84 & x85 ) | ( x84 & n1356 ) | ( x85 & n1356 ) ;
  assign n1419 = n1418 ^ x86 ^ x85 ;
  assign n1420 = n880 & n1419 ;
  assign n1421 = n1417 | n1420 ;
  assign n1422 = ( x85 & x86 ) | ( x85 & n1418 ) | ( x86 & n1418 ) ;
  assign n1423 = n1421 ^ x44 ^ 1'b0 ;
  assign n1424 = n1423 ^ n1402 ^ n1353 ;
  assign n1425 = ( n1353 & n1402 ) | ( n1353 & n1423 ) | ( n1402 & n1423 ) ;
  assign n1426 = x84 & n1058 ;
  assign n1427 = ( x86 & n1065 ) | ( x86 & n1426 ) | ( n1065 & n1426 ) ;
  assign n1428 = n1426 | n1427 ;
  assign n1429 = x85 & ~n1060 ;
  assign n1430 = ( x85 & n1428 ) | ( x85 & ~n1429 ) | ( n1428 & ~n1429 ) ;
  assign n1431 = n1063 & n1419 ;
  assign n1432 = n1430 | n1431 ;
  assign n1433 = n1432 ^ x41 ^ 1'b0 ;
  assign n1434 = n1433 ^ n1414 ^ n1339 ;
  assign n1435 = ( n1339 & n1414 ) | ( n1339 & n1433 ) | ( n1414 & n1433 ) ;
  assign n1436 = x68 & n208 ;
  assign n1437 = ( x70 & n194 ) | ( x70 & n1436 ) | ( n194 & n1436 ) ;
  assign n1438 = x67 & ~n242 ;
  assign n1439 = n1436 | n1437 ;
  assign n1440 = x71 & n133 ;
  assign n1441 = x66 & n325 ;
  assign n1442 = ( x67 & ~n1438 ) | ( x67 & n1441 ) | ( ~n1438 & n1441 ) ;
  assign n1443 = x69 & ~n192 ;
  assign n1444 = ( x69 & n1439 ) | ( x69 & ~n1443 ) | ( n1439 & ~n1443 ) ;
  assign n1445 = ( n168 & n197 ) | ( n168 & n1444 ) | ( n197 & n1444 ) ;
  assign n1446 = n1444 | n1445 ;
  assign n1447 = n1446 ^ x62 ^ 1'b0 ;
  assign n1448 = n1447 ^ n1442 ^ x2 ;
  assign n1449 = ( x2 & n1442 ) | ( x2 & n1447 ) | ( n1442 & n1447 ) ;
  assign n1450 = ( x73 & n142 ) | ( x73 & n1440 ) | ( n142 & n1440 ) ;
  assign n1451 = n1440 | n1450 ;
  assign n1452 = x72 & ~n134 ;
  assign n1453 = ( x72 & n1451 ) | ( x72 & ~n1452 ) | ( n1451 & ~n1452 ) ;
  assign n1454 = n140 & n370 ;
  assign n1455 = n1453 | n1454 ;
  assign n1456 = n1455 ^ x59 ^ 1'b0 ;
  assign n1457 = n1456 ^ n1448 ^ n363 ;
  assign n1458 = ( n363 & n1448 ) | ( n363 & n1456 ) | ( n1448 & n1456 ) ;
  assign n1459 = x74 & n263 ;
  assign n1460 = ( x76 & n264 ) | ( x76 & n1459 ) | ( n264 & n1459 ) ;
  assign n1461 = n1459 | n1460 ;
  assign n1462 = x75 & ~n260 ;
  assign n1463 = ( x75 & n1461 ) | ( x75 & ~n1462 ) | ( n1461 & ~n1462 ) ;
  assign n1464 = n272 & n664 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = n1465 ^ x56 ^ 1'b0 ;
  assign n1467 = ( n387 & n1457 ) | ( n387 & n1466 ) | ( n1457 & n1466 ) ;
  assign n1468 = n1466 ^ n1457 ^ n387 ;
  assign n1469 = x77 & n408 ;
  assign n1470 = ( x79 & n403 ) | ( x79 & n1469 ) | ( n403 & n1469 ) ;
  assign n1471 = n1469 | n1470 ;
  assign n1472 = x78 & ~n410 ;
  assign n1473 = ( x78 & n1471 ) | ( x78 & ~n1472 ) | ( n1471 & ~n1472 ) ;
  assign n1474 = n402 & n1015 ;
  assign n1475 = n1473 | n1474 ;
  assign n1476 = n1475 ^ x53 ^ 1'b0 ;
  assign n1477 = ( n540 & n1468 ) | ( n540 & n1476 ) | ( n1468 & n1476 ) ;
  assign n1478 = n1476 ^ n1468 ^ n540 ;
  assign n1479 = x85 & n888 ;
  assign n1480 = ( x87 & n878 ) | ( x87 & n1479 ) | ( n878 & n1479 ) ;
  assign n1481 = n1479 | n1480 ;
  assign n1482 = x86 & ~n877 ;
  assign n1483 = ( x86 & n1481 ) | ( x86 & ~n1482 ) | ( n1481 & ~n1482 ) ;
  assign n1484 = n1422 ^ x87 ^ x86 ;
  assign n1485 = n880 & n1484 ;
  assign n1486 = n1483 | n1485 ;
  assign n1487 = n1486 ^ x44 ^ 1'b0 ;
  assign n1488 = n1487 ^ n1425 ^ n1361 ;
  assign n1489 = ( n1361 & n1425 ) | ( n1361 & n1487 ) | ( n1425 & n1487 ) ;
  assign n1490 = x85 & n1058 ;
  assign n1491 = ( x87 & n1065 ) | ( x87 & n1490 ) | ( n1065 & n1490 ) ;
  assign n1492 = n1490 | n1491 ;
  assign n1493 = x86 & ~n1060 ;
  assign n1494 = ( x86 & n1492 ) | ( x86 & ~n1493 ) | ( n1492 & ~n1493 ) ;
  assign n1495 = ( x86 & x87 ) | ( x86 & n1422 ) | ( x87 & n1422 ) ;
  assign n1496 = n1063 & n1484 ;
  assign n1497 = n1494 | n1496 ;
  assign n1498 = n1497 ^ x41 ^ 1'b0 ;
  assign n1499 = ( n1370 & n1435 ) | ( n1370 & n1498 ) | ( n1435 & n1498 ) ;
  assign n1500 = n1498 ^ n1435 ^ n1370 ;
  assign n1501 = x80 & n561 ;
  assign n1502 = ( x82 & n551 ) | ( x82 & n1501 ) | ( n551 & n1501 ) ;
  assign n1503 = n1501 | n1502 ;
  assign n1504 = x81 & ~n550 ;
  assign n1505 = ( x81 & n1503 ) | ( x81 & ~n1504 ) | ( n1503 & ~n1504 ) ;
  assign n1506 = n553 & n1301 ;
  assign n1507 = n1505 | n1506 ;
  assign n1508 = n1507 ^ x50 ^ 1'b0 ;
  assign n1509 = ( n713 & n1478 ) | ( n713 & n1508 ) | ( n1478 & n1508 ) ;
  assign n1510 = n1508 ^ n1478 ^ n713 ;
  assign n1511 = x83 & n744 ;
  assign n1512 = ( x85 & n730 ) | ( x85 & n1511 ) | ( n730 & n1511 ) ;
  assign n1513 = n1511 | n1512 ;
  assign n1514 = x84 & ~n732 ;
  assign n1515 = ( x84 & n1513 ) | ( x84 & ~n1514 ) | ( n1513 & ~n1514 ) ;
  assign n1516 = n731 & n1392 ;
  assign n1517 = n1515 | n1516 ;
  assign n1518 = n1517 ^ x47 ^ 1'b0 ;
  assign n1519 = ( n1274 & n1510 ) | ( n1274 & n1518 ) | ( n1510 & n1518 ) ;
  assign n1520 = n1518 ^ n1510 ^ n1274 ;
  assign n1521 = x69 & n208 ;
  assign n1522 = ( x71 & n194 ) | ( x71 & n1521 ) | ( n194 & n1521 ) ;
  assign n1523 = x70 & ~n192 ;
  assign n1524 = x68 & ~n242 ;
  assign n1525 = n1521 | n1522 ;
  assign n1526 = ( x70 & ~n1523 ) | ( x70 & n1525 ) | ( ~n1523 & n1525 ) ;
  assign n1527 = n197 & n328 ;
  assign n1528 = x72 & n133 ;
  assign n1529 = n1526 | n1527 ;
  assign n1530 = ( x74 & n142 ) | ( x74 & n1528 ) | ( n142 & n1528 ) ;
  assign n1531 = n1528 | n1530 ;
  assign n1532 = x67 & n325 ;
  assign n1533 = n1529 ^ x62 ^ 1'b0 ;
  assign n1534 = ( x68 & ~n1524 ) | ( x68 & n1532 ) | ( ~n1524 & n1532 ) ;
  assign n1535 = ( x2 & n1533 ) | ( x2 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1536 = n1534 ^ n1533 ^ x2 ;
  assign n1537 = x73 & ~n134 ;
  assign n1538 = ( x73 & n1531 ) | ( x73 & ~n1537 ) | ( n1531 & ~n1537 ) ;
  assign n1539 = n140 & n504 ;
  assign n1540 = n1538 | n1539 ;
  assign n1541 = n1540 ^ x59 ^ 1'b0 ;
  assign n1542 = ( n1449 & n1536 ) | ( n1449 & n1541 ) | ( n1536 & n1541 ) ;
  assign n1543 = n1541 ^ n1536 ^ n1449 ;
  assign n1544 = x75 & n263 ;
  assign n1545 = ( x77 & n264 ) | ( x77 & n1544 ) | ( n264 & n1544 ) ;
  assign n1546 = n1544 | n1545 ;
  assign n1547 = x76 & ~n260 ;
  assign n1548 = ( x76 & n1546 ) | ( x76 & ~n1547 ) | ( n1546 & ~n1547 ) ;
  assign n1549 = n272 & n690 ;
  assign n1550 = n1548 | n1549 ;
  assign n1551 = n1550 ^ x56 ^ 1'b0 ;
  assign n1552 = ( n1458 & n1543 ) | ( n1458 & n1551 ) | ( n1543 & n1551 ) ;
  assign n1553 = n1551 ^ n1543 ^ n1458 ;
  assign n1554 = x78 & n408 ;
  assign n1555 = ( x80 & n403 ) | ( x80 & n1554 ) | ( n403 & n1554 ) ;
  assign n1556 = n1554 | n1555 ;
  assign n1557 = x79 & ~n410 ;
  assign n1558 = ( x79 & n1556 ) | ( x79 & ~n1557 ) | ( n1556 & ~n1557 ) ;
  assign n1559 = n402 & n1216 ;
  assign n1560 = n1558 | n1559 ;
  assign n1561 = n1560 ^ x53 ^ 1'b0 ;
  assign n1562 = n1561 ^ n1553 ^ n1467 ;
  assign n1563 = ( n1467 & n1553 ) | ( n1467 & n1561 ) | ( n1553 & n1561 ) ;
  assign n1564 = x86 & n888 ;
  assign n1565 = ( x88 & n878 ) | ( x88 & n1564 ) | ( n878 & n1564 ) ;
  assign n1566 = n1564 | n1565 ;
  assign n1567 = x87 & ~n877 ;
  assign n1568 = ( x87 & n1566 ) | ( x87 & ~n1567 ) | ( n1566 & ~n1567 ) ;
  assign n1569 = n1495 ^ x88 ^ x87 ;
  assign n1570 = n880 & n1569 ;
  assign n1571 = n1568 | n1570 ;
  assign n1572 = n1571 ^ x44 ^ 1'b0 ;
  assign n1573 = n1572 ^ n1520 ^ n1360 ;
  assign n1574 = ( n1360 & n1520 ) | ( n1360 & n1572 ) | ( n1520 & n1572 ) ;
  assign n1575 = x86 & n1058 ;
  assign n1576 = ( x88 & n1065 ) | ( x88 & n1575 ) | ( n1065 & n1575 ) ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = x87 & ~n1060 ;
  assign n1579 = ( x87 & n1577 ) | ( x87 & ~n1578 ) | ( n1577 & ~n1578 ) ;
  assign n1580 = ( x87 & x88 ) | ( x87 & n1495 ) | ( x88 & n1495 ) ;
  assign n1581 = n1063 & n1569 ;
  assign n1582 = n1579 | n1581 ;
  assign n1583 = n1582 ^ x41 ^ 1'b0 ;
  assign n1584 = ( n1401 & n1499 ) | ( n1401 & n1583 ) | ( n1499 & n1583 ) ;
  assign n1585 = n1583 ^ n1499 ^ n1401 ;
  assign n1586 = x81 & n561 ;
  assign n1587 = ( x83 & n551 ) | ( x83 & n1586 ) | ( n551 & n1586 ) ;
  assign n1588 = n1586 | n1587 ;
  assign n1589 = x82 & ~n550 ;
  assign n1590 = ( x82 & n1588 ) | ( x82 & ~n1589 ) | ( n1588 & ~n1589 ) ;
  assign n1591 = n553 & n1329 ;
  assign n1592 = n1590 | n1591 ;
  assign n1593 = n1592 ^ x50 ^ 1'b0 ;
  assign n1594 = ( n1477 & n1562 ) | ( n1477 & n1593 ) | ( n1562 & n1593 ) ;
  assign n1595 = n1593 ^ n1562 ^ n1477 ;
  assign n1596 = x84 & n744 ;
  assign n1597 = ( x86 & n730 ) | ( x86 & n1596 ) | ( n730 & n1596 ) ;
  assign n1598 = n1596 | n1597 ;
  assign n1599 = x85 & ~n732 ;
  assign n1600 = ( x85 & n1598 ) | ( x85 & ~n1599 ) | ( n1598 & ~n1599 ) ;
  assign n1601 = n731 & n1419 ;
  assign n1602 = n1600 | n1601 ;
  assign n1603 = n1602 ^ x47 ^ 1'b0 ;
  assign n1604 = ( n1509 & n1595 ) | ( n1509 & n1603 ) | ( n1595 & n1603 ) ;
  assign n1605 = n1603 ^ n1595 ^ n1509 ;
  assign n1606 = x70 & n208 ;
  assign n1607 = ( x72 & n194 ) | ( x72 & n1606 ) | ( n194 & n1606 ) ;
  assign n1608 = x71 & ~n192 ;
  assign n1609 = x69 & ~n242 ;
  assign n1610 = n1606 | n1607 ;
  assign n1611 = ( x71 & ~n1608 ) | ( x71 & n1610 ) | ( ~n1608 & n1610 ) ;
  assign n1612 = n197 & n349 ;
  assign n1613 = x73 & n133 ;
  assign n1614 = n1611 | n1612 ;
  assign n1615 = ( x75 & n142 ) | ( x75 & n1613 ) | ( n142 & n1613 ) ;
  assign n1616 = n1613 | n1615 ;
  assign n1617 = x68 & n325 ;
  assign n1618 = n1614 ^ x62 ^ 1'b0 ;
  assign n1619 = ( x69 & ~n1609 ) | ( x69 & n1617 ) | ( ~n1609 & n1617 ) ;
  assign n1620 = ( x2 & n1618 ) | ( x2 & n1619 ) | ( n1618 & n1619 ) ;
  assign n1621 = n1619 ^ n1618 ^ x2 ;
  assign n1622 = x74 & ~n134 ;
  assign n1623 = ( x74 & n1616 ) | ( x74 & ~n1622 ) | ( n1616 & ~n1622 ) ;
  assign n1624 = n140 & n525 ;
  assign n1625 = n1623 | n1624 ;
  assign n1626 = n1625 ^ x59 ^ 1'b0 ;
  assign n1627 = ( n1535 & n1621 ) | ( n1535 & n1626 ) | ( n1621 & n1626 ) ;
  assign n1628 = n1626 ^ n1621 ^ n1535 ;
  assign n1629 = x76 & n263 ;
  assign n1630 = ( x78 & n264 ) | ( x78 & n1629 ) | ( n264 & n1629 ) ;
  assign n1631 = n1629 | n1630 ;
  assign n1632 = x77 & ~n260 ;
  assign n1633 = ( x77 & n1631 ) | ( x77 & ~n1632 ) | ( n1631 & ~n1632 ) ;
  assign n1634 = n272 & n709 ;
  assign n1635 = n1633 | n1634 ;
  assign n1636 = n1635 ^ x56 ^ 1'b0 ;
  assign n1637 = ( n1542 & n1628 ) | ( n1542 & n1636 ) | ( n1628 & n1636 ) ;
  assign n1638 = n1636 ^ n1628 ^ n1542 ;
  assign n1639 = x79 & n408 ;
  assign n1640 = ( x81 & n403 ) | ( x81 & n1639 ) | ( n403 & n1639 ) ;
  assign n1641 = n1639 | n1640 ;
  assign n1642 = x80 & ~n410 ;
  assign n1643 = ( x80 & n1641 ) | ( x80 & ~n1642 ) | ( n1641 & ~n1642 ) ;
  assign n1644 = n402 & n1258 ;
  assign n1645 = n1643 | n1644 ;
  assign n1646 = n1645 ^ x53 ^ 1'b0 ;
  assign n1647 = n1646 ^ n1638 ^ n1552 ;
  assign n1648 = ( n1552 & n1638 ) | ( n1552 & n1646 ) | ( n1638 & n1646 ) ;
  assign n1649 = x87 & n888 ;
  assign n1650 = ( x89 & n878 ) | ( x89 & n1649 ) | ( n878 & n1649 ) ;
  assign n1651 = n1649 | n1650 ;
  assign n1652 = x88 & ~n877 ;
  assign n1653 = ( x88 & n1651 ) | ( x88 & ~n1652 ) | ( n1651 & ~n1652 ) ;
  assign n1654 = n1580 ^ x89 ^ x88 ;
  assign n1655 = n880 & n1654 ;
  assign n1656 = n1653 | n1655 ;
  assign n1657 = n1656 ^ x44 ^ 1'b0 ;
  assign n1658 = n1657 ^ n1605 ^ n1519 ;
  assign n1659 = ( n1519 & n1605 ) | ( n1519 & n1657 ) | ( n1605 & n1657 ) ;
  assign n1660 = x87 & n1058 ;
  assign n1661 = ( x89 & n1065 ) | ( x89 & n1660 ) | ( n1065 & n1660 ) ;
  assign n1662 = n1660 | n1661 ;
  assign n1663 = x88 & ~n1060 ;
  assign n1664 = ( x88 & n1662 ) | ( x88 & ~n1663 ) | ( n1662 & ~n1663 ) ;
  assign n1665 = ( x88 & x89 ) | ( x88 & n1580 ) | ( x89 & n1580 ) ;
  assign n1666 = n1063 & n1654 ;
  assign n1667 = n1664 | n1666 ;
  assign n1668 = n1667 ^ x41 ^ 1'b0 ;
  assign n1669 = ( n1424 & n1584 ) | ( n1424 & n1668 ) | ( n1584 & n1668 ) ;
  assign n1670 = n1668 ^ n1584 ^ n1424 ;
  assign n1671 = x82 & n561 ;
  assign n1672 = ( x84 & n551 ) | ( x84 & n1671 ) | ( n551 & n1671 ) ;
  assign n1673 = n1671 | n1672 ;
  assign n1674 = x83 & ~n550 ;
  assign n1675 = ( x83 & n1673 ) | ( x83 & ~n1674 ) | ( n1673 & ~n1674 ) ;
  assign n1676 = n553 & n1355 ;
  assign n1677 = n1675 | n1676 ;
  assign n1678 = n1677 ^ x50 ^ 1'b0 ;
  assign n1679 = ( n1563 & n1647 ) | ( n1563 & n1678 ) | ( n1647 & n1678 ) ;
  assign n1680 = n1678 ^ n1647 ^ n1563 ;
  assign n1681 = x85 & n744 ;
  assign n1682 = ( x87 & n730 ) | ( x87 & n1681 ) | ( n730 & n1681 ) ;
  assign n1683 = n1681 | n1682 ;
  assign n1684 = x86 & ~n732 ;
  assign n1685 = ( x86 & n1683 ) | ( x86 & ~n1684 ) | ( n1683 & ~n1684 ) ;
  assign n1686 = n731 & n1484 ;
  assign n1687 = n1685 | n1686 ;
  assign n1688 = n1687 ^ x47 ^ 1'b0 ;
  assign n1689 = ( n1594 & n1680 ) | ( n1594 & n1688 ) | ( n1680 & n1688 ) ;
  assign n1690 = n1688 ^ n1680 ^ n1594 ;
  assign n1691 = x72 & ~n192 ;
  assign n1692 = x71 & n208 ;
  assign n1693 = x69 & n325 ;
  assign n1694 = ( x73 & n194 ) | ( x73 & n1692 ) | ( n194 & n1692 ) ;
  assign n1695 = n1692 | n1694 ;
  assign n1696 = ( x72 & ~n1691 ) | ( x72 & n1695 ) | ( ~n1691 & n1695 ) ;
  assign n1697 = n197 & n370 ;
  assign n1698 = n1696 | n1697 ;
  assign n1699 = n1698 ^ x62 ^ 1'b0 ;
  assign n1700 = x70 & ~n242 ;
  assign n1701 = ( x70 & n1693 ) | ( x70 & ~n1700 ) | ( n1693 & ~n1700 ) ;
  assign n1702 = n1701 ^ x5 ^ x2 ;
  assign n1703 = ( n1620 & n1699 ) | ( n1620 & n1702 ) | ( n1699 & n1702 ) ;
  assign n1704 = n1702 ^ n1699 ^ n1620 ;
  assign n1705 = x74 & n133 ;
  assign n1706 = ( x76 & n142 ) | ( x76 & n1705 ) | ( n142 & n1705 ) ;
  assign n1707 = n1705 | n1706 ;
  assign n1708 = x75 & ~n134 ;
  assign n1709 = ( x75 & n1707 ) | ( x75 & ~n1708 ) | ( n1707 & ~n1708 ) ;
  assign n1710 = n140 & n664 ;
  assign n1711 = n1709 | n1710 ;
  assign n1712 = n1711 ^ x59 ^ 1'b0 ;
  assign n1713 = ( n1627 & n1704 ) | ( n1627 & n1712 ) | ( n1704 & n1712 ) ;
  assign n1714 = n1712 ^ n1704 ^ n1627 ;
  assign n1715 = x77 & n263 ;
  assign n1716 = ( x2 & x5 ) | ( x2 & ~n1701 ) | ( x5 & ~n1701 ) ;
  assign n1717 = ( x79 & n264 ) | ( x79 & n1715 ) | ( n264 & n1715 ) ;
  assign n1718 = n1715 | n1717 ;
  assign n1719 = x78 & ~n260 ;
  assign n1720 = ( x78 & n1718 ) | ( x78 & ~n1719 ) | ( n1718 & ~n1719 ) ;
  assign n1721 = n272 & n1015 ;
  assign n1722 = n1720 | n1721 ;
  assign n1723 = n1722 ^ x56 ^ 1'b0 ;
  assign n1724 = ( n1637 & n1714 ) | ( n1637 & n1723 ) | ( n1714 & n1723 ) ;
  assign n1725 = n1723 ^ n1714 ^ n1637 ;
  assign n1726 = x80 & n408 ;
  assign n1727 = ( x82 & n403 ) | ( x82 & n1726 ) | ( n403 & n1726 ) ;
  assign n1728 = n1726 | n1727 ;
  assign n1729 = x81 & ~n410 ;
  assign n1730 = ( x81 & n1728 ) | ( x81 & ~n1729 ) | ( n1728 & ~n1729 ) ;
  assign n1731 = n402 & n1301 ;
  assign n1732 = n1730 | n1731 ;
  assign n1733 = n1732 ^ x53 ^ 1'b0 ;
  assign n1734 = n1733 ^ n1725 ^ n1648 ;
  assign n1735 = ( n1648 & n1725 ) | ( n1648 & n1733 ) | ( n1725 & n1733 ) ;
  assign n1736 = x88 & n888 ;
  assign n1737 = ( x90 & n878 ) | ( x90 & n1736 ) | ( n878 & n1736 ) ;
  assign n1738 = n1736 | n1737 ;
  assign n1739 = x89 & ~n877 ;
  assign n1740 = ( x89 & n1738 ) | ( x89 & ~n1739 ) | ( n1738 & ~n1739 ) ;
  assign n1741 = n1665 ^ x90 ^ x89 ;
  assign n1742 = n880 & n1741 ;
  assign n1743 = n1740 | n1742 ;
  assign n1744 = n1743 ^ x44 ^ 1'b0 ;
  assign n1745 = n1744 ^ n1690 ^ n1604 ;
  assign n1746 = ( n1604 & n1690 ) | ( n1604 & n1744 ) | ( n1690 & n1744 ) ;
  assign n1747 = x88 & n1058 ;
  assign n1748 = ( x90 & n1065 ) | ( x90 & n1747 ) | ( n1065 & n1747 ) ;
  assign n1749 = n1747 | n1748 ;
  assign n1750 = x89 & ~n1060 ;
  assign n1751 = ( x89 & n1749 ) | ( x89 & ~n1750 ) | ( n1749 & ~n1750 ) ;
  assign n1752 = ( x89 & x90 ) | ( x89 & n1665 ) | ( x90 & n1665 ) ;
  assign n1753 = n1063 & n1741 ;
  assign n1754 = n1751 | n1753 ;
  assign n1755 = n1754 ^ x41 ^ 1'b0 ;
  assign n1756 = ( n1488 & n1669 ) | ( n1488 & n1755 ) | ( n1669 & n1755 ) ;
  assign n1757 = n1755 ^ n1669 ^ n1488 ;
  assign n1758 = x83 & n561 ;
  assign n1759 = ( x85 & n551 ) | ( x85 & n1758 ) | ( n551 & n1758 ) ;
  assign n1760 = n1758 | n1759 ;
  assign n1761 = x84 & ~n550 ;
  assign n1762 = ( x84 & n1760 ) | ( x84 & ~n1761 ) | ( n1760 & ~n1761 ) ;
  assign n1763 = n553 & n1392 ;
  assign n1764 = n1762 | n1763 ;
  assign n1765 = n1764 ^ x50 ^ 1'b0 ;
  assign n1766 = ( n1679 & n1734 ) | ( n1679 & n1765 ) | ( n1734 & n1765 ) ;
  assign n1767 = n1765 ^ n1734 ^ n1679 ;
  assign n1768 = x86 & n744 ;
  assign n1769 = ( x88 & n730 ) | ( x88 & n1768 ) | ( n730 & n1768 ) ;
  assign n1770 = n1768 | n1769 ;
  assign n1771 = x87 & ~n732 ;
  assign n1772 = ( x87 & n1770 ) | ( x87 & ~n1771 ) | ( n1770 & ~n1771 ) ;
  assign n1773 = n731 & n1569 ;
  assign n1774 = n1772 | n1773 ;
  assign n1775 = n1774 ^ x47 ^ 1'b0 ;
  assign n1776 = ( n1689 & n1767 ) | ( n1689 & n1775 ) | ( n1767 & n1775 ) ;
  assign n1777 = n1775 ^ n1767 ^ n1689 ;
  assign n1778 = x72 & n208 ;
  assign n1779 = ( x74 & n194 ) | ( x74 & n1778 ) | ( n194 & n1778 ) ;
  assign n1780 = x71 & ~n242 ;
  assign n1781 = n1778 | n1779 ;
  assign n1782 = x70 & n325 ;
  assign n1783 = x73 & ~n192 ;
  assign n1784 = ( x73 & n1781 ) | ( x73 & ~n1783 ) | ( n1781 & ~n1783 ) ;
  assign n1785 = ( x71 & ~n1780 ) | ( x71 & n1782 ) | ( ~n1780 & n1782 ) ;
  assign n1786 = x75 & n133 ;
  assign n1787 = ( x77 & n142 ) | ( x77 & n1786 ) | ( n142 & n1786 ) ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = ( n197 & n504 ) | ( n197 & n1784 ) | ( n504 & n1784 ) ;
  assign n1790 = n1784 | n1789 ;
  assign n1791 = n1790 ^ x62 ^ 1'b0 ;
  assign n1792 = n1791 ^ n1785 ^ n1716 ;
  assign n1793 = ( n1716 & n1785 ) | ( n1716 & ~n1791 ) | ( n1785 & ~n1791 ) ;
  assign n1794 = x76 & ~n134 ;
  assign n1795 = ( x76 & n1788 ) | ( x76 & ~n1794 ) | ( n1788 & ~n1794 ) ;
  assign n1796 = n140 & n690 ;
  assign n1797 = n1795 | n1796 ;
  assign n1798 = n1797 ^ x59 ^ 1'b0 ;
  assign n1799 = ( n1703 & n1792 ) | ( n1703 & n1798 ) | ( n1792 & n1798 ) ;
  assign n1800 = n1798 ^ n1792 ^ n1703 ;
  assign n1801 = x78 & n263 ;
  assign n1802 = ( x80 & n264 ) | ( x80 & n1801 ) | ( n264 & n1801 ) ;
  assign n1803 = n1801 | n1802 ;
  assign n1804 = x79 & ~n260 ;
  assign n1805 = ( x79 & n1803 ) | ( x79 & ~n1804 ) | ( n1803 & ~n1804 ) ;
  assign n1806 = n272 & n1216 ;
  assign n1807 = n1805 | n1806 ;
  assign n1808 = n1807 ^ x56 ^ 1'b0 ;
  assign n1809 = n1808 ^ n1800 ^ n1713 ;
  assign n1810 = ( n1713 & n1800 ) | ( n1713 & n1808 ) | ( n1800 & n1808 ) ;
  assign n1811 = x81 & n408 ;
  assign n1812 = ( x83 & n403 ) | ( x83 & n1811 ) | ( n403 & n1811 ) ;
  assign n1813 = n1811 | n1812 ;
  assign n1814 = x82 & ~n410 ;
  assign n1815 = ( x82 & n1813 ) | ( x82 & ~n1814 ) | ( n1813 & ~n1814 ) ;
  assign n1816 = n402 & n1329 ;
  assign n1817 = n1815 | n1816 ;
  assign n1818 = n1817 ^ x53 ^ 1'b0 ;
  assign n1819 = n1818 ^ n1809 ^ n1724 ;
  assign n1820 = ( n1724 & n1809 ) | ( n1724 & n1818 ) | ( n1809 & n1818 ) ;
  assign n1821 = n731 & n1654 ;
  assign n1822 = x84 & n561 ;
  assign n1823 = ( x86 & n551 ) | ( x86 & n1822 ) | ( n551 & n1822 ) ;
  assign n1824 = n553 & n1419 ;
  assign n1825 = n1822 | n1823 ;
  assign n1826 = x85 & ~n550 ;
  assign n1827 = ( x85 & n1825 ) | ( x85 & ~n1826 ) | ( n1825 & ~n1826 ) ;
  assign n1828 = n1824 | n1827 ;
  assign n1829 = x72 & ~n242 ;
  assign n1830 = n1828 ^ x50 ^ 1'b0 ;
  assign n1831 = n1830 ^ n1819 ^ n1735 ;
  assign n1832 = ( n1735 & n1819 ) | ( n1735 & n1830 ) | ( n1819 & n1830 ) ;
  assign n1833 = x87 & n744 ;
  assign n1834 = ( x89 & n730 ) | ( x89 & n1833 ) | ( n730 & n1833 ) ;
  assign n1835 = n1833 | n1834 ;
  assign n1836 = x88 & ~n732 ;
  assign n1837 = ( x88 & n1835 ) | ( x88 & ~n1836 ) | ( n1835 & ~n1836 ) ;
  assign n1838 = n1821 | n1837 ;
  assign n1839 = n1838 ^ x47 ^ 1'b0 ;
  assign n1840 = x71 & n325 ;
  assign n1841 = ( x72 & ~n1829 ) | ( x72 & n1840 ) | ( ~n1829 & n1840 ) ;
  assign n1842 = x74 & n208 ;
  assign n1843 = ( x76 & n194 ) | ( x76 & n1842 ) | ( n194 & n1842 ) ;
  assign n1844 = n1842 | n1843 ;
  assign n1845 = x75 & ~n192 ;
  assign n1846 = ( x75 & n1844 ) | ( x75 & ~n1845 ) | ( n1844 & ~n1845 ) ;
  assign n1847 = n197 & n664 ;
  assign n1848 = n1846 | n1847 ;
  assign n1849 = n1848 ^ x62 ^ 1'b0 ;
  assign n1850 = ( ~n1785 & n1793 ) | ( ~n1785 & n1841 ) | ( n1793 & n1841 ) ;
  assign n1851 = n1841 ^ n1793 ^ n1785 ;
  assign n1852 = ( n1766 & n1831 ) | ( n1766 & n1839 ) | ( n1831 & n1839 ) ;
  assign n1853 = n1839 ^ n1831 ^ n1766 ;
  assign n1854 = x73 & ~n242 ;
  assign n1855 = x72 & n325 ;
  assign n1856 = ( x73 & ~n1854 ) | ( x73 & n1855 ) | ( ~n1854 & n1855 ) ;
  assign n1857 = n1856 ^ n1841 ^ x8 ;
  assign n1858 = ( ~x8 & n1841 ) | ( ~x8 & n1856 ) | ( n1841 & n1856 ) ;
  assign n1859 = n1857 ^ n1850 ^ n1849 ;
  assign n1860 = ( ~n1849 & n1850 ) | ( ~n1849 & n1857 ) | ( n1850 & n1857 ) ;
  assign n1861 = x76 & n133 ;
  assign n1862 = ( x78 & n142 ) | ( x78 & n1861 ) | ( n142 & n1861 ) ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = x77 & ~n134 ;
  assign n1865 = ( x77 & n1863 ) | ( x77 & ~n1864 ) | ( n1863 & ~n1864 ) ;
  assign n1866 = x73 & n208 ;
  assign n1867 = ( x75 & n194 ) | ( x75 & n1866 ) | ( n194 & n1866 ) ;
  assign n1868 = n1866 | n1867 ;
  assign n1869 = n140 & n709 ;
  assign n1870 = n1865 | n1869 ;
  assign n1871 = x74 & ~n192 ;
  assign n1872 = ( x74 & n1868 ) | ( x74 & ~n1871 ) | ( n1868 & ~n1871 ) ;
  assign n1873 = n197 & n525 ;
  assign n1874 = n1872 | n1873 ;
  assign n1875 = n1870 ^ x59 ^ 1'b0 ;
  assign n1876 = n1874 ^ x62 ^ 1'b0 ;
  assign n1877 = n1876 ^ n1875 ^ n1851 ;
  assign n1878 = ( n1851 & n1875 ) | ( n1851 & n1876 ) | ( n1875 & n1876 ) ;
  assign n1879 = x79 & n263 ;
  assign n1880 = ( x81 & n264 ) | ( x81 & n1879 ) | ( n264 & n1879 ) ;
  assign n1881 = n1879 | n1880 ;
  assign n1882 = x80 & ~n260 ;
  assign n1883 = ( x80 & n1881 ) | ( x80 & ~n1882 ) | ( n1881 & ~n1882 ) ;
  assign n1884 = n272 & n1258 ;
  assign n1885 = n1883 | n1884 ;
  assign n1886 = n1885 ^ x56 ^ 1'b0 ;
  assign n1887 = ( n1799 & n1877 ) | ( n1799 & n1886 ) | ( n1877 & n1886 ) ;
  assign n1888 = n1886 ^ n1877 ^ n1799 ;
  assign n1889 = x82 & n408 ;
  assign n1890 = ( x84 & n403 ) | ( x84 & n1889 ) | ( n403 & n1889 ) ;
  assign n1891 = n1889 | n1890 ;
  assign n1892 = x83 & ~n410 ;
  assign n1893 = ( x83 & n1891 ) | ( x83 & ~n1892 ) | ( n1891 & ~n1892 ) ;
  assign n1894 = n402 & n1355 ;
  assign n1895 = n1893 | n1894 ;
  assign n1896 = n1895 ^ x53 ^ 1'b0 ;
  assign n1897 = n1896 ^ n1888 ^ n1810 ;
  assign n1898 = ( n1810 & n1888 ) | ( n1810 & n1896 ) | ( n1888 & n1896 ) ;
  assign n1899 = x85 & n561 ;
  assign n1900 = ( x87 & n551 ) | ( x87 & n1899 ) | ( n551 & n1899 ) ;
  assign n1901 = n1899 | n1900 ;
  assign n1902 = x86 & ~n550 ;
  assign n1903 = ( x86 & n1901 ) | ( x86 & ~n1902 ) | ( n1901 & ~n1902 ) ;
  assign n1904 = n553 & n1484 ;
  assign n1905 = n1903 | n1904 ;
  assign n1906 = n1905 ^ x50 ^ 1'b0 ;
  assign n1907 = n1906 ^ n1897 ^ n1820 ;
  assign n1908 = ( n1820 & n1897 ) | ( n1820 & n1906 ) | ( n1897 & n1906 ) ;
  assign n1909 = x77 & n133 ;
  assign n1910 = ( x79 & n142 ) | ( x79 & n1909 ) | ( n142 & n1909 ) ;
  assign n1911 = n1909 | n1910 ;
  assign n1912 = x78 & ~n134 ;
  assign n1913 = ( x78 & n1911 ) | ( x78 & ~n1912 ) | ( n1911 & ~n1912 ) ;
  assign n1914 = n140 & n1015 ;
  assign n1915 = n1913 | n1914 ;
  assign n1916 = n1915 ^ x59 ^ 1'b0 ;
  assign n1917 = ( n1859 & n1878 ) | ( n1859 & n1916 ) | ( n1878 & n1916 ) ;
  assign n1918 = n1916 ^ n1878 ^ n1859 ;
  assign n1919 = x80 & n263 ;
  assign n1920 = ( x82 & n264 ) | ( x82 & n1919 ) | ( n264 & n1919 ) ;
  assign n1921 = n1919 | n1920 ;
  assign n1922 = x81 & ~n260 ;
  assign n1923 = ( x81 & n1921 ) | ( x81 & ~n1922 ) | ( n1921 & ~n1922 ) ;
  assign n1924 = n272 & n1301 ;
  assign n1925 = n1923 | n1924 ;
  assign n1926 = n1925 ^ x56 ^ 1'b0 ;
  assign n1927 = ( n1887 & n1918 ) | ( n1887 & n1926 ) | ( n1918 & n1926 ) ;
  assign n1928 = n1926 ^ n1918 ^ n1887 ;
  assign n1929 = x83 & n408 ;
  assign n1930 = ( x85 & n403 ) | ( x85 & n1929 ) | ( n403 & n1929 ) ;
  assign n1931 = n1929 | n1930 ;
  assign n1932 = x84 & ~n410 ;
  assign n1933 = ( x84 & n1931 ) | ( x84 & ~n1932 ) | ( n1931 & ~n1932 ) ;
  assign n1934 = n402 & n1392 ;
  assign n1935 = n1933 | n1934 ;
  assign n1936 = n1935 ^ x53 ^ 1'b0 ;
  assign n1937 = ( n1898 & n1928 ) | ( n1898 & n1936 ) | ( n1928 & n1936 ) ;
  assign n1938 = n1936 ^ n1928 ^ n1898 ;
  assign n1939 = x88 & n744 ;
  assign n1940 = ( x90 & n730 ) | ( x90 & n1939 ) | ( n730 & n1939 ) ;
  assign n1941 = n1939 | n1940 ;
  assign n1942 = x89 & ~n732 ;
  assign n1943 = ( x89 & n1941 ) | ( x89 & ~n1942 ) | ( n1941 & ~n1942 ) ;
  assign n1944 = n731 & n1741 ;
  assign n1945 = n1943 | n1944 ;
  assign n1946 = n1945 ^ x47 ^ 1'b0 ;
  assign n1947 = ( n1832 & n1907 ) | ( n1832 & n1946 ) | ( n1907 & n1946 ) ;
  assign n1948 = n1946 ^ n1907 ^ n1832 ;
  assign n1949 = x86 & n561 ;
  assign n1950 = ( x88 & n551 ) | ( x88 & n1949 ) | ( n551 & n1949 ) ;
  assign n1951 = n1949 | n1950 ;
  assign n1952 = x87 & ~n550 ;
  assign n1953 = ( x87 & n1951 ) | ( x87 & ~n1952 ) | ( n1951 & ~n1952 ) ;
  assign n1954 = n553 & n1569 ;
  assign n1955 = n1953 | n1954 ;
  assign n1956 = n1955 ^ x50 ^ 1'b0 ;
  assign n1957 = ( n1908 & n1938 ) | ( n1908 & n1956 ) | ( n1938 & n1956 ) ;
  assign n1958 = n1956 ^ n1938 ^ n1908 ;
  assign n1959 = x78 & n133 ;
  assign n1960 = x79 & ~n134 ;
  assign n1961 = n140 & n1216 ;
  assign n1962 = ( x80 & n142 ) | ( x80 & n1959 ) | ( n142 & n1959 ) ;
  assign n1963 = n1959 | n1962 ;
  assign n1964 = x73 & n325 ;
  assign n1965 = ( x79 & ~n1960 ) | ( x79 & n1963 ) | ( ~n1960 & n1963 ) ;
  assign n1966 = n1961 | n1965 ;
  assign n1967 = x74 & ~n242 ;
  assign n1968 = ( x74 & n1964 ) | ( x74 & ~n1967 ) | ( n1964 & ~n1967 ) ;
  assign n1969 = x75 & n208 ;
  assign n1970 = ( x77 & n194 ) | ( x77 & n1969 ) | ( n194 & n1969 ) ;
  assign n1971 = n1969 | n1970 ;
  assign n1972 = x76 & ~n192 ;
  assign n1973 = n1966 ^ x59 ^ 1'b0 ;
  assign n1974 = ( x76 & n1971 ) | ( x76 & ~n1972 ) | ( n1971 & ~n1972 ) ;
  assign n1975 = n197 & n690 ;
  assign n1976 = n1974 | n1975 ;
  assign n1977 = n1976 ^ x62 ^ 1'b0 ;
  assign n1978 = n1977 ^ n1968 ^ n1858 ;
  assign n1979 = ( n1858 & ~n1968 ) | ( n1858 & n1977 ) | ( ~n1968 & n1977 ) ;
  assign n1980 = ( n1860 & ~n1973 ) | ( n1860 & n1978 ) | ( ~n1973 & n1978 ) ;
  assign n1981 = n1978 ^ n1973 ^ n1860 ;
  assign n1982 = x81 & n263 ;
  assign n1983 = ( x83 & n264 ) | ( x83 & n1982 ) | ( n264 & n1982 ) ;
  assign n1984 = n1982 | n1983 ;
  assign n1985 = x82 & ~n260 ;
  assign n1986 = ( x82 & n1984 ) | ( x82 & ~n1985 ) | ( n1984 & ~n1985 ) ;
  assign n1987 = n272 & n1329 ;
  assign n1988 = n1986 | n1987 ;
  assign n1989 = n1988 ^ x56 ^ 1'b0 ;
  assign n1990 = n1989 ^ n1981 ^ n1917 ;
  assign n1991 = ( n1917 & n1981 ) | ( n1917 & n1989 ) | ( n1981 & n1989 ) ;
  assign n1992 = x84 & n408 ;
  assign n1993 = ( x86 & n403 ) | ( x86 & n1992 ) | ( n403 & n1992 ) ;
  assign n1994 = n1992 | n1993 ;
  assign n1995 = x85 & ~n410 ;
  assign n1996 = ( x85 & n1994 ) | ( x85 & ~n1995 ) | ( n1994 & ~n1995 ) ;
  assign n1997 = n402 & n1419 ;
  assign n1998 = n1996 | n1997 ;
  assign n1999 = n1998 ^ x53 ^ 1'b0 ;
  assign n2000 = n1999 ^ n1990 ^ n1927 ;
  assign n2001 = ( n1927 & n1990 ) | ( n1927 & n1999 ) | ( n1990 & n1999 ) ;
  assign n2002 = x87 & n561 ;
  assign n2003 = ( x89 & n551 ) | ( x89 & n2002 ) | ( n551 & n2002 ) ;
  assign n2004 = n2002 | n2003 ;
  assign n2005 = x88 & ~n550 ;
  assign n2006 = ( x88 & n2004 ) | ( x88 & ~n2005 ) | ( n2004 & ~n2005 ) ;
  assign n2007 = n553 & n1654 ;
  assign n2008 = n2006 | n2007 ;
  assign n2009 = n2008 ^ x50 ^ 1'b0 ;
  assign n2010 = n2009 ^ n2000 ^ n1937 ;
  assign n2011 = ( n1937 & n2000 ) | ( n1937 & n2009 ) | ( n2000 & n2009 ) ;
  assign n2012 = x74 & n325 ;
  assign n2013 = x79 & n133 ;
  assign n2014 = ( x81 & n142 ) | ( x81 & n2013 ) | ( n142 & n2013 ) ;
  assign n2015 = n2013 | n2014 ;
  assign n2016 = x80 & ~n134 ;
  assign n2017 = ( x80 & n2015 ) | ( x80 & ~n2016 ) | ( n2015 & ~n2016 ) ;
  assign n2018 = n140 & n1258 ;
  assign n2019 = x75 & ~n242 ;
  assign n2020 = ( x75 & n2012 ) | ( x75 & ~n2019 ) | ( n2012 & ~n2019 ) ;
  assign n2021 = ( ~n1968 & n1979 ) | ( ~n1968 & n2020 ) | ( n1979 & n2020 ) ;
  assign n2022 = n2017 | n2018 ;
  assign n2023 = n2020 ^ n1979 ^ n1968 ;
  assign n2024 = n2022 ^ x59 ^ 1'b0 ;
  assign n2025 = x76 & n208 ;
  assign n2026 = ( x78 & n194 ) | ( x78 & n2025 ) | ( n194 & n2025 ) ;
  assign n2027 = n2025 | n2026 ;
  assign n2028 = x77 & ~n192 ;
  assign n2029 = ( x77 & n2027 ) | ( x77 & ~n2028 ) | ( n2027 & ~n2028 ) ;
  assign n2030 = n197 & n709 ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = n2031 ^ x62 ^ 1'b0 ;
  assign n2033 = ( ~n2023 & n2024 ) | ( ~n2023 & n2032 ) | ( n2024 & n2032 ) ;
  assign n2034 = n2032 ^ n2024 ^ n2023 ;
  assign n2035 = x82 & n263 ;
  assign n2036 = ( x84 & n264 ) | ( x84 & n2035 ) | ( n264 & n2035 ) ;
  assign n2037 = n2035 | n2036 ;
  assign n2038 = x83 & ~n260 ;
  assign n2039 = ( x83 & n2037 ) | ( x83 & ~n2038 ) | ( n2037 & ~n2038 ) ;
  assign n2040 = n272 & n1355 ;
  assign n2041 = n2039 | n2040 ;
  assign n2042 = n2041 ^ x56 ^ 1'b0 ;
  assign n2043 = n2042 ^ n2034 ^ n1980 ;
  assign n2044 = ( n1980 & n2034 ) | ( n1980 & ~n2042 ) | ( n2034 & ~n2042 ) ;
  assign n2045 = x85 & n408 ;
  assign n2046 = ( x87 & n403 ) | ( x87 & n2045 ) | ( n403 & n2045 ) ;
  assign n2047 = n2045 | n2046 ;
  assign n2048 = x86 & ~n410 ;
  assign n2049 = ( x86 & n2047 ) | ( x86 & ~n2048 ) | ( n2047 & ~n2048 ) ;
  assign n2050 = n402 & n1484 ;
  assign n2051 = n2049 | n2050 ;
  assign n2052 = n2051 ^ x53 ^ 1'b0 ;
  assign n2053 = ( n1991 & n2043 ) | ( n1991 & n2052 ) | ( n2043 & n2052 ) ;
  assign n2054 = n2052 ^ n2043 ^ n1991 ;
  assign n2055 = x88 & n561 ;
  assign n2056 = ( x90 & n551 ) | ( x90 & n2055 ) | ( n551 & n2055 ) ;
  assign n2057 = n2055 | n2056 ;
  assign n2058 = x89 & ~n550 ;
  assign n2059 = ( x89 & n2057 ) | ( x89 & ~n2058 ) | ( n2057 & ~n2058 ) ;
  assign n2060 = n553 & n1741 ;
  assign n2061 = n2059 | n2060 ;
  assign n2062 = n2061 ^ x50 ^ 1'b0 ;
  assign n2063 = n2062 ^ n2054 ^ n2001 ;
  assign n2064 = ( n2001 & n2054 ) | ( n2001 & n2062 ) | ( n2054 & n2062 ) ;
  assign n2065 = x77 & n208 ;
  assign n2066 = ( x79 & n194 ) | ( x79 & n2065 ) | ( n194 & n2065 ) ;
  assign n2067 = n2065 | n2066 ;
  assign n2068 = x76 & ~n242 ;
  assign n2069 = x75 & n325 ;
  assign n2070 = ( x76 & ~n2068 ) | ( x76 & n2069 ) | ( ~n2068 & n2069 ) ;
  assign n2071 = x78 & ~n192 ;
  assign n2072 = ( x78 & n2067 ) | ( x78 & ~n2071 ) | ( n2067 & ~n2071 ) ;
  assign n2073 = n2070 ^ n1968 ^ x11 ;
  assign n2074 = ( ~x11 & n1968 ) | ( ~x11 & n2070 ) | ( n1968 & n2070 ) ;
  assign n2075 = n197 & n1015 ;
  assign n2076 = n2072 | n2075 ;
  assign n2077 = n2076 ^ x62 ^ 1'b0 ;
  assign n2078 = ( n2021 & ~n2073 ) | ( n2021 & n2077 ) | ( ~n2073 & n2077 ) ;
  assign n2079 = n2077 ^ n2073 ^ n2021 ;
  assign n2080 = x80 & n133 ;
  assign n2081 = ( x82 & n142 ) | ( x82 & n2080 ) | ( n142 & n2080 ) ;
  assign n2082 = n2080 | n2081 ;
  assign n2083 = x81 & ~n134 ;
  assign n2084 = ( x81 & n2082 ) | ( x81 & ~n2083 ) | ( n2082 & ~n2083 ) ;
  assign n2085 = n140 & n1301 ;
  assign n2086 = n2084 | n2085 ;
  assign n2087 = n2086 ^ x59 ^ 1'b0 ;
  assign n2088 = ( n2033 & ~n2079 ) | ( n2033 & n2087 ) | ( ~n2079 & n2087 ) ;
  assign n2089 = n2087 ^ n2079 ^ n2033 ;
  assign n2090 = x83 & n263 ;
  assign n2091 = ( x85 & n264 ) | ( x85 & n2090 ) | ( n264 & n2090 ) ;
  assign n2092 = n2090 | n2091 ;
  assign n2093 = x84 & ~n260 ;
  assign n2094 = ( x84 & n2092 ) | ( x84 & ~n2093 ) | ( n2092 & ~n2093 ) ;
  assign n2095 = n272 & n1392 ;
  assign n2096 = n2094 | n2095 ;
  assign n2097 = n2096 ^ x56 ^ 1'b0 ;
  assign n2098 = ( n2044 & n2089 ) | ( n2044 & ~n2097 ) | ( n2089 & ~n2097 ) ;
  assign n2099 = n2097 ^ n2089 ^ n2044 ;
  assign n2100 = x86 & n408 ;
  assign n2101 = ( x88 & n403 ) | ( x88 & n2100 ) | ( n403 & n2100 ) ;
  assign n2102 = n2100 | n2101 ;
  assign n2103 = x87 & ~n410 ;
  assign n2104 = ( x87 & n2102 ) | ( x87 & ~n2103 ) | ( n2102 & ~n2103 ) ;
  assign n2105 = n402 & n1569 ;
  assign n2106 = n2104 | n2105 ;
  assign n2107 = n2106 ^ x53 ^ 1'b0 ;
  assign n2108 = n2107 ^ n2099 ^ n2053 ;
  assign n2109 = ( n2053 & n2099 ) | ( n2053 & n2107 ) | ( n2099 & n2107 ) ;
  assign n2110 = x90 & ~n732 ;
  assign n2111 = x89 & n744 ;
  assign n2112 = ( x91 & n730 ) | ( x91 & n2111 ) | ( n730 & n2111 ) ;
  assign n2113 = n2111 | n2112 ;
  assign n2114 = n1752 ^ x91 ^ x90 ;
  assign n2115 = ( x90 & ~n2110 ) | ( x90 & n2113 ) | ( ~n2110 & n2113 ) ;
  assign n2116 = n731 & n2114 ;
  assign n2117 = n2115 | n2116 ;
  assign n2118 = n2117 ^ x47 ^ 1'b0 ;
  assign n2119 = ( n1947 & n1958 ) | ( n1947 & n2118 ) | ( n1958 & n2118 ) ;
  assign n2120 = n2118 ^ n1958 ^ n1947 ;
  assign n2121 = x89 & n561 ;
  assign n2122 = ( x91 & n551 ) | ( x91 & n2121 ) | ( n551 & n2121 ) ;
  assign n2123 = ( x90 & x91 ) | ( x90 & n1752 ) | ( x91 & n1752 ) ;
  assign n2124 = n2121 | n2122 ;
  assign n2125 = x90 & ~n550 ;
  assign n2126 = ( x90 & n2124 ) | ( x90 & ~n2125 ) | ( n2124 & ~n2125 ) ;
  assign n2127 = n553 & n2114 ;
  assign n2128 = n2126 | n2127 ;
  assign n2129 = n2128 ^ x50 ^ 1'b0 ;
  assign n2130 = ( n2064 & n2108 ) | ( n2064 & n2129 ) | ( n2108 & n2129 ) ;
  assign n2131 = n2129 ^ n2108 ^ n2064 ;
  assign n2132 = x89 & n1058 ;
  assign n2133 = ( x91 & n1065 ) | ( x91 & n2132 ) | ( n1065 & n2132 ) ;
  assign n2134 = n2132 | n2133 ;
  assign n2135 = x90 & ~n1060 ;
  assign n2136 = ( x90 & n2134 ) | ( x90 & ~n2135 ) | ( n2134 & ~n2135 ) ;
  assign n2137 = n1063 & n2114 ;
  assign n2138 = n2136 | n2137 ;
  assign n2139 = n2138 ^ x41 ^ 1'b0 ;
  assign n2140 = ( n1489 & n1573 ) | ( n1489 & n2139 ) | ( n1573 & n2139 ) ;
  assign n2141 = n2139 ^ n1573 ^ n1489 ;
  assign n2142 = x89 & n888 ;
  assign n2143 = ( x91 & n878 ) | ( x91 & n2142 ) | ( n878 & n2142 ) ;
  assign n2144 = n2142 | n2143 ;
  assign n2145 = x90 & ~n877 ;
  assign n2146 = ( x90 & n2144 ) | ( x90 & ~n2145 ) | ( n2144 & ~n2145 ) ;
  assign n2147 = n880 & n2114 ;
  assign n2148 = n2146 | n2147 ;
  assign n2149 = n2148 ^ x44 ^ 1'b0 ;
  assign n2150 = n2149 ^ n1777 ^ n1746 ;
  assign n2151 = ( n1746 & n1777 ) | ( n1746 & n2149 ) | ( n1777 & n2149 ) ;
  assign n2152 = x38 ^ x37 ^ 1'b0 ;
  assign n2153 = x36 ^ x35 ^ 1'b0 ;
  assign n2154 = x37 ^ x36 ^ 1'b0 ;
  assign n2155 = ( n2152 & ~n2153 ) | ( n2152 & n2154 ) | ( ~n2153 & n2154 ) ;
  assign n2156 = ~n2154 & n2155 ;
  assign n2157 = x64 & n2156 ;
  assign n2158 = ~n2153 & n2154 ;
  assign n2159 = x65 & ~n2158 ;
  assign n2160 = x64 & n2158 ;
  assign n2161 = n2152 & n2153 ;
  assign n2162 = ( n190 & n2160 ) | ( n190 & n2161 ) | ( n2160 & n2161 ) ;
  assign n2163 = ~n2152 & n2153 ;
  assign n2164 = ~x65 & n2163 ;
  assign n2165 = ( n2160 & n2163 ) | ( n2160 & ~n2164 ) | ( n2163 & ~n2164 ) ;
  assign n2166 = n2162 | n2165 ;
  assign n2167 = ( x66 & n2157 ) | ( x66 & n2163 ) | ( n2157 & n2163 ) ;
  assign n2168 = n139 & n2161 ;
  assign n2169 = n2157 | n2167 ;
  assign n2170 = ( x65 & ~n2159 ) | ( x65 & n2169 ) | ( ~n2159 & n2169 ) ;
  assign n2171 = x66 & ~n2158 ;
  assign n2172 = x65 & n2156 ;
  assign n2173 = n2168 | n2170 ;
  assign n2174 = ( x67 & n2163 ) | ( x67 & n2172 ) | ( n2163 & n2172 ) ;
  assign n2175 = n2172 | n2174 ;
  assign n2176 = n161 & n2161 ;
  assign n2177 = n2173 ^ x38 ^ 1'b0 ;
  assign n2178 = ( x66 & ~n2171 ) | ( x66 & n2175 ) | ( ~n2171 & n2175 ) ;
  assign n2179 = n2176 | n2178 ;
  assign n2180 = n2179 ^ x38 ^ 1'b0 ;
  assign n2181 = x64 & n2153 ;
  assign n2182 = n2166 ^ x38 ^ 1'b0 ;
  assign n2183 = x38 & ~n2181 ;
  assign n2184 = n2183 ^ n2182 ^ 1'b0 ;
  assign n2185 = n2182 & n2183 ;
  assign n2186 = n2185 ^ n2177 ^ 1'b0 ;
  assign n2187 = n2177 & n2185 ;
  assign n2188 = n2187 ^ n2180 ^ n1083 ;
  assign n2189 = ( n1083 & n2180 ) | ( n1083 & n2187 ) | ( n2180 & n2187 ) ;
  assign n2190 = x66 & n2156 ;
  assign n2191 = ( x68 & n2163 ) | ( x68 & n2190 ) | ( n2163 & n2190 ) ;
  assign n2192 = n2190 | n2191 ;
  assign n2193 = x67 & ~n2158 ;
  assign n2194 = ( x67 & n2192 ) | ( x67 & ~n2193 ) | ( n2192 & ~n2193 ) ;
  assign n2195 = n175 & n2161 ;
  assign n2196 = n2194 | n2195 ;
  assign n2197 = n2196 ^ x38 ^ 1'b0 ;
  assign n2198 = n2197 ^ n2189 ^ n1086 ;
  assign n2199 = ( n1086 & n2189 ) | ( n1086 & n2197 ) | ( n2189 & n2197 ) ;
  assign n2200 = x67 & n2156 ;
  assign n2201 = ( x69 & n2163 ) | ( x69 & n2200 ) | ( n2163 & n2200 ) ;
  assign n2202 = n2200 | n2201 ;
  assign n2203 = x68 & ~n2158 ;
  assign n2204 = ( x68 & n2202 ) | ( x68 & ~n2203 ) | ( n2202 & ~n2203 ) ;
  assign n2205 = n172 & n2161 ;
  assign n2206 = n2204 | n2205 ;
  assign n2207 = n2206 ^ x38 ^ 1'b0 ;
  assign n2208 = ( n1088 & n2199 ) | ( n1088 & n2207 ) | ( n2199 & n2207 ) ;
  assign n2209 = n2207 ^ n2199 ^ n1088 ;
  assign n2210 = x68 & n2156 ;
  assign n2211 = ( x70 & n2163 ) | ( x70 & n2210 ) | ( n2163 & n2210 ) ;
  assign n2212 = n2210 | n2211 ;
  assign n2213 = x69 & ~n2158 ;
  assign n2214 = ( x69 & n2212 ) | ( x69 & ~n2213 ) | ( n2212 & ~n2213 ) ;
  assign n2215 = n168 & n2161 ;
  assign n2216 = n2214 | n2215 ;
  assign n2217 = n2216 ^ x38 ^ 1'b0 ;
  assign n2218 = ( n1090 & n2208 ) | ( n1090 & n2217 ) | ( n2208 & n2217 ) ;
  assign n2219 = n2217 ^ n2208 ^ n1090 ;
  assign n2220 = x69 & n2156 ;
  assign n2221 = ( x71 & n2163 ) | ( x71 & n2220 ) | ( n2163 & n2220 ) ;
  assign n2222 = n2220 | n2221 ;
  assign n2223 = x70 & ~n2158 ;
  assign n2224 = ( x70 & n2222 ) | ( x70 & ~n2223 ) | ( n2222 & ~n2223 ) ;
  assign n2225 = n328 & n2161 ;
  assign n2226 = n2224 | n2225 ;
  assign n2227 = n2226 ^ x38 ^ 1'b0 ;
  assign n2228 = n2227 ^ n2218 ^ n1100 ;
  assign n2229 = ( n1100 & n2218 ) | ( n1100 & n2227 ) | ( n2218 & n2227 ) ;
  assign n2230 = x70 & n2156 ;
  assign n2231 = ( x72 & n2163 ) | ( x72 & n2230 ) | ( n2163 & n2230 ) ;
  assign n2232 = n2230 | n2231 ;
  assign n2233 = x71 & ~n2158 ;
  assign n2234 = ( x71 & n2232 ) | ( x71 & ~n2233 ) | ( n2232 & ~n2233 ) ;
  assign n2235 = n349 & n2161 ;
  assign n2236 = n2234 | n2235 ;
  assign n2237 = n2236 ^ x38 ^ 1'b0 ;
  assign n2238 = ( n1111 & n2229 ) | ( n1111 & n2237 ) | ( n2229 & n2237 ) ;
  assign n2239 = n2237 ^ n2229 ^ n1111 ;
  assign n2240 = x71 & n2156 ;
  assign n2241 = ( x73 & n2163 ) | ( x73 & n2240 ) | ( n2163 & n2240 ) ;
  assign n2242 = n2240 | n2241 ;
  assign n2243 = x72 & ~n2158 ;
  assign n2244 = ( x72 & n2242 ) | ( x72 & ~n2243 ) | ( n2242 & ~n2243 ) ;
  assign n2245 = n370 & n2161 ;
  assign n2246 = n2244 | n2245 ;
  assign n2247 = n2246 ^ x38 ^ 1'b0 ;
  assign n2248 = ( n1121 & n2238 ) | ( n1121 & n2247 ) | ( n2238 & n2247 ) ;
  assign n2249 = n2247 ^ n2238 ^ n1121 ;
  assign n2250 = x72 & n2156 ;
  assign n2251 = ( x74 & n2163 ) | ( x74 & n2250 ) | ( n2163 & n2250 ) ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = x73 & ~n2158 ;
  assign n2254 = ( x73 & n2252 ) | ( x73 & ~n2253 ) | ( n2252 & ~n2253 ) ;
  assign n2255 = n504 & n2161 ;
  assign n2256 = n2254 | n2255 ;
  assign n2257 = n2256 ^ x38 ^ 1'b0 ;
  assign n2258 = n2257 ^ n2248 ^ n1130 ;
  assign n2259 = ( n1130 & n2248 ) | ( n1130 & n2257 ) | ( n2248 & n2257 ) ;
  assign n2260 = x73 & n2156 ;
  assign n2261 = ( x75 & n2163 ) | ( x75 & n2260 ) | ( n2163 & n2260 ) ;
  assign n2262 = n2260 | n2261 ;
  assign n2263 = x74 & ~n2158 ;
  assign n2264 = ( x74 & n2262 ) | ( x74 & ~n2263 ) | ( n2262 & ~n2263 ) ;
  assign n2265 = n525 & n2161 ;
  assign n2266 = n2264 | n2265 ;
  assign n2267 = n2266 ^ x38 ^ 1'b0 ;
  assign n2268 = ( n1141 & n2259 ) | ( n1141 & n2267 ) | ( n2259 & n2267 ) ;
  assign n2269 = n2267 ^ n2259 ^ n1141 ;
  assign n2270 = x74 & n2156 ;
  assign n2271 = ( x76 & n2163 ) | ( x76 & n2270 ) | ( n2163 & n2270 ) ;
  assign n2272 = n2270 | n2271 ;
  assign n2273 = x75 & ~n2158 ;
  assign n2274 = ( x75 & n2272 ) | ( x75 & ~n2273 ) | ( n2272 & ~n2273 ) ;
  assign n2275 = n664 & n2161 ;
  assign n2276 = n2274 | n2275 ;
  assign n2277 = n2276 ^ x38 ^ 1'b0 ;
  assign n2278 = ( n1151 & n2268 ) | ( n1151 & n2277 ) | ( n2268 & n2277 ) ;
  assign n2279 = n2277 ^ n2268 ^ n1151 ;
  assign n2280 = x75 & n2156 ;
  assign n2281 = ( x77 & n2163 ) | ( x77 & n2280 ) | ( n2163 & n2280 ) ;
  assign n2282 = n2280 | n2281 ;
  assign n2283 = x76 & ~n2158 ;
  assign n2284 = ( x76 & n2282 ) | ( x76 & ~n2283 ) | ( n2282 & ~n2283 ) ;
  assign n2285 = n690 & n2161 ;
  assign n2286 = n2284 | n2285 ;
  assign n2287 = n2286 ^ x38 ^ 1'b0 ;
  assign n2288 = n2287 ^ n2278 ^ n1160 ;
  assign n2289 = ( n1160 & n2278 ) | ( n1160 & n2287 ) | ( n2278 & n2287 ) ;
  assign n2290 = x76 & n2156 ;
  assign n2291 = ( x78 & n2163 ) | ( x78 & n2290 ) | ( n2163 & n2290 ) ;
  assign n2292 = n2290 | n2291 ;
  assign n2293 = x77 & ~n2158 ;
  assign n2294 = ( x77 & n2292 ) | ( x77 & ~n2293 ) | ( n2292 & ~n2293 ) ;
  assign n2295 = n709 & n2161 ;
  assign n2296 = n2294 | n2295 ;
  assign n2297 = n2296 ^ x38 ^ 1'b0 ;
  assign n2298 = n2297 ^ n2289 ^ n1170 ;
  assign n2299 = ( n1170 & n2289 ) | ( n1170 & n2297 ) | ( n2289 & n2297 ) ;
  assign n2300 = x77 & n2156 ;
  assign n2301 = ( x79 & n2163 ) | ( x79 & n2300 ) | ( n2163 & n2300 ) ;
  assign n2302 = n2300 | n2301 ;
  assign n2303 = x78 & ~n2158 ;
  assign n2304 = ( x78 & n2302 ) | ( x78 & ~n2303 ) | ( n2302 & ~n2303 ) ;
  assign n2305 = n1015 & n2161 ;
  assign n2306 = n2304 | n2305 ;
  assign n2307 = n2306 ^ x38 ^ 1'b0 ;
  assign n2308 = ( n1180 & n2299 ) | ( n1180 & n2307 ) | ( n2299 & n2307 ) ;
  assign n2309 = n2307 ^ n2299 ^ n1180 ;
  assign n2310 = x78 & n2156 ;
  assign n2311 = ( x80 & n2163 ) | ( x80 & n2310 ) | ( n2163 & n2310 ) ;
  assign n2312 = n2310 | n2311 ;
  assign n2313 = x79 & ~n2158 ;
  assign n2314 = ( x79 & n2312 ) | ( x79 & ~n2313 ) | ( n2312 & ~n2313 ) ;
  assign n2315 = n1216 & n2161 ;
  assign n2316 = n2314 | n2315 ;
  assign n2317 = n2316 ^ x38 ^ 1'b0 ;
  assign n2318 = ( n1190 & n2308 ) | ( n1190 & n2317 ) | ( n2308 & n2317 ) ;
  assign n2319 = n2317 ^ n2308 ^ n1190 ;
  assign n2320 = x79 & n2156 ;
  assign n2321 = ( x81 & n2163 ) | ( x81 & n2320 ) | ( n2163 & n2320 ) ;
  assign n2322 = n2320 | n2321 ;
  assign n2323 = x80 & ~n2158 ;
  assign n2324 = ( x80 & n2322 ) | ( x80 & ~n2323 ) | ( n2322 & ~n2323 ) ;
  assign n2325 = n1258 & n2161 ;
  assign n2326 = n2324 | n2325 ;
  assign n2327 = n2326 ^ x38 ^ 1'b0 ;
  assign n2328 = n2327 ^ n2318 ^ n1201 ;
  assign n2329 = ( n1201 & n2318 ) | ( n1201 & n2327 ) | ( n2318 & n2327 ) ;
  assign n2330 = x80 & n2156 ;
  assign n2331 = ( x82 & n2163 ) | ( x82 & n2330 ) | ( n2163 & n2330 ) ;
  assign n2332 = n2330 | n2331 ;
  assign n2333 = x81 & ~n2158 ;
  assign n2334 = ( x81 & n2332 ) | ( x81 & ~n2333 ) | ( n2332 & ~n2333 ) ;
  assign n2335 = n1301 & n2161 ;
  assign n2336 = n2334 | n2335 ;
  assign n2337 = n2336 ^ x38 ^ 1'b0 ;
  assign n2338 = ( n1211 & n2329 ) | ( n1211 & n2337 ) | ( n2329 & n2337 ) ;
  assign n2339 = n2337 ^ n2329 ^ n1211 ;
  assign n2340 = x81 & n2156 ;
  assign n2341 = ( x83 & n2163 ) | ( x83 & n2340 ) | ( n2163 & n2340 ) ;
  assign n2342 = n2340 | n2341 ;
  assign n2343 = x82 & ~n2158 ;
  assign n2344 = ( x82 & n2342 ) | ( x82 & ~n2343 ) | ( n2342 & ~n2343 ) ;
  assign n2345 = n1329 & n2161 ;
  assign n2346 = n2344 | n2345 ;
  assign n2347 = n2346 ^ x38 ^ 1'b0 ;
  assign n2348 = n2347 ^ n2338 ^ n1243 ;
  assign n2349 = ( n1243 & n2338 ) | ( n1243 & n2347 ) | ( n2338 & n2347 ) ;
  assign n2350 = x82 & n2156 ;
  assign n2351 = ( x84 & n2163 ) | ( x84 & n2350 ) | ( n2163 & n2350 ) ;
  assign n2352 = n2350 | n2351 ;
  assign n2353 = x83 & ~n2158 ;
  assign n2354 = ( x83 & n2352 ) | ( x83 & ~n2353 ) | ( n2352 & ~n2353 ) ;
  assign n2355 = n1355 & n2161 ;
  assign n2356 = n2354 | n2355 ;
  assign n2357 = n2356 ^ x38 ^ 1'b0 ;
  assign n2358 = ( n1285 & n2349 ) | ( n1285 & n2357 ) | ( n2349 & n2357 ) ;
  assign n2359 = n2357 ^ n2349 ^ n1285 ;
  assign n2360 = x83 & n2156 ;
  assign n2361 = ( x85 & n2163 ) | ( x85 & n2360 ) | ( n2163 & n2360 ) ;
  assign n2362 = n2360 | n2361 ;
  assign n2363 = x84 & ~n2158 ;
  assign n2364 = ( x84 & n2362 ) | ( x84 & ~n2363 ) | ( n2362 & ~n2363 ) ;
  assign n2365 = n1392 & n2161 ;
  assign n2366 = n2364 | n2365 ;
  assign n2367 = n2366 ^ x38 ^ 1'b0 ;
  assign n2368 = ( n1308 & n2358 ) | ( n1308 & n2367 ) | ( n2358 & n2367 ) ;
  assign n2369 = n2367 ^ n2358 ^ n1308 ;
  assign n2370 = x84 & n2156 ;
  assign n2371 = ( x86 & n2163 ) | ( x86 & n2370 ) | ( n2163 & n2370 ) ;
  assign n2372 = n2370 | n2371 ;
  assign n2373 = x85 & ~n2158 ;
  assign n2374 = ( x85 & n2372 ) | ( x85 & ~n2373 ) | ( n2372 & ~n2373 ) ;
  assign n2375 = n1419 & n2161 ;
  assign n2376 = n2374 | n2375 ;
  assign n2377 = n2376 ^ x38 ^ 1'b0 ;
  assign n2378 = ( n1381 & n2368 ) | ( n1381 & n2377 ) | ( n2368 & n2377 ) ;
  assign n2379 = n2377 ^ n2368 ^ n1381 ;
  assign n2380 = x85 & n2156 ;
  assign n2381 = ( x87 & n2163 ) | ( x87 & n2380 ) | ( n2163 & n2380 ) ;
  assign n2382 = n2380 | n2381 ;
  assign n2383 = x86 & ~n2158 ;
  assign n2384 = ( x86 & n2382 ) | ( x86 & ~n2383 ) | ( n2382 & ~n2383 ) ;
  assign n2385 = n1484 & n2161 ;
  assign n2386 = n2384 | n2385 ;
  assign n2387 = n2386 ^ x38 ^ 1'b0 ;
  assign n2388 = n2387 ^ n2378 ^ n1390 ;
  assign n2389 = ( n1390 & n2378 ) | ( n1390 & n2387 ) | ( n2378 & n2387 ) ;
  assign n2390 = x86 & n2156 ;
  assign n2391 = ( x88 & n2163 ) | ( x88 & n2390 ) | ( n2163 & n2390 ) ;
  assign n2392 = n2390 | n2391 ;
  assign n2393 = x87 & ~n2158 ;
  assign n2394 = ( x87 & n2392 ) | ( x87 & ~n2393 ) | ( n2392 & ~n2393 ) ;
  assign n2395 = n1569 & n2161 ;
  assign n2396 = n2394 | n2395 ;
  assign n2397 = n2396 ^ x38 ^ 1'b0 ;
  assign n2398 = ( n1415 & n2389 ) | ( n1415 & n2397 ) | ( n2389 & n2397 ) ;
  assign n2399 = n2397 ^ n2389 ^ n1415 ;
  assign n2400 = x87 & n2156 ;
  assign n2401 = ( x89 & n2163 ) | ( x89 & n2400 ) | ( n2163 & n2400 ) ;
  assign n2402 = n2400 | n2401 ;
  assign n2403 = x88 & ~n2158 ;
  assign n2404 = ( x88 & n2402 ) | ( x88 & ~n2403 ) | ( n2402 & ~n2403 ) ;
  assign n2405 = n1654 & n2161 ;
  assign n2406 = n2404 | n2405 ;
  assign n2407 = n2406 ^ x38 ^ 1'b0 ;
  assign n2408 = ( n1434 & n2398 ) | ( n1434 & n2407 ) | ( n2398 & n2407 ) ;
  assign n2409 = n2407 ^ n2398 ^ n1434 ;
  assign n2410 = x88 & n2156 ;
  assign n2411 = ( x90 & n2163 ) | ( x90 & n2410 ) | ( n2163 & n2410 ) ;
  assign n2412 = n2410 | n2411 ;
  assign n2413 = x89 & ~n2158 ;
  assign n2414 = ( x89 & n2412 ) | ( x89 & ~n2413 ) | ( n2412 & ~n2413 ) ;
  assign n2415 = n1741 & n2161 ;
  assign n2416 = n2414 | n2415 ;
  assign n2417 = n2416 ^ x38 ^ 1'b0 ;
  assign n2418 = ( n1500 & n2408 ) | ( n1500 & n2417 ) | ( n2408 & n2417 ) ;
  assign n2419 = n2417 ^ n2408 ^ n1500 ;
  assign n2420 = n2123 ^ x92 ^ x91 ;
  assign n2421 = x90 & n888 ;
  assign n2422 = ( x92 & n878 ) | ( x92 & n2421 ) | ( n878 & n2421 ) ;
  assign n2423 = n2421 | n2422 ;
  assign n2424 = x91 & ~n877 ;
  assign n2425 = ( x91 & n2423 ) | ( x91 & ~n2424 ) | ( n2423 & ~n2424 ) ;
  assign n2426 = n880 & n2420 ;
  assign n2427 = n2425 | n2426 ;
  assign n2428 = n2427 ^ x44 ^ 1'b0 ;
  assign n2429 = n2428 ^ n1853 ^ n1776 ;
  assign n2430 = ( n1776 & n1853 ) | ( n1776 & n2428 ) | ( n1853 & n2428 ) ;
  assign n2431 = ( x91 & x92 ) | ( x91 & n2123 ) | ( x92 & n2123 ) ;
  assign n2432 = x90 & n1058 ;
  assign n2433 = ( x92 & n1065 ) | ( x92 & n2432 ) | ( n1065 & n2432 ) ;
  assign n2434 = n2432 | n2433 ;
  assign n2435 = x91 & ~n1060 ;
  assign n2436 = ( x91 & n2434 ) | ( x91 & ~n2435 ) | ( n2434 & ~n2435 ) ;
  assign n2437 = n1063 & n2420 ;
  assign n2438 = n2436 | n2437 ;
  assign n2439 = n2438 ^ x41 ^ 1'b0 ;
  assign n2440 = ( n1574 & n1658 ) | ( n1574 & n2439 ) | ( n1658 & n2439 ) ;
  assign n2441 = n2439 ^ n1658 ^ n1574 ;
  assign n2442 = x89 & n2156 ;
  assign n2443 = ( x91 & n2163 ) | ( x91 & n2442 ) | ( n2163 & n2442 ) ;
  assign n2444 = n2442 | n2443 ;
  assign n2445 = x90 & ~n2158 ;
  assign n2446 = ( x90 & n2444 ) | ( x90 & ~n2445 ) | ( n2444 & ~n2445 ) ;
  assign n2447 = n2114 & n2161 ;
  assign n2448 = n2446 | n2447 ;
  assign n2449 = n2448 ^ x38 ^ 1'b0 ;
  assign n2450 = ( n1585 & n2418 ) | ( n1585 & n2449 ) | ( n2418 & n2449 ) ;
  assign n2451 = n2449 ^ n2418 ^ n1585 ;
  assign n2452 = x90 & n744 ;
  assign n2453 = ( x92 & n730 ) | ( x92 & n2452 ) | ( n730 & n2452 ) ;
  assign n2454 = n2452 | n2453 ;
  assign n2455 = x91 & ~n732 ;
  assign n2456 = ( x91 & n2454 ) | ( x91 & ~n2455 ) | ( n2454 & ~n2455 ) ;
  assign n2457 = n731 & n2420 ;
  assign n2458 = n2456 | n2457 ;
  assign n2459 = n2458 ^ x47 ^ 1'b0 ;
  assign n2460 = n2459 ^ n2010 ^ n1957 ;
  assign n2461 = ( n1957 & n2010 ) | ( n1957 & n2459 ) | ( n2010 & n2459 ) ;
  assign n2462 = x90 & n2156 ;
  assign n2463 = ( x92 & n2163 ) | ( x92 & n2462 ) | ( n2163 & n2462 ) ;
  assign n2464 = n2462 | n2463 ;
  assign n2465 = x91 & ~n2158 ;
  assign n2466 = ( x91 & n2464 ) | ( x91 & ~n2465 ) | ( n2464 & ~n2465 ) ;
  assign n2467 = n2161 & n2420 ;
  assign n2468 = n2466 | n2467 ;
  assign n2469 = n2468 ^ x38 ^ 1'b0 ;
  assign n2470 = ( n1670 & n2450 ) | ( n1670 & n2469 ) | ( n2450 & n2469 ) ;
  assign n2471 = n2469 ^ n2450 ^ n1670 ;
  assign n2472 = x92 & ~n877 ;
  assign n2473 = x91 & n888 ;
  assign n2474 = ( x93 & n878 ) | ( x93 & n2473 ) | ( n878 & n2473 ) ;
  assign n2475 = n2473 | n2474 ;
  assign n2476 = n2431 ^ x93 ^ x92 ;
  assign n2477 = ( x92 & ~n2472 ) | ( x92 & n2475 ) | ( ~n2472 & n2475 ) ;
  assign n2478 = n880 & n2476 ;
  assign n2479 = n2477 | n2478 ;
  assign n2480 = n2479 ^ x44 ^ 1'b0 ;
  assign n2481 = ( n1852 & n1948 ) | ( n1852 & n2480 ) | ( n1948 & n2480 ) ;
  assign n2482 = n2480 ^ n1948 ^ n1852 ;
  assign n2483 = x91 & n744 ;
  assign n2484 = ( x93 & n730 ) | ( x93 & n2483 ) | ( n730 & n2483 ) ;
  assign n2485 = ( x92 & x93 ) | ( x92 & n2431 ) | ( x93 & n2431 ) ;
  assign n2486 = n2483 | n2484 ;
  assign n2487 = x92 & ~n732 ;
  assign n2488 = ( x92 & n2486 ) | ( x92 & ~n2487 ) | ( n2486 & ~n2487 ) ;
  assign n2489 = n731 & n2476 ;
  assign n2490 = n2488 | n2489 ;
  assign n2491 = n2490 ^ x47 ^ 1'b0 ;
  assign n2492 = ( n2011 & n2063 ) | ( n2011 & n2491 ) | ( n2063 & n2491 ) ;
  assign n2493 = n2491 ^ n2063 ^ n2011 ;
  assign n2494 = x91 & n2156 ;
  assign n2495 = ( x93 & n2163 ) | ( x93 & n2494 ) | ( n2163 & n2494 ) ;
  assign n2496 = n2494 | n2495 ;
  assign n2497 = x92 & ~n2158 ;
  assign n2498 = ( x92 & n2496 ) | ( x92 & ~n2497 ) | ( n2496 & ~n2497 ) ;
  assign n2499 = n2161 & n2476 ;
  assign n2500 = n2498 | n2499 ;
  assign n2501 = n2500 ^ x38 ^ 1'b0 ;
  assign n2502 = ( n1757 & n2470 ) | ( n1757 & n2501 ) | ( n2470 & n2501 ) ;
  assign n2503 = n2501 ^ n2470 ^ n1757 ;
  assign n2504 = x91 & n1058 ;
  assign n2505 = ( x93 & n1065 ) | ( x93 & n2504 ) | ( n1065 & n2504 ) ;
  assign n2506 = n2504 | n2505 ;
  assign n2507 = x92 & ~n1060 ;
  assign n2508 = ( x92 & n2506 ) | ( x92 & ~n2507 ) | ( n2506 & ~n2507 ) ;
  assign n2509 = n1063 & n2476 ;
  assign n2510 = n2508 | n2509 ;
  assign n2511 = n2510 ^ x41 ^ 1'b0 ;
  assign n2512 = n2511 ^ n1745 ^ n1659 ;
  assign n2513 = ( n1659 & n1745 ) | ( n1659 & n2511 ) | ( n1745 & n2511 ) ;
  assign n2514 = x93 & ~n877 ;
  assign n2515 = x92 & n888 ;
  assign n2516 = ( x94 & n878 ) | ( x94 & n2515 ) | ( n878 & n2515 ) ;
  assign n2517 = n2515 | n2516 ;
  assign n2518 = n2485 ^ x94 ^ x93 ;
  assign n2519 = ( x93 & ~n2514 ) | ( x93 & n2517 ) | ( ~n2514 & n2517 ) ;
  assign n2520 = n880 & n2518 ;
  assign n2521 = n2519 | n2520 ;
  assign n2522 = n2521 ^ x44 ^ 1'b0 ;
  assign n2523 = ( n2120 & n2481 ) | ( n2120 & n2522 ) | ( n2481 & n2522 ) ;
  assign n2524 = n2522 ^ n2481 ^ n2120 ;
  assign n2525 = x92 & n744 ;
  assign n2526 = ( x94 & n730 ) | ( x94 & n2525 ) | ( n730 & n2525 ) ;
  assign n2527 = ( x93 & x94 ) | ( x93 & n2485 ) | ( x94 & n2485 ) ;
  assign n2528 = n2525 | n2526 ;
  assign n2529 = x93 & ~n732 ;
  assign n2530 = ( x93 & n2528 ) | ( x93 & ~n2529 ) | ( n2528 & ~n2529 ) ;
  assign n2531 = n731 & n2518 ;
  assign n2532 = n2530 | n2531 ;
  assign n2533 = n2532 ^ x47 ^ 1'b0 ;
  assign n2534 = ( n2131 & n2492 ) | ( n2131 & n2533 ) | ( n2492 & n2533 ) ;
  assign n2535 = n2533 ^ n2492 ^ n2131 ;
  assign n2536 = x92 & n2156 ;
  assign n2537 = ( x94 & n2163 ) | ( x94 & n2536 ) | ( n2163 & n2536 ) ;
  assign n2538 = n2536 | n2537 ;
  assign n2539 = x93 & ~n2158 ;
  assign n2540 = ( x93 & n2538 ) | ( x93 & ~n2539 ) | ( n2538 & ~n2539 ) ;
  assign n2541 = n2161 & n2518 ;
  assign n2542 = n2540 | n2541 ;
  assign n2543 = n2542 ^ x38 ^ 1'b0 ;
  assign n2544 = ( n1756 & n2141 ) | ( n1756 & n2543 ) | ( n2141 & n2543 ) ;
  assign n2545 = n2543 ^ n2141 ^ n1756 ;
  assign n2546 = x92 & n1058 ;
  assign n2547 = ( x94 & n1065 ) | ( x94 & n2546 ) | ( n1065 & n2546 ) ;
  assign n2548 = n2546 | n2547 ;
  assign n2549 = x93 & ~n1060 ;
  assign n2550 = ( x93 & n2548 ) | ( x93 & ~n2549 ) | ( n2548 & ~n2549 ) ;
  assign n2551 = n1063 & n2518 ;
  assign n2552 = n2550 | n2551 ;
  assign n2553 = n2552 ^ x41 ^ 1'b0 ;
  assign n2554 = n2553 ^ n2513 ^ n2150 ;
  assign n2555 = ( n2150 & n2513 ) | ( n2150 & n2553 ) | ( n2513 & n2553 ) ;
  assign n2556 = x35 ^ x34 ^ 1'b0 ;
  assign n2557 = x33 ^ x32 ^ 1'b0 ;
  assign n2558 = x34 ^ x33 ^ 1'b0 ;
  assign n2559 = ( n2556 & ~n2557 ) | ( n2556 & n2558 ) | ( ~n2557 & n2558 ) ;
  assign n2560 = ~n2558 & n2559 ;
  assign n2561 = x64 & n2560 ;
  assign n2562 = ~n2557 & n2558 ;
  assign n2563 = x65 & ~n2562 ;
  assign n2564 = x64 & n2562 ;
  assign n2565 = n2556 & n2557 ;
  assign n2566 = ( n190 & n2564 ) | ( n190 & n2565 ) | ( n2564 & n2565 ) ;
  assign n2567 = ~n2556 & n2557 ;
  assign n2568 = ~x65 & n2567 ;
  assign n2569 = ( n2564 & n2567 ) | ( n2564 & ~n2568 ) | ( n2567 & ~n2568 ) ;
  assign n2570 = n2566 | n2569 ;
  assign n2571 = ( x66 & n2561 ) | ( x66 & n2567 ) | ( n2561 & n2567 ) ;
  assign n2572 = n139 & n2565 ;
  assign n2573 = n2561 | n2571 ;
  assign n2574 = ( x65 & ~n2563 ) | ( x65 & n2573 ) | ( ~n2563 & n2573 ) ;
  assign n2575 = x66 & ~n2562 ;
  assign n2576 = x65 & n2560 ;
  assign n2577 = n2572 | n2574 ;
  assign n2578 = ( x67 & n2567 ) | ( x67 & n2576 ) | ( n2567 & n2576 ) ;
  assign n2579 = n2576 | n2578 ;
  assign n2580 = n161 & n2565 ;
  assign n2581 = n2577 ^ x35 ^ 1'b0 ;
  assign n2582 = ( x66 & ~n2575 ) | ( x66 & n2579 ) | ( ~n2575 & n2579 ) ;
  assign n2583 = n2580 | n2582 ;
  assign n2584 = n2583 ^ x35 ^ 1'b0 ;
  assign n2585 = x64 & n2557 ;
  assign n2586 = n2570 ^ x35 ^ 1'b0 ;
  assign n2587 = x35 & ~n2585 ;
  assign n2588 = n2587 ^ n2586 ^ 1'b0 ;
  assign n2589 = n2586 & n2587 ;
  assign n2590 = n2589 ^ n2581 ^ 1'b0 ;
  assign n2591 = n2581 & n2589 ;
  assign n2592 = n2591 ^ n2584 ^ n2181 ;
  assign n2593 = ( n2181 & n2584 ) | ( n2181 & n2591 ) | ( n2584 & n2591 ) ;
  assign n2594 = x66 & n2560 ;
  assign n2595 = ( x68 & n2567 ) | ( x68 & n2594 ) | ( n2567 & n2594 ) ;
  assign n2596 = n2594 | n2595 ;
  assign n2597 = x67 & ~n2562 ;
  assign n2598 = ( x67 & n2596 ) | ( x67 & ~n2597 ) | ( n2596 & ~n2597 ) ;
  assign n2599 = n175 & n2565 ;
  assign n2600 = n2598 | n2599 ;
  assign n2601 = n2600 ^ x35 ^ 1'b0 ;
  assign n2602 = n2601 ^ n2593 ^ n2184 ;
  assign n2603 = ( n2184 & n2593 ) | ( n2184 & n2601 ) | ( n2593 & n2601 ) ;
  assign n2604 = x67 & n2560 ;
  assign n2605 = ( x69 & n2567 ) | ( x69 & n2604 ) | ( n2567 & n2604 ) ;
  assign n2606 = n2604 | n2605 ;
  assign n2607 = x68 & ~n2562 ;
  assign n2608 = ( x68 & n2606 ) | ( x68 & ~n2607 ) | ( n2606 & ~n2607 ) ;
  assign n2609 = n172 & n2565 ;
  assign n2610 = n2608 | n2609 ;
  assign n2611 = n2610 ^ x35 ^ 1'b0 ;
  assign n2612 = ( n2186 & n2603 ) | ( n2186 & n2611 ) | ( n2603 & n2611 ) ;
  assign n2613 = n2611 ^ n2603 ^ n2186 ;
  assign n2614 = x68 & n2560 ;
  assign n2615 = ( x70 & n2567 ) | ( x70 & n2614 ) | ( n2567 & n2614 ) ;
  assign n2616 = n2614 | n2615 ;
  assign n2617 = x69 & ~n2562 ;
  assign n2618 = ( x69 & n2616 ) | ( x69 & ~n2617 ) | ( n2616 & ~n2617 ) ;
  assign n2619 = n168 & n2565 ;
  assign n2620 = n2618 | n2619 ;
  assign n2621 = n2620 ^ x35 ^ 1'b0 ;
  assign n2622 = ( n2188 & n2612 ) | ( n2188 & n2621 ) | ( n2612 & n2621 ) ;
  assign n2623 = n2621 ^ n2612 ^ n2188 ;
  assign n2624 = x69 & n2560 ;
  assign n2625 = ( x71 & n2567 ) | ( x71 & n2624 ) | ( n2567 & n2624 ) ;
  assign n2626 = n2624 | n2625 ;
  assign n2627 = x70 & ~n2562 ;
  assign n2628 = ( x70 & n2626 ) | ( x70 & ~n2627 ) | ( n2626 & ~n2627 ) ;
  assign n2629 = n328 & n2565 ;
  assign n2630 = n2628 | n2629 ;
  assign n2631 = n2630 ^ x35 ^ 1'b0 ;
  assign n2632 = ( n2198 & n2622 ) | ( n2198 & n2631 ) | ( n2622 & n2631 ) ;
  assign n2633 = n2631 ^ n2622 ^ n2198 ;
  assign n2634 = x70 & n2560 ;
  assign n2635 = ( x72 & n2567 ) | ( x72 & n2634 ) | ( n2567 & n2634 ) ;
  assign n2636 = n2634 | n2635 ;
  assign n2637 = x71 & ~n2562 ;
  assign n2638 = ( x71 & n2636 ) | ( x71 & ~n2637 ) | ( n2636 & ~n2637 ) ;
  assign n2639 = n349 & n2565 ;
  assign n2640 = n2638 | n2639 ;
  assign n2641 = n2640 ^ x35 ^ 1'b0 ;
  assign n2642 = n2641 ^ n2632 ^ n2209 ;
  assign n2643 = ( n2209 & n2632 ) | ( n2209 & n2641 ) | ( n2632 & n2641 ) ;
  assign n2644 = x71 & n2560 ;
  assign n2645 = ( x73 & n2567 ) | ( x73 & n2644 ) | ( n2567 & n2644 ) ;
  assign n2646 = n2644 | n2645 ;
  assign n2647 = x72 & ~n2562 ;
  assign n2648 = ( x72 & n2646 ) | ( x72 & ~n2647 ) | ( n2646 & ~n2647 ) ;
  assign n2649 = n370 & n2565 ;
  assign n2650 = n2648 | n2649 ;
  assign n2651 = n2650 ^ x35 ^ 1'b0 ;
  assign n2652 = ( n2219 & n2643 ) | ( n2219 & n2651 ) | ( n2643 & n2651 ) ;
  assign n2653 = n2651 ^ n2643 ^ n2219 ;
  assign n2654 = x72 & n2560 ;
  assign n2655 = ( x74 & n2567 ) | ( x74 & n2654 ) | ( n2567 & n2654 ) ;
  assign n2656 = n2654 | n2655 ;
  assign n2657 = x73 & ~n2562 ;
  assign n2658 = ( x73 & n2656 ) | ( x73 & ~n2657 ) | ( n2656 & ~n2657 ) ;
  assign n2659 = n504 & n2565 ;
  assign n2660 = n2658 | n2659 ;
  assign n2661 = n2660 ^ x35 ^ 1'b0 ;
  assign n2662 = n2661 ^ n2652 ^ n2228 ;
  assign n2663 = ( n2228 & n2652 ) | ( n2228 & n2661 ) | ( n2652 & n2661 ) ;
  assign n2664 = x73 & n2560 ;
  assign n2665 = ( x75 & n2567 ) | ( x75 & n2664 ) | ( n2567 & n2664 ) ;
  assign n2666 = n2664 | n2665 ;
  assign n2667 = x74 & ~n2562 ;
  assign n2668 = ( x74 & n2666 ) | ( x74 & ~n2667 ) | ( n2666 & ~n2667 ) ;
  assign n2669 = n525 & n2565 ;
  assign n2670 = n2668 | n2669 ;
  assign n2671 = n2670 ^ x35 ^ 1'b0 ;
  assign n2672 = n2671 ^ n2663 ^ n2239 ;
  assign n2673 = ( n2239 & n2663 ) | ( n2239 & n2671 ) | ( n2663 & n2671 ) ;
  assign n2674 = x74 & n2560 ;
  assign n2675 = ( x76 & n2567 ) | ( x76 & n2674 ) | ( n2567 & n2674 ) ;
  assign n2676 = n2674 | n2675 ;
  assign n2677 = x75 & ~n2562 ;
  assign n2678 = ( x75 & n2676 ) | ( x75 & ~n2677 ) | ( n2676 & ~n2677 ) ;
  assign n2679 = n664 & n2565 ;
  assign n2680 = n2678 | n2679 ;
  assign n2681 = n2680 ^ x35 ^ 1'b0 ;
  assign n2682 = n2681 ^ n2673 ^ n2249 ;
  assign n2683 = ( n2249 & n2673 ) | ( n2249 & n2681 ) | ( n2673 & n2681 ) ;
  assign n2684 = x75 & n2560 ;
  assign n2685 = ( x77 & n2567 ) | ( x77 & n2684 ) | ( n2567 & n2684 ) ;
  assign n2686 = n2684 | n2685 ;
  assign n2687 = x76 & ~n2562 ;
  assign n2688 = ( x76 & n2686 ) | ( x76 & ~n2687 ) | ( n2686 & ~n2687 ) ;
  assign n2689 = n690 & n2565 ;
  assign n2690 = n2688 | n2689 ;
  assign n2691 = n2690 ^ x35 ^ 1'b0 ;
  assign n2692 = ( n2258 & n2683 ) | ( n2258 & n2691 ) | ( n2683 & n2691 ) ;
  assign n2693 = n2691 ^ n2683 ^ n2258 ;
  assign n2694 = x76 & n2560 ;
  assign n2695 = ( x78 & n2567 ) | ( x78 & n2694 ) | ( n2567 & n2694 ) ;
  assign n2696 = n2694 | n2695 ;
  assign n2697 = x77 & ~n2562 ;
  assign n2698 = ( x77 & n2696 ) | ( x77 & ~n2697 ) | ( n2696 & ~n2697 ) ;
  assign n2699 = n709 & n2565 ;
  assign n2700 = n2698 | n2699 ;
  assign n2701 = n2700 ^ x35 ^ 1'b0 ;
  assign n2702 = n2701 ^ n2692 ^ n2269 ;
  assign n2703 = ( n2269 & n2692 ) | ( n2269 & n2701 ) | ( n2692 & n2701 ) ;
  assign n2704 = x77 & n2560 ;
  assign n2705 = ( x79 & n2567 ) | ( x79 & n2704 ) | ( n2567 & n2704 ) ;
  assign n2706 = n2704 | n2705 ;
  assign n2707 = x78 & ~n2562 ;
  assign n2708 = ( x78 & n2706 ) | ( x78 & ~n2707 ) | ( n2706 & ~n2707 ) ;
  assign n2709 = n1015 & n2565 ;
  assign n2710 = n2708 | n2709 ;
  assign n2711 = n2710 ^ x35 ^ 1'b0 ;
  assign n2712 = n2711 ^ n2703 ^ n2279 ;
  assign n2713 = ( n2279 & n2703 ) | ( n2279 & n2711 ) | ( n2703 & n2711 ) ;
  assign n2714 = x78 & n2560 ;
  assign n2715 = ( x80 & n2567 ) | ( x80 & n2714 ) | ( n2567 & n2714 ) ;
  assign n2716 = n2714 | n2715 ;
  assign n2717 = x79 & ~n2562 ;
  assign n2718 = ( x79 & n2716 ) | ( x79 & ~n2717 ) | ( n2716 & ~n2717 ) ;
  assign n2719 = n1216 & n2565 ;
  assign n2720 = n2718 | n2719 ;
  assign n2721 = n2720 ^ x35 ^ 1'b0 ;
  assign n2722 = ( n2288 & n2713 ) | ( n2288 & n2721 ) | ( n2713 & n2721 ) ;
  assign n2723 = n2721 ^ n2713 ^ n2288 ;
  assign n2724 = x79 & n2560 ;
  assign n2725 = ( x81 & n2567 ) | ( x81 & n2724 ) | ( n2567 & n2724 ) ;
  assign n2726 = n2724 | n2725 ;
  assign n2727 = x80 & ~n2562 ;
  assign n2728 = ( x80 & n2726 ) | ( x80 & ~n2727 ) | ( n2726 & ~n2727 ) ;
  assign n2729 = n1258 & n2565 ;
  assign n2730 = n2728 | n2729 ;
  assign n2731 = n2730 ^ x35 ^ 1'b0 ;
  assign n2732 = ( n2298 & n2722 ) | ( n2298 & n2731 ) | ( n2722 & n2731 ) ;
  assign n2733 = n2731 ^ n2722 ^ n2298 ;
  assign n2734 = x80 & n2560 ;
  assign n2735 = ( x82 & n2567 ) | ( x82 & n2734 ) | ( n2567 & n2734 ) ;
  assign n2736 = n2734 | n2735 ;
  assign n2737 = x81 & ~n2562 ;
  assign n2738 = ( x81 & n2736 ) | ( x81 & ~n2737 ) | ( n2736 & ~n2737 ) ;
  assign n2739 = n1301 & n2565 ;
  assign n2740 = n2738 | n2739 ;
  assign n2741 = n2740 ^ x35 ^ 1'b0 ;
  assign n2742 = n2741 ^ n2732 ^ n2309 ;
  assign n2743 = ( n2309 & n2732 ) | ( n2309 & n2741 ) | ( n2732 & n2741 ) ;
  assign n2744 = x81 & n2560 ;
  assign n2745 = ( x83 & n2567 ) | ( x83 & n2744 ) | ( n2567 & n2744 ) ;
  assign n2746 = n2744 | n2745 ;
  assign n2747 = x82 & ~n2562 ;
  assign n2748 = ( x82 & n2746 ) | ( x82 & ~n2747 ) | ( n2746 & ~n2747 ) ;
  assign n2749 = n1329 & n2565 ;
  assign n2750 = n2748 | n2749 ;
  assign n2751 = n2750 ^ x35 ^ 1'b0 ;
  assign n2752 = n2751 ^ n2743 ^ n2319 ;
  assign n2753 = ( n2319 & n2743 ) | ( n2319 & n2751 ) | ( n2743 & n2751 ) ;
  assign n2754 = x82 & n2560 ;
  assign n2755 = ( x84 & n2567 ) | ( x84 & n2754 ) | ( n2567 & n2754 ) ;
  assign n2756 = n2754 | n2755 ;
  assign n2757 = x83 & ~n2562 ;
  assign n2758 = ( x83 & n2756 ) | ( x83 & ~n2757 ) | ( n2756 & ~n2757 ) ;
  assign n2759 = n1355 & n2565 ;
  assign n2760 = n2758 | n2759 ;
  assign n2761 = n2760 ^ x35 ^ 1'b0 ;
  assign n2762 = n2761 ^ n2753 ^ n2328 ;
  assign n2763 = ( n2328 & n2753 ) | ( n2328 & n2761 ) | ( n2753 & n2761 ) ;
  assign n2764 = x83 & n2560 ;
  assign n2765 = ( x85 & n2567 ) | ( x85 & n2764 ) | ( n2567 & n2764 ) ;
  assign n2766 = n2764 | n2765 ;
  assign n2767 = x84 & ~n2562 ;
  assign n2768 = ( x84 & n2766 ) | ( x84 & ~n2767 ) | ( n2766 & ~n2767 ) ;
  assign n2769 = n1392 & n2565 ;
  assign n2770 = n2768 | n2769 ;
  assign n2771 = n2770 ^ x35 ^ 1'b0 ;
  assign n2772 = n2771 ^ n2763 ^ n2339 ;
  assign n2773 = ( n2339 & n2763 ) | ( n2339 & n2771 ) | ( n2763 & n2771 ) ;
  assign n2774 = x84 & n2560 ;
  assign n2775 = ( x86 & n2567 ) | ( x86 & n2774 ) | ( n2567 & n2774 ) ;
  assign n2776 = n2774 | n2775 ;
  assign n2777 = x85 & ~n2562 ;
  assign n2778 = ( x85 & n2776 ) | ( x85 & ~n2777 ) | ( n2776 & ~n2777 ) ;
  assign n2779 = n1419 & n2565 ;
  assign n2780 = n2778 | n2779 ;
  assign n2781 = n2780 ^ x35 ^ 1'b0 ;
  assign n2782 = ( n2348 & n2773 ) | ( n2348 & n2781 ) | ( n2773 & n2781 ) ;
  assign n2783 = n2781 ^ n2773 ^ n2348 ;
  assign n2784 = x85 & n2560 ;
  assign n2785 = ( x87 & n2567 ) | ( x87 & n2784 ) | ( n2567 & n2784 ) ;
  assign n2786 = n2784 | n2785 ;
  assign n2787 = x86 & ~n2562 ;
  assign n2788 = ( x86 & n2786 ) | ( x86 & ~n2787 ) | ( n2786 & ~n2787 ) ;
  assign n2789 = n1484 & n2565 ;
  assign n2790 = n2788 | n2789 ;
  assign n2791 = n2790 ^ x35 ^ 1'b0 ;
  assign n2792 = ( n2359 & n2782 ) | ( n2359 & n2791 ) | ( n2782 & n2791 ) ;
  assign n2793 = n2791 ^ n2782 ^ n2359 ;
  assign n2794 = x86 & n2560 ;
  assign n2795 = ( x88 & n2567 ) | ( x88 & n2794 ) | ( n2567 & n2794 ) ;
  assign n2796 = n2794 | n2795 ;
  assign n2797 = x87 & ~n2562 ;
  assign n2798 = ( x87 & n2796 ) | ( x87 & ~n2797 ) | ( n2796 & ~n2797 ) ;
  assign n2799 = n1569 & n2565 ;
  assign n2800 = n2798 | n2799 ;
  assign n2801 = n2800 ^ x35 ^ 1'b0 ;
  assign n2802 = n2801 ^ n2792 ^ n2369 ;
  assign n2803 = ( n2369 & n2792 ) | ( n2369 & n2801 ) | ( n2792 & n2801 ) ;
  assign n2804 = x87 & n2560 ;
  assign n2805 = ( x89 & n2567 ) | ( x89 & n2804 ) | ( n2567 & n2804 ) ;
  assign n2806 = n2804 | n2805 ;
  assign n2807 = x88 & ~n2562 ;
  assign n2808 = ( x88 & n2806 ) | ( x88 & ~n2807 ) | ( n2806 & ~n2807 ) ;
  assign n2809 = n1654 & n2565 ;
  assign n2810 = n2808 | n2809 ;
  assign n2811 = n2810 ^ x35 ^ 1'b0 ;
  assign n2812 = ( n2379 & n2803 ) | ( n2379 & n2811 ) | ( n2803 & n2811 ) ;
  assign n2813 = n2811 ^ n2803 ^ n2379 ;
  assign n2814 = x88 & n2560 ;
  assign n2815 = ( x90 & n2567 ) | ( x90 & n2814 ) | ( n2567 & n2814 ) ;
  assign n2816 = n2814 | n2815 ;
  assign n2817 = x89 & ~n2562 ;
  assign n2818 = ( x89 & n2816 ) | ( x89 & ~n2817 ) | ( n2816 & ~n2817 ) ;
  assign n2819 = n1741 & n2565 ;
  assign n2820 = n2818 | n2819 ;
  assign n2821 = n2820 ^ x35 ^ 1'b0 ;
  assign n2822 = ( n2388 & n2812 ) | ( n2388 & n2821 ) | ( n2812 & n2821 ) ;
  assign n2823 = n2821 ^ n2812 ^ n2388 ;
  assign n2824 = x89 & n2560 ;
  assign n2825 = ( x91 & n2567 ) | ( x91 & n2824 ) | ( n2567 & n2824 ) ;
  assign n2826 = n2824 | n2825 ;
  assign n2827 = x90 & ~n2562 ;
  assign n2828 = ( x90 & n2826 ) | ( x90 & ~n2827 ) | ( n2826 & ~n2827 ) ;
  assign n2829 = n2114 & n2565 ;
  assign n2830 = n2828 | n2829 ;
  assign n2831 = n2830 ^ x35 ^ 1'b0 ;
  assign n2832 = n2831 ^ n2822 ^ n2399 ;
  assign n2833 = ( n2399 & n2822 ) | ( n2399 & n2831 ) | ( n2822 & n2831 ) ;
  assign n2834 = x90 & n2560 ;
  assign n2835 = ( x92 & n2567 ) | ( x92 & n2834 ) | ( n2567 & n2834 ) ;
  assign n2836 = n2834 | n2835 ;
  assign n2837 = x91 & ~n2562 ;
  assign n2838 = ( x91 & n2836 ) | ( x91 & ~n2837 ) | ( n2836 & ~n2837 ) ;
  assign n2839 = n2420 & n2565 ;
  assign n2840 = n2838 | n2839 ;
  assign n2841 = n2840 ^ x35 ^ 1'b0 ;
  assign n2842 = n2841 ^ n2833 ^ n2409 ;
  assign n2843 = ( n2409 & n2833 ) | ( n2409 & n2841 ) | ( n2833 & n2841 ) ;
  assign n2844 = x91 & n2560 ;
  assign n2845 = ( x93 & n2567 ) | ( x93 & n2844 ) | ( n2567 & n2844 ) ;
  assign n2846 = n2844 | n2845 ;
  assign n2847 = x92 & ~n2562 ;
  assign n2848 = ( x92 & n2846 ) | ( x92 & ~n2847 ) | ( n2846 & ~n2847 ) ;
  assign n2849 = n2476 & n2565 ;
  assign n2850 = n2848 | n2849 ;
  assign n2851 = n2850 ^ x35 ^ 1'b0 ;
  assign n2852 = n2851 ^ n2843 ^ n2419 ;
  assign n2853 = ( n2419 & n2843 ) | ( n2419 & n2851 ) | ( n2843 & n2851 ) ;
  assign n2854 = n2527 ^ x95 ^ x94 ;
  assign n2855 = x93 & n1058 ;
  assign n2856 = ( x95 & n1065 ) | ( x95 & n2855 ) | ( n1065 & n2855 ) ;
  assign n2857 = n2855 | n2856 ;
  assign n2858 = x94 & ~n1060 ;
  assign n2859 = ( x94 & n2857 ) | ( x94 & ~n2858 ) | ( n2857 & ~n2858 ) ;
  assign n2860 = n1063 & n2854 ;
  assign n2861 = n2859 | n2860 ;
  assign n2862 = n2861 ^ x41 ^ 1'b0 ;
  assign n2863 = n2862 ^ n2429 ^ n2151 ;
  assign n2864 = ( n2151 & n2429 ) | ( n2151 & n2862 ) | ( n2429 & n2862 ) ;
  assign n2865 = ( x94 & x95 ) | ( x94 & n2527 ) | ( x95 & n2527 ) ;
  assign n2866 = x93 & n2156 ;
  assign n2867 = ( x95 & n2163 ) | ( x95 & n2866 ) | ( n2163 & n2866 ) ;
  assign n2868 = n2866 | n2867 ;
  assign n2869 = x94 & ~n2158 ;
  assign n2870 = ( x94 & n2868 ) | ( x94 & ~n2869 ) | ( n2868 & ~n2869 ) ;
  assign n2871 = n2161 & n2854 ;
  assign n2872 = n2870 | n2871 ;
  assign n2873 = n2872 ^ x38 ^ 1'b0 ;
  assign n2874 = ( n2140 & n2441 ) | ( n2140 & n2873 ) | ( n2441 & n2873 ) ;
  assign n2875 = n2873 ^ n2441 ^ n2140 ;
  assign n2876 = x92 & n2560 ;
  assign n2877 = ( x94 & n2567 ) | ( x94 & n2876 ) | ( n2567 & n2876 ) ;
  assign n2878 = n2876 | n2877 ;
  assign n2879 = x93 & ~n2562 ;
  assign n2880 = ( x93 & n2878 ) | ( x93 & ~n2879 ) | ( n2878 & ~n2879 ) ;
  assign n2881 = n2518 & n2565 ;
  assign n2882 = n2880 | n2881 ;
  assign n2883 = n2882 ^ x35 ^ 1'b0 ;
  assign n2884 = ( n2451 & n2853 ) | ( n2451 & n2883 ) | ( n2853 & n2883 ) ;
  assign n2885 = n2883 ^ n2853 ^ n2451 ;
  assign n2886 = x93 & n888 ;
  assign n2887 = ( x95 & n878 ) | ( x95 & n2886 ) | ( n878 & n2886 ) ;
  assign n2888 = n2886 | n2887 ;
  assign n2889 = x94 & ~n877 ;
  assign n2890 = ( x94 & n2888 ) | ( x94 & ~n2889 ) | ( n2888 & ~n2889 ) ;
  assign n2891 = n880 & n2854 ;
  assign n2892 = n2890 | n2891 ;
  assign n2893 = n2892 ^ x44 ^ 1'b0 ;
  assign n2894 = n2893 ^ n2460 ^ n2119 ;
  assign n2895 = ( n2119 & n2460 ) | ( n2119 & n2893 ) | ( n2460 & n2893 ) ;
  assign n2896 = x93 & n2560 ;
  assign n2897 = ( x95 & n2567 ) | ( x95 & n2896 ) | ( n2567 & n2896 ) ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = x94 & ~n2562 ;
  assign n2900 = ( x94 & n2898 ) | ( x94 & ~n2899 ) | ( n2898 & ~n2899 ) ;
  assign n2901 = n2565 & n2854 ;
  assign n2902 = n2900 | n2901 ;
  assign n2903 = n2902 ^ x35 ^ 1'b0 ;
  assign n2904 = ( n2471 & n2884 ) | ( n2471 & n2903 ) | ( n2884 & n2903 ) ;
  assign n2905 = n2903 ^ n2884 ^ n2471 ;
  assign n2906 = x94 & n1058 ;
  assign n2907 = n2865 ^ x96 ^ x95 ;
  assign n2908 = ( x95 & x96 ) | ( x95 & n2865 ) | ( x96 & n2865 ) ;
  assign n2909 = ( x96 & n1065 ) | ( x96 & n2906 ) | ( n1065 & n2906 ) ;
  assign n2910 = n2906 | n2909 ;
  assign n2911 = x95 & ~n1060 ;
  assign n2912 = ( x95 & n2910 ) | ( x95 & ~n2911 ) | ( n2910 & ~n2911 ) ;
  assign n2913 = n1063 & n2907 ;
  assign n2914 = n2912 | n2913 ;
  assign n2915 = n2914 ^ x41 ^ 1'b0 ;
  assign n2916 = ( n2430 & n2482 ) | ( n2430 & n2915 ) | ( n2482 & n2915 ) ;
  assign n2917 = n2915 ^ n2482 ^ n2430 ;
  assign n2918 = x94 & n2560 ;
  assign n2919 = ( x96 & n2567 ) | ( x96 & n2918 ) | ( n2567 & n2918 ) ;
  assign n2920 = n2918 | n2919 ;
  assign n2921 = x95 & ~n2562 ;
  assign n2922 = ( x95 & n2920 ) | ( x95 & ~n2921 ) | ( n2920 & ~n2921 ) ;
  assign n2923 = n2565 & n2907 ;
  assign n2924 = n2922 | n2923 ;
  assign n2925 = n2924 ^ x35 ^ 1'b0 ;
  assign n2926 = ( n2503 & n2904 ) | ( n2503 & n2925 ) | ( n2904 & n2925 ) ;
  assign n2927 = n2925 ^ n2904 ^ n2503 ;
  assign n2928 = x94 & n2156 ;
  assign n2929 = ( x96 & n2163 ) | ( x96 & n2928 ) | ( n2163 & n2928 ) ;
  assign n2930 = n2928 | n2929 ;
  assign n2931 = x95 & ~n2158 ;
  assign n2932 = ( x95 & n2930 ) | ( x95 & ~n2931 ) | ( n2930 & ~n2931 ) ;
  assign n2933 = n2161 & n2907 ;
  assign n2934 = n2932 | n2933 ;
  assign n2935 = n2934 ^ x38 ^ 1'b0 ;
  assign n2936 = ( n2440 & n2512 ) | ( n2440 & n2935 ) | ( n2512 & n2935 ) ;
  assign n2937 = n2935 ^ n2512 ^ n2440 ;
  assign n2938 = x94 & n888 ;
  assign n2939 = ( x96 & n878 ) | ( x96 & n2938 ) | ( n878 & n2938 ) ;
  assign n2940 = n2938 | n2939 ;
  assign n2941 = x95 & ~n877 ;
  assign n2942 = ( x95 & n2940 ) | ( x95 & ~n2941 ) | ( n2940 & ~n2941 ) ;
  assign n2943 = n880 & n2907 ;
  assign n2944 = n2942 | n2943 ;
  assign n2945 = n2944 ^ x44 ^ 1'b0 ;
  assign n2946 = ( n2461 & n2493 ) | ( n2461 & n2945 ) | ( n2493 & n2945 ) ;
  assign n2947 = n2945 ^ n2493 ^ n2461 ;
  assign n2948 = x93 & n744 ;
  assign n2949 = ( x95 & n730 ) | ( x95 & n2948 ) | ( n730 & n2948 ) ;
  assign n2950 = n2948 | n2949 ;
  assign n2951 = x94 & ~n732 ;
  assign n2952 = ( x94 & n2950 ) | ( x94 & ~n2951 ) | ( n2950 & ~n2951 ) ;
  assign n2953 = n731 & n2854 ;
  assign n2954 = n2952 | n2953 ;
  assign n2955 = n140 & n1329 ;
  assign n2956 = x81 & n133 ;
  assign n2957 = ( x83 & n142 ) | ( x83 & n2956 ) | ( n142 & n2956 ) ;
  assign n2958 = x76 & n325 ;
  assign n2959 = n2956 | n2957 ;
  assign n2960 = x82 & ~n134 ;
  assign n2961 = ( x82 & n2959 ) | ( x82 & ~n2960 ) | ( n2959 & ~n2960 ) ;
  assign n2962 = x78 & n208 ;
  assign n2963 = n2955 | n2961 ;
  assign n2964 = ( x80 & n194 ) | ( x80 & n2962 ) | ( n194 & n2962 ) ;
  assign n2965 = n2962 | n2964 ;
  assign n2966 = x77 & ~n242 ;
  assign n2967 = ( x77 & n2958 ) | ( x77 & ~n2966 ) | ( n2958 & ~n2966 ) ;
  assign n2968 = x79 & ~n192 ;
  assign n2969 = ( x79 & n2965 ) | ( x79 & ~n2968 ) | ( n2965 & ~n2968 ) ;
  assign n2970 = n197 & n1216 ;
  assign n2971 = n2969 | n2970 ;
  assign n2972 = n2971 ^ x62 ^ 1'b0 ;
  assign n2973 = n2954 ^ x47 ^ 1'b0 ;
  assign n2974 = ( n2074 & ~n2967 ) | ( n2074 & n2972 ) | ( ~n2967 & n2972 ) ;
  assign n2975 = n2972 ^ n2967 ^ n2074 ;
  assign n2976 = n2963 ^ x59 ^ 1'b0 ;
  assign n2977 = n2976 ^ n2975 ^ n2078 ;
  assign n2978 = ( n2078 & ~n2975 ) | ( n2078 & n2976 ) | ( ~n2975 & n2976 ) ;
  assign n2979 = x84 & n263 ;
  assign n2980 = ( x86 & n264 ) | ( x86 & n2979 ) | ( n264 & n2979 ) ;
  assign n2981 = n2979 | n2980 ;
  assign n2982 = x85 & ~n260 ;
  assign n2983 = ( x85 & n2981 ) | ( x85 & ~n2982 ) | ( n2981 & ~n2982 ) ;
  assign n2984 = n272 & n1419 ;
  assign n2985 = n2983 | n2984 ;
  assign n2986 = n2985 ^ x56 ^ 1'b0 ;
  assign n2987 = n2986 ^ n2977 ^ n2088 ;
  assign n2988 = ( n2088 & ~n2977 ) | ( n2088 & n2986 ) | ( ~n2977 & n2986 ) ;
  assign n2989 = x87 & n408 ;
  assign n2990 = ( x89 & n403 ) | ( x89 & n2989 ) | ( n403 & n2989 ) ;
  assign n2991 = n2989 | n2990 ;
  assign n2992 = x88 & ~n410 ;
  assign n2993 = ( x88 & n2991 ) | ( x88 & ~n2992 ) | ( n2991 & ~n2992 ) ;
  assign n2994 = n402 & n1654 ;
  assign n2995 = n2993 | n2994 ;
  assign n2996 = n2995 ^ x53 ^ 1'b0 ;
  assign n2997 = n2996 ^ n2987 ^ n2098 ;
  assign n2998 = ( n2098 & n2987 ) | ( n2098 & ~n2996 ) | ( n2987 & ~n2996 ) ;
  assign n2999 = x90 & n561 ;
  assign n3000 = ( x92 & n551 ) | ( x92 & n2999 ) | ( n551 & n2999 ) ;
  assign n3001 = n2999 | n3000 ;
  assign n3002 = x91 & ~n550 ;
  assign n3003 = ( x91 & n3001 ) | ( x91 & ~n3002 ) | ( n3001 & ~n3002 ) ;
  assign n3004 = n553 & n2420 ;
  assign n3005 = n3003 | n3004 ;
  assign n3006 = n3005 ^ x50 ^ 1'b0 ;
  assign n3007 = ( n2109 & n2997 ) | ( n2109 & n3006 ) | ( n2997 & n3006 ) ;
  assign n3008 = n3006 ^ n2997 ^ n2109 ;
  assign n3009 = ( n2130 & n2973 ) | ( n2130 & n3008 ) | ( n2973 & n3008 ) ;
  assign n3010 = n3008 ^ n2973 ^ n2130 ;
  assign n3011 = x31 ^ x30 ^ 1'b0 ;
  assign n3012 = x30 ^ x29 ^ 1'b0 ;
  assign n3013 = x32 ^ x31 ^ 1'b0 ;
  assign n3014 = n3011 & ~n3012 ;
  assign n3015 = n3012 & ~n3013 ;
  assign n3016 = ~x65 & n3015 ;
  assign n3017 = n3012 & n3013 ;
  assign n3018 = x64 & n3014 ;
  assign n3019 = ( n3015 & ~n3016 ) | ( n3015 & n3018 ) | ( ~n3016 & n3018 ) ;
  assign n3020 = ( n190 & n3017 ) | ( n190 & n3018 ) | ( n3017 & n3018 ) ;
  assign n3021 = n139 & n3017 ;
  assign n3022 = n3019 | n3020 ;
  assign n3023 = x65 & ~n3014 ;
  assign n3024 = ( n3011 & ~n3012 ) | ( n3011 & n3013 ) | ( ~n3012 & n3013 ) ;
  assign n3025 = ~n3011 & n3024 ;
  assign n3026 = x64 & n3025 ;
  assign n3027 = ( x66 & n3015 ) | ( x66 & n3026 ) | ( n3015 & n3026 ) ;
  assign n3028 = n3026 | n3027 ;
  assign n3029 = x64 & n3012 ;
  assign n3030 = ( x65 & ~n3023 ) | ( x65 & n3028 ) | ( ~n3023 & n3028 ) ;
  assign n3031 = x32 & ~n3029 ;
  assign n3032 = n3021 | n3030 ;
  assign n3033 = n3032 ^ x32 ^ 1'b0 ;
  assign n3034 = n3022 ^ x32 ^ 1'b0 ;
  assign n3035 = n3031 & n3034 ;
  assign n3036 = n3035 ^ n3033 ^ 1'b0 ;
  assign n3037 = n3033 & n3035 ;
  assign n3038 = n3034 ^ n3031 ^ 1'b0 ;
  assign n3039 = x65 & n3025 ;
  assign n3040 = ( x67 & n3015 ) | ( x67 & n3039 ) | ( n3015 & n3039 ) ;
  assign n3041 = n3039 | n3040 ;
  assign n3042 = x66 & ~n3014 ;
  assign n3043 = ( x66 & n3041 ) | ( x66 & ~n3042 ) | ( n3041 & ~n3042 ) ;
  assign n3044 = n161 & n3017 ;
  assign n3045 = n3043 | n3044 ;
  assign n3046 = n3045 ^ x32 ^ 1'b0 ;
  assign n3047 = ( n2585 & n3037 ) | ( n2585 & n3046 ) | ( n3037 & n3046 ) ;
  assign n3048 = n3046 ^ n3037 ^ n2585 ;
  assign n3049 = x66 & n3025 ;
  assign n3050 = ( x68 & n3015 ) | ( x68 & n3049 ) | ( n3015 & n3049 ) ;
  assign n3051 = n3049 | n3050 ;
  assign n3052 = x67 & ~n3014 ;
  assign n3053 = ( x67 & n3051 ) | ( x67 & ~n3052 ) | ( n3051 & ~n3052 ) ;
  assign n3054 = n175 & n3017 ;
  assign n3055 = n3053 | n3054 ;
  assign n3056 = n3055 ^ x32 ^ 1'b0 ;
  assign n3057 = n3056 ^ n3047 ^ n2588 ;
  assign n3058 = ( n2588 & n3047 ) | ( n2588 & n3056 ) | ( n3047 & n3056 ) ;
  assign n3059 = x67 & n3025 ;
  assign n3060 = ( x69 & n3015 ) | ( x69 & n3059 ) | ( n3015 & n3059 ) ;
  assign n3061 = n3059 | n3060 ;
  assign n3062 = x68 & ~n3014 ;
  assign n3063 = ( x68 & n3061 ) | ( x68 & ~n3062 ) | ( n3061 & ~n3062 ) ;
  assign n3064 = n172 & n3017 ;
  assign n3065 = n3063 | n3064 ;
  assign n3066 = n3065 ^ x32 ^ 1'b0 ;
  assign n3067 = n3066 ^ n3058 ^ n2590 ;
  assign n3068 = ( n2590 & n3058 ) | ( n2590 & n3066 ) | ( n3058 & n3066 ) ;
  assign n3069 = x68 & n3025 ;
  assign n3070 = ( x70 & n3015 ) | ( x70 & n3069 ) | ( n3015 & n3069 ) ;
  assign n3071 = n3069 | n3070 ;
  assign n3072 = x69 & ~n3014 ;
  assign n3073 = ( x69 & n3071 ) | ( x69 & ~n3072 ) | ( n3071 & ~n3072 ) ;
  assign n3074 = n168 & n3017 ;
  assign n3075 = n3073 | n3074 ;
  assign n3076 = n3075 ^ x32 ^ 1'b0 ;
  assign n3077 = ( n2592 & n3068 ) | ( n2592 & n3076 ) | ( n3068 & n3076 ) ;
  assign n3078 = n3076 ^ n3068 ^ n2592 ;
  assign n3079 = x69 & n3025 ;
  assign n3080 = ( x71 & n3015 ) | ( x71 & n3079 ) | ( n3015 & n3079 ) ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = x70 & ~n3014 ;
  assign n3083 = ( x70 & n3081 ) | ( x70 & ~n3082 ) | ( n3081 & ~n3082 ) ;
  assign n3084 = n328 & n3017 ;
  assign n3085 = n3083 | n3084 ;
  assign n3086 = n3085 ^ x32 ^ 1'b0 ;
  assign n3087 = n3086 ^ n3077 ^ n2602 ;
  assign n3088 = ( n2602 & n3077 ) | ( n2602 & n3086 ) | ( n3077 & n3086 ) ;
  assign n3089 = x70 & n3025 ;
  assign n3090 = ( x72 & n3015 ) | ( x72 & n3089 ) | ( n3015 & n3089 ) ;
  assign n3091 = n3089 | n3090 ;
  assign n3092 = x71 & ~n3014 ;
  assign n3093 = ( x71 & n3091 ) | ( x71 & ~n3092 ) | ( n3091 & ~n3092 ) ;
  assign n3094 = n349 & n3017 ;
  assign n3095 = n3093 | n3094 ;
  assign n3096 = n3095 ^ x32 ^ 1'b0 ;
  assign n3097 = ( n2613 & n3088 ) | ( n2613 & n3096 ) | ( n3088 & n3096 ) ;
  assign n3098 = n3096 ^ n3088 ^ n2613 ;
  assign n3099 = x71 & n3025 ;
  assign n3100 = ( x73 & n3015 ) | ( x73 & n3099 ) | ( n3015 & n3099 ) ;
  assign n3101 = n3099 | n3100 ;
  assign n3102 = x72 & ~n3014 ;
  assign n3103 = ( x72 & n3101 ) | ( x72 & ~n3102 ) | ( n3101 & ~n3102 ) ;
  assign n3104 = n370 & n3017 ;
  assign n3105 = n3103 | n3104 ;
  assign n3106 = n3105 ^ x32 ^ 1'b0 ;
  assign n3107 = ( n2623 & n3097 ) | ( n2623 & n3106 ) | ( n3097 & n3106 ) ;
  assign n3108 = n3106 ^ n3097 ^ n2623 ;
  assign n3109 = x72 & n3025 ;
  assign n3110 = ( x74 & n3015 ) | ( x74 & n3109 ) | ( n3015 & n3109 ) ;
  assign n3111 = n3109 | n3110 ;
  assign n3112 = x73 & ~n3014 ;
  assign n3113 = ( x73 & n3111 ) | ( x73 & ~n3112 ) | ( n3111 & ~n3112 ) ;
  assign n3114 = n504 & n3017 ;
  assign n3115 = n3113 | n3114 ;
  assign n3116 = n3115 ^ x32 ^ 1'b0 ;
  assign n3117 = n3116 ^ n3107 ^ n2633 ;
  assign n3118 = ( n2633 & n3107 ) | ( n2633 & n3116 ) | ( n3107 & n3116 ) ;
  assign n3119 = x73 & n3025 ;
  assign n3120 = ( x75 & n3015 ) | ( x75 & n3119 ) | ( n3015 & n3119 ) ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = x74 & ~n3014 ;
  assign n3123 = ( x74 & n3121 ) | ( x74 & ~n3122 ) | ( n3121 & ~n3122 ) ;
  assign n3124 = n525 & n3017 ;
  assign n3125 = n3123 | n3124 ;
  assign n3126 = n3125 ^ x32 ^ 1'b0 ;
  assign n3127 = ( n2642 & n3118 ) | ( n2642 & n3126 ) | ( n3118 & n3126 ) ;
  assign n3128 = n3126 ^ n3118 ^ n2642 ;
  assign n3129 = x74 & n3025 ;
  assign n3130 = ( x76 & n3015 ) | ( x76 & n3129 ) | ( n3015 & n3129 ) ;
  assign n3131 = n3129 | n3130 ;
  assign n3132 = x75 & ~n3014 ;
  assign n3133 = ( x75 & n3131 ) | ( x75 & ~n3132 ) | ( n3131 & ~n3132 ) ;
  assign n3134 = n664 & n3017 ;
  assign n3135 = n3133 | n3134 ;
  assign n3136 = n3135 ^ x32 ^ 1'b0 ;
  assign n3137 = n3136 ^ n3127 ^ n2653 ;
  assign n3138 = ( n2653 & n3127 ) | ( n2653 & n3136 ) | ( n3127 & n3136 ) ;
  assign n3139 = x75 & n3025 ;
  assign n3140 = ( x77 & n3015 ) | ( x77 & n3139 ) | ( n3015 & n3139 ) ;
  assign n3141 = n3139 | n3140 ;
  assign n3142 = x76 & ~n3014 ;
  assign n3143 = ( x76 & n3141 ) | ( x76 & ~n3142 ) | ( n3141 & ~n3142 ) ;
  assign n3144 = n690 & n3017 ;
  assign n3145 = n3143 | n3144 ;
  assign n3146 = n3145 ^ x32 ^ 1'b0 ;
  assign n3147 = ( n2662 & n3138 ) | ( n2662 & n3146 ) | ( n3138 & n3146 ) ;
  assign n3148 = n3146 ^ n3138 ^ n2662 ;
  assign n3149 = x76 & n3025 ;
  assign n3150 = ( x78 & n3015 ) | ( x78 & n3149 ) | ( n3015 & n3149 ) ;
  assign n3151 = n3149 | n3150 ;
  assign n3152 = x77 & ~n3014 ;
  assign n3153 = ( x77 & n3151 ) | ( x77 & ~n3152 ) | ( n3151 & ~n3152 ) ;
  assign n3154 = n709 & n3017 ;
  assign n3155 = n3153 | n3154 ;
  assign n3156 = n3155 ^ x32 ^ 1'b0 ;
  assign n3157 = n3156 ^ n3147 ^ n2672 ;
  assign n3158 = ( n2672 & n3147 ) | ( n2672 & n3156 ) | ( n3147 & n3156 ) ;
  assign n3159 = x77 & n3025 ;
  assign n3160 = ( x79 & n3015 ) | ( x79 & n3159 ) | ( n3015 & n3159 ) ;
  assign n3161 = n3159 | n3160 ;
  assign n3162 = x78 & ~n3014 ;
  assign n3163 = ( x78 & n3161 ) | ( x78 & ~n3162 ) | ( n3161 & ~n3162 ) ;
  assign n3164 = n1015 & n3017 ;
  assign n3165 = n3163 | n3164 ;
  assign n3166 = n3165 ^ x32 ^ 1'b0 ;
  assign n3167 = n3166 ^ n3158 ^ n2682 ;
  assign n3168 = ( n2682 & n3158 ) | ( n2682 & n3166 ) | ( n3158 & n3166 ) ;
  assign n3169 = x78 & n3025 ;
  assign n3170 = ( x80 & n3015 ) | ( x80 & n3169 ) | ( n3015 & n3169 ) ;
  assign n3171 = n3169 | n3170 ;
  assign n3172 = x79 & ~n3014 ;
  assign n3173 = ( x79 & n3171 ) | ( x79 & ~n3172 ) | ( n3171 & ~n3172 ) ;
  assign n3174 = n1216 & n3017 ;
  assign n3175 = n3173 | n3174 ;
  assign n3176 = n3175 ^ x32 ^ 1'b0 ;
  assign n3177 = n3176 ^ n3168 ^ n2693 ;
  assign n3178 = ( n2693 & n3168 ) | ( n2693 & n3176 ) | ( n3168 & n3176 ) ;
  assign n3179 = x79 & n3025 ;
  assign n3180 = ( x81 & n3015 ) | ( x81 & n3179 ) | ( n3015 & n3179 ) ;
  assign n3181 = n3179 | n3180 ;
  assign n3182 = x80 & ~n3014 ;
  assign n3183 = ( x80 & n3181 ) | ( x80 & ~n3182 ) | ( n3181 & ~n3182 ) ;
  assign n3184 = n1258 & n3017 ;
  assign n3185 = n3183 | n3184 ;
  assign n3186 = n3185 ^ x32 ^ 1'b0 ;
  assign n3187 = n3186 ^ n3178 ^ n2702 ;
  assign n3188 = ( n2702 & n3178 ) | ( n2702 & n3186 ) | ( n3178 & n3186 ) ;
  assign n3189 = x80 & n3025 ;
  assign n3190 = ( x82 & n3015 ) | ( x82 & n3189 ) | ( n3015 & n3189 ) ;
  assign n3191 = n3189 | n3190 ;
  assign n3192 = x81 & ~n3014 ;
  assign n3193 = ( x81 & n3191 ) | ( x81 & ~n3192 ) | ( n3191 & ~n3192 ) ;
  assign n3194 = n1301 & n3017 ;
  assign n3195 = n3193 | n3194 ;
  assign n3196 = n3195 ^ x32 ^ 1'b0 ;
  assign n3197 = n3196 ^ n3188 ^ n2712 ;
  assign n3198 = ( n2712 & n3188 ) | ( n2712 & n3196 ) | ( n3188 & n3196 ) ;
  assign n3199 = x81 & n3025 ;
  assign n3200 = ( x83 & n3015 ) | ( x83 & n3199 ) | ( n3015 & n3199 ) ;
  assign n3201 = n3199 | n3200 ;
  assign n3202 = x82 & ~n3014 ;
  assign n3203 = ( x82 & n3201 ) | ( x82 & ~n3202 ) | ( n3201 & ~n3202 ) ;
  assign n3204 = n1329 & n3017 ;
  assign n3205 = n3203 | n3204 ;
  assign n3206 = n3205 ^ x32 ^ 1'b0 ;
  assign n3207 = ( n2723 & n3198 ) | ( n2723 & n3206 ) | ( n3198 & n3206 ) ;
  assign n3208 = n3206 ^ n3198 ^ n2723 ;
  assign n3209 = x82 & n3025 ;
  assign n3210 = ( x84 & n3015 ) | ( x84 & n3209 ) | ( n3015 & n3209 ) ;
  assign n3211 = n3209 | n3210 ;
  assign n3212 = x83 & ~n3014 ;
  assign n3213 = ( x83 & n3211 ) | ( x83 & ~n3212 ) | ( n3211 & ~n3212 ) ;
  assign n3214 = n1355 & n3017 ;
  assign n3215 = n3213 | n3214 ;
  assign n3216 = n3215 ^ x32 ^ 1'b0 ;
  assign n3217 = ( n2733 & n3207 ) | ( n2733 & n3216 ) | ( n3207 & n3216 ) ;
  assign n3218 = n3216 ^ n3207 ^ n2733 ;
  assign n3219 = x83 & n3025 ;
  assign n3220 = ( x85 & n3015 ) | ( x85 & n3219 ) | ( n3015 & n3219 ) ;
  assign n3221 = n3219 | n3220 ;
  assign n3222 = x84 & ~n3014 ;
  assign n3223 = ( x84 & n3221 ) | ( x84 & ~n3222 ) | ( n3221 & ~n3222 ) ;
  assign n3224 = n1392 & n3017 ;
  assign n3225 = n3223 | n3224 ;
  assign n3226 = n3225 ^ x32 ^ 1'b0 ;
  assign n3227 = n3226 ^ n3217 ^ n2742 ;
  assign n3228 = ( n2742 & n3217 ) | ( n2742 & n3226 ) | ( n3217 & n3226 ) ;
  assign n3229 = x84 & n3025 ;
  assign n3230 = ( x86 & n3015 ) | ( x86 & n3229 ) | ( n3015 & n3229 ) ;
  assign n3231 = n3229 | n3230 ;
  assign n3232 = x85 & ~n3014 ;
  assign n3233 = ( x85 & n3231 ) | ( x85 & ~n3232 ) | ( n3231 & ~n3232 ) ;
  assign n3234 = n1419 & n3017 ;
  assign n3235 = n3233 | n3234 ;
  assign n3236 = n3235 ^ x32 ^ 1'b0 ;
  assign n3237 = ( n2752 & n3228 ) | ( n2752 & n3236 ) | ( n3228 & n3236 ) ;
  assign n3238 = n3236 ^ n3228 ^ n2752 ;
  assign n3239 = x85 & n3025 ;
  assign n3240 = ( x87 & n3015 ) | ( x87 & n3239 ) | ( n3015 & n3239 ) ;
  assign n3241 = n3239 | n3240 ;
  assign n3242 = x86 & ~n3014 ;
  assign n3243 = ( x86 & n3241 ) | ( x86 & ~n3242 ) | ( n3241 & ~n3242 ) ;
  assign n3244 = n1484 & n3017 ;
  assign n3245 = n3243 | n3244 ;
  assign n3246 = n3245 ^ x32 ^ 1'b0 ;
  assign n3247 = n3246 ^ n3237 ^ n2762 ;
  assign n3248 = ( n2762 & n3237 ) | ( n2762 & n3246 ) | ( n3237 & n3246 ) ;
  assign n3249 = x86 & n3025 ;
  assign n3250 = ( x88 & n3015 ) | ( x88 & n3249 ) | ( n3015 & n3249 ) ;
  assign n3251 = n3249 | n3250 ;
  assign n3252 = x87 & ~n3014 ;
  assign n3253 = ( x87 & n3251 ) | ( x87 & ~n3252 ) | ( n3251 & ~n3252 ) ;
  assign n3254 = n1569 & n3017 ;
  assign n3255 = n3253 | n3254 ;
  assign n3256 = n3255 ^ x32 ^ 1'b0 ;
  assign n3257 = ( n2772 & n3248 ) | ( n2772 & n3256 ) | ( n3248 & n3256 ) ;
  assign n3258 = n3256 ^ n3248 ^ n2772 ;
  assign n3259 = x87 & n3025 ;
  assign n3260 = ( x89 & n3015 ) | ( x89 & n3259 ) | ( n3015 & n3259 ) ;
  assign n3261 = n3259 | n3260 ;
  assign n3262 = x88 & ~n3014 ;
  assign n3263 = ( x88 & n3261 ) | ( x88 & ~n3262 ) | ( n3261 & ~n3262 ) ;
  assign n3264 = n1654 & n3017 ;
  assign n3265 = n3263 | n3264 ;
  assign n3266 = n3265 ^ x32 ^ 1'b0 ;
  assign n3267 = n3266 ^ n3257 ^ n2783 ;
  assign n3268 = ( n2783 & n3257 ) | ( n2783 & n3266 ) | ( n3257 & n3266 ) ;
  assign n3269 = x88 & n3025 ;
  assign n3270 = ( x90 & n3015 ) | ( x90 & n3269 ) | ( n3015 & n3269 ) ;
  assign n3271 = n3269 | n3270 ;
  assign n3272 = x89 & ~n3014 ;
  assign n3273 = ( x89 & n3271 ) | ( x89 & ~n3272 ) | ( n3271 & ~n3272 ) ;
  assign n3274 = n1741 & n3017 ;
  assign n3275 = n3273 | n3274 ;
  assign n3276 = n3275 ^ x32 ^ 1'b0 ;
  assign n3277 = ( n2793 & n3268 ) | ( n2793 & n3276 ) | ( n3268 & n3276 ) ;
  assign n3278 = n3276 ^ n3268 ^ n2793 ;
  assign n3279 = x89 & n3025 ;
  assign n3280 = ( x91 & n3015 ) | ( x91 & n3279 ) | ( n3015 & n3279 ) ;
  assign n3281 = n3279 | n3280 ;
  assign n3282 = x90 & ~n3014 ;
  assign n3283 = ( x90 & n3281 ) | ( x90 & ~n3282 ) | ( n3281 & ~n3282 ) ;
  assign n3284 = n2114 & n3017 ;
  assign n3285 = n3283 | n3284 ;
  assign n3286 = n3285 ^ x32 ^ 1'b0 ;
  assign n3287 = ( n2802 & n3277 ) | ( n2802 & n3286 ) | ( n3277 & n3286 ) ;
  assign n3288 = n3286 ^ n3277 ^ n2802 ;
  assign n3289 = x90 & n3025 ;
  assign n3290 = ( x92 & n3015 ) | ( x92 & n3289 ) | ( n3015 & n3289 ) ;
  assign n3291 = n3289 | n3290 ;
  assign n3292 = x91 & ~n3014 ;
  assign n3293 = ( x91 & n3291 ) | ( x91 & ~n3292 ) | ( n3291 & ~n3292 ) ;
  assign n3294 = n2420 & n3017 ;
  assign n3295 = n3293 | n3294 ;
  assign n3296 = n3295 ^ x32 ^ 1'b0 ;
  assign n3297 = n3296 ^ n3287 ^ n2813 ;
  assign n3298 = ( n2813 & n3287 ) | ( n2813 & n3296 ) | ( n3287 & n3296 ) ;
  assign n3299 = x91 & n3025 ;
  assign n3300 = ( x93 & n3015 ) | ( x93 & n3299 ) | ( n3015 & n3299 ) ;
  assign n3301 = n3299 | n3300 ;
  assign n3302 = x92 & ~n3014 ;
  assign n3303 = ( x92 & n3301 ) | ( x92 & ~n3302 ) | ( n3301 & ~n3302 ) ;
  assign n3304 = n2476 & n3017 ;
  assign n3305 = n3303 | n3304 ;
  assign n3306 = n3305 ^ x32 ^ 1'b0 ;
  assign n3307 = ( n2823 & n3298 ) | ( n2823 & n3306 ) | ( n3298 & n3306 ) ;
  assign n3308 = n3306 ^ n3298 ^ n2823 ;
  assign n3309 = x92 & n3025 ;
  assign n3310 = ( x94 & n3015 ) | ( x94 & n3309 ) | ( n3015 & n3309 ) ;
  assign n3311 = n3309 | n3310 ;
  assign n3312 = x93 & ~n3014 ;
  assign n3313 = ( x93 & n3311 ) | ( x93 & ~n3312 ) | ( n3311 & ~n3312 ) ;
  assign n3314 = n2518 & n3017 ;
  assign n3315 = n3313 | n3314 ;
  assign n3316 = n3315 ^ x32 ^ 1'b0 ;
  assign n3317 = n3316 ^ n3307 ^ n2832 ;
  assign n3318 = ( n2832 & n3307 ) | ( n2832 & n3316 ) | ( n3307 & n3316 ) ;
  assign n3319 = x93 & n3025 ;
  assign n3320 = ( x95 & n3015 ) | ( x95 & n3319 ) | ( n3015 & n3319 ) ;
  assign n3321 = n3319 | n3320 ;
  assign n3322 = x94 & ~n3014 ;
  assign n3323 = ( x94 & n3321 ) | ( x94 & ~n3322 ) | ( n3321 & ~n3322 ) ;
  assign n3324 = n2854 & n3017 ;
  assign n3325 = n3323 | n3324 ;
  assign n3326 = n3325 ^ x32 ^ 1'b0 ;
  assign n3327 = n3326 ^ n3318 ^ n2842 ;
  assign n3328 = ( n2842 & n3318 ) | ( n2842 & n3326 ) | ( n3318 & n3326 ) ;
  assign n3329 = x94 & n3025 ;
  assign n3330 = ( x96 & n3015 ) | ( x96 & n3329 ) | ( n3015 & n3329 ) ;
  assign n3331 = n3329 | n3330 ;
  assign n3332 = x95 & ~n3014 ;
  assign n3333 = ( x95 & n3331 ) | ( x95 & ~n3332 ) | ( n3331 & ~n3332 ) ;
  assign n3334 = n2907 & n3017 ;
  assign n3335 = n3333 | n3334 ;
  assign n3336 = n3335 ^ x32 ^ 1'b0 ;
  assign n3337 = ( n2852 & n3328 ) | ( n2852 & n3336 ) | ( n3328 & n3336 ) ;
  assign n3338 = n3336 ^ n3328 ^ n2852 ;
  assign n3339 = x27 ^ x26 ^ 1'b0 ;
  assign n3340 = x29 ^ x28 ^ 1'b0 ;
  assign n3341 = x28 ^ x27 ^ 1'b0 ;
  assign n3342 = n3339 & ~n3340 ;
  assign n3343 = ( ~n3339 & n3340 ) | ( ~n3339 & n3341 ) | ( n3340 & n3341 ) ;
  assign n3344 = ~n3341 & n3343 ;
  assign n3345 = x64 & n3344 ;
  assign n3346 = n3339 & n3340 ;
  assign n3347 = ~n3339 & n3341 ;
  assign n3348 = n139 & n3346 ;
  assign n3349 = x65 & ~n3347 ;
  assign n3350 = x64 & n3339 ;
  assign n3351 = ( x66 & n3342 ) | ( x66 & n3345 ) | ( n3342 & n3345 ) ;
  assign n3352 = n3345 | n3351 ;
  assign n3353 = ( x65 & ~n3349 ) | ( x65 & n3352 ) | ( ~n3349 & n3352 ) ;
  assign n3354 = n3348 | n3353 ;
  assign n3355 = x65 & n3344 ;
  assign n3356 = x64 & n3347 ;
  assign n3357 = ( x67 & n3342 ) | ( x67 & n3355 ) | ( n3342 & n3355 ) ;
  assign n3358 = n3355 | n3357 ;
  assign n3359 = ~x65 & n3342 ;
  assign n3360 = ( n3342 & n3356 ) | ( n3342 & ~n3359 ) | ( n3356 & ~n3359 ) ;
  assign n3361 = x29 & ~n3350 ;
  assign n3362 = ( n190 & n3346 ) | ( n190 & n3356 ) | ( n3346 & n3356 ) ;
  assign n3363 = n3360 | n3362 ;
  assign n3364 = n3363 ^ x29 ^ 1'b0 ;
  assign n3365 = n3364 ^ n3361 ^ 1'b0 ;
  assign n3366 = n3361 & n3364 ;
  assign n3367 = x66 & ~n3347 ;
  assign n3368 = ( x66 & n3358 ) | ( x66 & ~n3367 ) | ( n3358 & ~n3367 ) ;
  assign n3369 = n3354 ^ x29 ^ 1'b0 ;
  assign n3370 = n161 & n3346 ;
  assign n3371 = n3368 | n3370 ;
  assign n3372 = n3366 & n3369 ;
  assign n3373 = n3371 ^ x29 ^ 1'b0 ;
  assign n3374 = n3369 ^ n3366 ^ 1'b0 ;
  assign n3375 = n3373 ^ n3372 ^ n3029 ;
  assign n3376 = ( n3029 & n3372 ) | ( n3029 & n3373 ) | ( n3372 & n3373 ) ;
  assign n3377 = x66 & n3344 ;
  assign n3378 = ( x68 & n3342 ) | ( x68 & n3377 ) | ( n3342 & n3377 ) ;
  assign n3379 = n3377 | n3378 ;
  assign n3380 = x67 & ~n3347 ;
  assign n3381 = ( x67 & n3379 ) | ( x67 & ~n3380 ) | ( n3379 & ~n3380 ) ;
  assign n3382 = n175 & n3346 ;
  assign n3383 = n3381 | n3382 ;
  assign n3384 = n3383 ^ x29 ^ 1'b0 ;
  assign n3385 = n3384 ^ n3376 ^ n3038 ;
  assign n3386 = ( n3038 & n3376 ) | ( n3038 & n3384 ) | ( n3376 & n3384 ) ;
  assign n3387 = x67 & n3344 ;
  assign n3388 = ( x69 & n3342 ) | ( x69 & n3387 ) | ( n3342 & n3387 ) ;
  assign n3389 = n3387 | n3388 ;
  assign n3390 = x68 & ~n3347 ;
  assign n3391 = ( x68 & n3389 ) | ( x68 & ~n3390 ) | ( n3389 & ~n3390 ) ;
  assign n3392 = n172 & n3346 ;
  assign n3393 = n3391 | n3392 ;
  assign n3394 = n3393 ^ x29 ^ 1'b0 ;
  assign n3395 = ( n3036 & n3386 ) | ( n3036 & n3394 ) | ( n3386 & n3394 ) ;
  assign n3396 = n3394 ^ n3386 ^ n3036 ;
  assign n3397 = x68 & n3344 ;
  assign n3398 = ( x70 & n3342 ) | ( x70 & n3397 ) | ( n3342 & n3397 ) ;
  assign n3399 = n3397 | n3398 ;
  assign n3400 = x69 & ~n3347 ;
  assign n3401 = ( x69 & n3399 ) | ( x69 & ~n3400 ) | ( n3399 & ~n3400 ) ;
  assign n3402 = n168 & n3346 ;
  assign n3403 = n3401 | n3402 ;
  assign n3404 = n3403 ^ x29 ^ 1'b0 ;
  assign n3405 = n3404 ^ n3395 ^ n3048 ;
  assign n3406 = ( n3048 & n3395 ) | ( n3048 & n3404 ) | ( n3395 & n3404 ) ;
  assign n3407 = x69 & n3344 ;
  assign n3408 = ( x71 & n3342 ) | ( x71 & n3407 ) | ( n3342 & n3407 ) ;
  assign n3409 = n3407 | n3408 ;
  assign n3410 = x70 & ~n3347 ;
  assign n3411 = ( x70 & n3409 ) | ( x70 & ~n3410 ) | ( n3409 & ~n3410 ) ;
  assign n3412 = n328 & n3346 ;
  assign n3413 = n3411 | n3412 ;
  assign n3414 = n3413 ^ x29 ^ 1'b0 ;
  assign n3415 = n3414 ^ n3406 ^ n3057 ;
  assign n3416 = ( n3057 & n3406 ) | ( n3057 & n3414 ) | ( n3406 & n3414 ) ;
  assign n3417 = x70 & n3344 ;
  assign n3418 = ( x72 & n3342 ) | ( x72 & n3417 ) | ( n3342 & n3417 ) ;
  assign n3419 = n3417 | n3418 ;
  assign n3420 = x71 & ~n3347 ;
  assign n3421 = ( x71 & n3419 ) | ( x71 & ~n3420 ) | ( n3419 & ~n3420 ) ;
  assign n3422 = n349 & n3346 ;
  assign n3423 = n3421 | n3422 ;
  assign n3424 = n3423 ^ x29 ^ 1'b0 ;
  assign n3425 = n3424 ^ n3416 ^ n3067 ;
  assign n3426 = ( n3067 & n3416 ) | ( n3067 & n3424 ) | ( n3416 & n3424 ) ;
  assign n3427 = x71 & n3344 ;
  assign n3428 = ( x73 & n3342 ) | ( x73 & n3427 ) | ( n3342 & n3427 ) ;
  assign n3429 = n3427 | n3428 ;
  assign n3430 = x72 & ~n3347 ;
  assign n3431 = ( x72 & n3429 ) | ( x72 & ~n3430 ) | ( n3429 & ~n3430 ) ;
  assign n3432 = n370 & n3346 ;
  assign n3433 = n3431 | n3432 ;
  assign n3434 = n3433 ^ x29 ^ 1'b0 ;
  assign n3435 = ( n3078 & n3426 ) | ( n3078 & n3434 ) | ( n3426 & n3434 ) ;
  assign n3436 = n3434 ^ n3426 ^ n3078 ;
  assign n3437 = x72 & n3344 ;
  assign n3438 = ( x74 & n3342 ) | ( x74 & n3437 ) | ( n3342 & n3437 ) ;
  assign n3439 = n3437 | n3438 ;
  assign n3440 = x73 & ~n3347 ;
  assign n3441 = ( x73 & n3439 ) | ( x73 & ~n3440 ) | ( n3439 & ~n3440 ) ;
  assign n3442 = n504 & n3346 ;
  assign n3443 = n3441 | n3442 ;
  assign n3444 = n3443 ^ x29 ^ 1'b0 ;
  assign n3445 = ( n3087 & n3435 ) | ( n3087 & n3444 ) | ( n3435 & n3444 ) ;
  assign n3446 = n3444 ^ n3435 ^ n3087 ;
  assign n3447 = x73 & n3344 ;
  assign n3448 = ( x75 & n3342 ) | ( x75 & n3447 ) | ( n3342 & n3447 ) ;
  assign n3449 = n3447 | n3448 ;
  assign n3450 = x74 & ~n3347 ;
  assign n3451 = ( x74 & n3449 ) | ( x74 & ~n3450 ) | ( n3449 & ~n3450 ) ;
  assign n3452 = n525 & n3346 ;
  assign n3453 = n3451 | n3452 ;
  assign n3454 = n3453 ^ x29 ^ 1'b0 ;
  assign n3455 = n3454 ^ n3445 ^ n3098 ;
  assign n3456 = ( n3098 & n3445 ) | ( n3098 & n3454 ) | ( n3445 & n3454 ) ;
  assign n3457 = x74 & n3344 ;
  assign n3458 = ( x76 & n3342 ) | ( x76 & n3457 ) | ( n3342 & n3457 ) ;
  assign n3459 = n3457 | n3458 ;
  assign n3460 = x75 & ~n3347 ;
  assign n3461 = ( x75 & n3459 ) | ( x75 & ~n3460 ) | ( n3459 & ~n3460 ) ;
  assign n3462 = n664 & n3346 ;
  assign n3463 = n3461 | n3462 ;
  assign n3464 = n3463 ^ x29 ^ 1'b0 ;
  assign n3465 = n3464 ^ n3456 ^ n3108 ;
  assign n3466 = ( n3108 & n3456 ) | ( n3108 & n3464 ) | ( n3456 & n3464 ) ;
  assign n3467 = x75 & n3344 ;
  assign n3468 = ( x77 & n3342 ) | ( x77 & n3467 ) | ( n3342 & n3467 ) ;
  assign n3469 = n3467 | n3468 ;
  assign n3470 = x76 & ~n3347 ;
  assign n3471 = ( x76 & n3469 ) | ( x76 & ~n3470 ) | ( n3469 & ~n3470 ) ;
  assign n3472 = n690 & n3346 ;
  assign n3473 = n3471 | n3472 ;
  assign n3474 = n3473 ^ x29 ^ 1'b0 ;
  assign n3475 = ( n3117 & n3466 ) | ( n3117 & n3474 ) | ( n3466 & n3474 ) ;
  assign n3476 = n3474 ^ n3466 ^ n3117 ;
  assign n3477 = x76 & n3344 ;
  assign n3478 = ( x78 & n3342 ) | ( x78 & n3477 ) | ( n3342 & n3477 ) ;
  assign n3479 = n3477 | n3478 ;
  assign n3480 = x77 & ~n3347 ;
  assign n3481 = ( x77 & n3479 ) | ( x77 & ~n3480 ) | ( n3479 & ~n3480 ) ;
  assign n3482 = n709 & n3346 ;
  assign n3483 = n3481 | n3482 ;
  assign n3484 = n3483 ^ x29 ^ 1'b0 ;
  assign n3485 = ( n3128 & n3475 ) | ( n3128 & n3484 ) | ( n3475 & n3484 ) ;
  assign n3486 = n3484 ^ n3475 ^ n3128 ;
  assign n3487 = x77 & n3344 ;
  assign n3488 = ( x79 & n3342 ) | ( x79 & n3487 ) | ( n3342 & n3487 ) ;
  assign n3489 = n3487 | n3488 ;
  assign n3490 = x78 & ~n3347 ;
  assign n3491 = ( x78 & n3489 ) | ( x78 & ~n3490 ) | ( n3489 & ~n3490 ) ;
  assign n3492 = n1015 & n3346 ;
  assign n3493 = n3491 | n3492 ;
  assign n3494 = n3493 ^ x29 ^ 1'b0 ;
  assign n3495 = ( n3137 & n3485 ) | ( n3137 & n3494 ) | ( n3485 & n3494 ) ;
  assign n3496 = n3494 ^ n3485 ^ n3137 ;
  assign n3497 = x78 & n3344 ;
  assign n3498 = ( x80 & n3342 ) | ( x80 & n3497 ) | ( n3342 & n3497 ) ;
  assign n3499 = n3497 | n3498 ;
  assign n3500 = x79 & ~n3347 ;
  assign n3501 = ( x79 & n3499 ) | ( x79 & ~n3500 ) | ( n3499 & ~n3500 ) ;
  assign n3502 = n1216 & n3346 ;
  assign n3503 = n3501 | n3502 ;
  assign n3504 = n3503 ^ x29 ^ 1'b0 ;
  assign n3505 = n3504 ^ n3495 ^ n3148 ;
  assign n3506 = ( n3148 & n3495 ) | ( n3148 & n3504 ) | ( n3495 & n3504 ) ;
  assign n3507 = x79 & n3344 ;
  assign n3508 = ( x81 & n3342 ) | ( x81 & n3507 ) | ( n3342 & n3507 ) ;
  assign n3509 = n3507 | n3508 ;
  assign n3510 = x80 & ~n3347 ;
  assign n3511 = ( x80 & n3509 ) | ( x80 & ~n3510 ) | ( n3509 & ~n3510 ) ;
  assign n3512 = n1258 & n3346 ;
  assign n3513 = n3511 | n3512 ;
  assign n3514 = n3513 ^ x29 ^ 1'b0 ;
  assign n3515 = n3514 ^ n3506 ^ n3157 ;
  assign n3516 = ( n3157 & n3506 ) | ( n3157 & n3514 ) | ( n3506 & n3514 ) ;
  assign n3517 = x80 & n3344 ;
  assign n3518 = ( x82 & n3342 ) | ( x82 & n3517 ) | ( n3342 & n3517 ) ;
  assign n3519 = n3517 | n3518 ;
  assign n3520 = x81 & ~n3347 ;
  assign n3521 = ( x81 & n3519 ) | ( x81 & ~n3520 ) | ( n3519 & ~n3520 ) ;
  assign n3522 = n1301 & n3346 ;
  assign n3523 = n3521 | n3522 ;
  assign n3524 = n3523 ^ x29 ^ 1'b0 ;
  assign n3525 = n3524 ^ n3516 ^ n3167 ;
  assign n3526 = ( n3167 & n3516 ) | ( n3167 & n3524 ) | ( n3516 & n3524 ) ;
  assign n3527 = x81 & n3344 ;
  assign n3528 = ( x83 & n3342 ) | ( x83 & n3527 ) | ( n3342 & n3527 ) ;
  assign n3529 = n3527 | n3528 ;
  assign n3530 = x82 & ~n3347 ;
  assign n3531 = ( x82 & n3529 ) | ( x82 & ~n3530 ) | ( n3529 & ~n3530 ) ;
  assign n3532 = n1329 & n3346 ;
  assign n3533 = n3531 | n3532 ;
  assign n3534 = n3533 ^ x29 ^ 1'b0 ;
  assign n3535 = n3534 ^ n3526 ^ n3177 ;
  assign n3536 = ( n3177 & n3526 ) | ( n3177 & n3534 ) | ( n3526 & n3534 ) ;
  assign n3537 = x82 & n3344 ;
  assign n3538 = ( x84 & n3342 ) | ( x84 & n3537 ) | ( n3342 & n3537 ) ;
  assign n3539 = n3537 | n3538 ;
  assign n3540 = x83 & ~n3347 ;
  assign n3541 = ( x83 & n3539 ) | ( x83 & ~n3540 ) | ( n3539 & ~n3540 ) ;
  assign n3542 = n1355 & n3346 ;
  assign n3543 = n3541 | n3542 ;
  assign n3544 = n3543 ^ x29 ^ 1'b0 ;
  assign n3545 = ( n3187 & n3536 ) | ( n3187 & n3544 ) | ( n3536 & n3544 ) ;
  assign n3546 = n3544 ^ n3536 ^ n3187 ;
  assign n3547 = x83 & n3344 ;
  assign n3548 = ( x85 & n3342 ) | ( x85 & n3547 ) | ( n3342 & n3547 ) ;
  assign n3549 = n3547 | n3548 ;
  assign n3550 = x84 & ~n3347 ;
  assign n3551 = ( x84 & n3549 ) | ( x84 & ~n3550 ) | ( n3549 & ~n3550 ) ;
  assign n3552 = n1392 & n3346 ;
  assign n3553 = n3551 | n3552 ;
  assign n3554 = n3553 ^ x29 ^ 1'b0 ;
  assign n3555 = ( n3197 & n3545 ) | ( n3197 & n3554 ) | ( n3545 & n3554 ) ;
  assign n3556 = n3554 ^ n3545 ^ n3197 ;
  assign n3557 = x84 & n3344 ;
  assign n3558 = ( x86 & n3342 ) | ( x86 & n3557 ) | ( n3342 & n3557 ) ;
  assign n3559 = n3557 | n3558 ;
  assign n3560 = x85 & ~n3347 ;
  assign n3561 = ( x85 & n3559 ) | ( x85 & ~n3560 ) | ( n3559 & ~n3560 ) ;
  assign n3562 = n1419 & n3346 ;
  assign n3563 = n3561 | n3562 ;
  assign n3564 = n3563 ^ x29 ^ 1'b0 ;
  assign n3565 = ( n3208 & n3555 ) | ( n3208 & n3564 ) | ( n3555 & n3564 ) ;
  assign n3566 = n3564 ^ n3555 ^ n3208 ;
  assign n3567 = x85 & n3344 ;
  assign n3568 = ( x87 & n3342 ) | ( x87 & n3567 ) | ( n3342 & n3567 ) ;
  assign n3569 = n3567 | n3568 ;
  assign n3570 = x86 & ~n3347 ;
  assign n3571 = ( x86 & n3569 ) | ( x86 & ~n3570 ) | ( n3569 & ~n3570 ) ;
  assign n3572 = n1484 & n3346 ;
  assign n3573 = n3571 | n3572 ;
  assign n3574 = n3573 ^ x29 ^ 1'b0 ;
  assign n3575 = ( n3218 & n3565 ) | ( n3218 & n3574 ) | ( n3565 & n3574 ) ;
  assign n3576 = n3574 ^ n3565 ^ n3218 ;
  assign n3577 = x86 & n3344 ;
  assign n3578 = ( x88 & n3342 ) | ( x88 & n3577 ) | ( n3342 & n3577 ) ;
  assign n3579 = n3577 | n3578 ;
  assign n3580 = x87 & ~n3347 ;
  assign n3581 = ( x87 & n3579 ) | ( x87 & ~n3580 ) | ( n3579 & ~n3580 ) ;
  assign n3582 = n1569 & n3346 ;
  assign n3583 = n3581 | n3582 ;
  assign n3584 = n3583 ^ x29 ^ 1'b0 ;
  assign n3585 = n3584 ^ n3575 ^ n3227 ;
  assign n3586 = ( n3227 & n3575 ) | ( n3227 & n3584 ) | ( n3575 & n3584 ) ;
  assign n3587 = x87 & n3344 ;
  assign n3588 = ( x89 & n3342 ) | ( x89 & n3587 ) | ( n3342 & n3587 ) ;
  assign n3589 = n3587 | n3588 ;
  assign n3590 = x88 & ~n3347 ;
  assign n3591 = ( x88 & n3589 ) | ( x88 & ~n3590 ) | ( n3589 & ~n3590 ) ;
  assign n3592 = n1654 & n3346 ;
  assign n3593 = n3591 | n3592 ;
  assign n3594 = n3593 ^ x29 ^ 1'b0 ;
  assign n3595 = n3594 ^ n3586 ^ n3238 ;
  assign n3596 = ( n3238 & n3586 ) | ( n3238 & n3594 ) | ( n3586 & n3594 ) ;
  assign n3597 = x88 & n3344 ;
  assign n3598 = ( x90 & n3342 ) | ( x90 & n3597 ) | ( n3342 & n3597 ) ;
  assign n3599 = n3597 | n3598 ;
  assign n3600 = x89 & ~n3347 ;
  assign n3601 = ( x89 & n3599 ) | ( x89 & ~n3600 ) | ( n3599 & ~n3600 ) ;
  assign n3602 = n1741 & n3346 ;
  assign n3603 = n3601 | n3602 ;
  assign n3604 = n3603 ^ x29 ^ 1'b0 ;
  assign n3605 = n3604 ^ n3596 ^ n3247 ;
  assign n3606 = ( n3247 & n3596 ) | ( n3247 & n3604 ) | ( n3596 & n3604 ) ;
  assign n3607 = x89 & n3344 ;
  assign n3608 = ( x91 & n3342 ) | ( x91 & n3607 ) | ( n3342 & n3607 ) ;
  assign n3609 = n3607 | n3608 ;
  assign n3610 = x90 & ~n3347 ;
  assign n3611 = ( x90 & n3609 ) | ( x90 & ~n3610 ) | ( n3609 & ~n3610 ) ;
  assign n3612 = n2114 & n3346 ;
  assign n3613 = n3611 | n3612 ;
  assign n3614 = n3613 ^ x29 ^ 1'b0 ;
  assign n3615 = ( n3258 & n3606 ) | ( n3258 & n3614 ) | ( n3606 & n3614 ) ;
  assign n3616 = n3614 ^ n3606 ^ n3258 ;
  assign n3617 = x90 & n3344 ;
  assign n3618 = ( x92 & n3342 ) | ( x92 & n3617 ) | ( n3342 & n3617 ) ;
  assign n3619 = n3617 | n3618 ;
  assign n3620 = x91 & ~n3347 ;
  assign n3621 = ( x91 & n3619 ) | ( x91 & ~n3620 ) | ( n3619 & ~n3620 ) ;
  assign n3622 = n2420 & n3346 ;
  assign n3623 = n3621 | n3622 ;
  assign n3624 = n3623 ^ x29 ^ 1'b0 ;
  assign n3625 = ( n3267 & n3615 ) | ( n3267 & n3624 ) | ( n3615 & n3624 ) ;
  assign n3626 = n3624 ^ n3615 ^ n3267 ;
  assign n3627 = x91 & n3344 ;
  assign n3628 = ( x93 & n3342 ) | ( x93 & n3627 ) | ( n3342 & n3627 ) ;
  assign n3629 = n3627 | n3628 ;
  assign n3630 = x92 & ~n3347 ;
  assign n3631 = ( x92 & n3629 ) | ( x92 & ~n3630 ) | ( n3629 & ~n3630 ) ;
  assign n3632 = n2476 & n3346 ;
  assign n3633 = n3631 | n3632 ;
  assign n3634 = n3633 ^ x29 ^ 1'b0 ;
  assign n3635 = ( n3278 & n3625 ) | ( n3278 & n3634 ) | ( n3625 & n3634 ) ;
  assign n3636 = n3634 ^ n3625 ^ n3278 ;
  assign n3637 = x94 & ~n3347 ;
  assign n3638 = x93 & n3344 ;
  assign n3639 = ( x95 & n3342 ) | ( x95 & n3638 ) | ( n3342 & n3638 ) ;
  assign n3640 = n3638 | n3639 ;
  assign n3641 = ( x94 & ~n3637 ) | ( x94 & n3640 ) | ( ~n3637 & n3640 ) ;
  assign n3642 = x92 & n3344 ;
  assign n3643 = ( x94 & n3342 ) | ( x94 & n3642 ) | ( n3342 & n3642 ) ;
  assign n3644 = n3642 | n3643 ;
  assign n3645 = x93 & ~n3347 ;
  assign n3646 = ( x93 & n3644 ) | ( x93 & ~n3645 ) | ( n3644 & ~n3645 ) ;
  assign n3647 = n2518 & n3346 ;
  assign n3648 = n3646 | n3647 ;
  assign n3649 = n3648 ^ x29 ^ 1'b0 ;
  assign n3650 = ( n3288 & n3635 ) | ( n3288 & n3649 ) | ( n3635 & n3649 ) ;
  assign n3651 = n3649 ^ n3635 ^ n3288 ;
  assign n3652 = n2854 & n3346 ;
  assign n3653 = x94 & n3344 ;
  assign n3654 = n3641 | n3652 ;
  assign n3655 = n3654 ^ x29 ^ 1'b0 ;
  assign n3656 = n3655 ^ n3650 ^ n3297 ;
  assign n3657 = ( n3297 & n3650 ) | ( n3297 & n3655 ) | ( n3650 & n3655 ) ;
  assign n3658 = ( x96 & n3342 ) | ( x96 & n3653 ) | ( n3342 & n3653 ) ;
  assign n3659 = ( x96 & x97 ) | ( x96 & n2908 ) | ( x97 & n2908 ) ;
  assign n3660 = n3653 | n3658 ;
  assign n3661 = x95 & ~n3347 ;
  assign n3662 = ( x95 & n3660 ) | ( x95 & ~n3661 ) | ( n3660 & ~n3661 ) ;
  assign n3663 = n2907 & n3346 ;
  assign n3664 = n3662 | n3663 ;
  assign n3665 = n3664 ^ x29 ^ 1'b0 ;
  assign n3666 = n3665 ^ n3657 ^ n3308 ;
  assign n3667 = ( n3308 & n3657 ) | ( n3308 & n3665 ) | ( n3657 & n3665 ) ;
  assign n3668 = n2908 ^ x97 ^ x96 ;
  assign n3669 = x95 & n3344 ;
  assign n3670 = ( x97 & n3342 ) | ( x97 & n3669 ) | ( n3342 & n3669 ) ;
  assign n3671 = n3669 | n3670 ;
  assign n3672 = x96 & ~n3347 ;
  assign n3673 = ( x96 & n3671 ) | ( x96 & ~n3672 ) | ( n3671 & ~n3672 ) ;
  assign n3674 = n3346 & n3668 ;
  assign n3675 = n3673 | n3674 ;
  assign n3676 = n3675 ^ x29 ^ 1'b0 ;
  assign n3677 = ( n3317 & n3667 ) | ( n3317 & n3676 ) | ( n3667 & n3676 ) ;
  assign n3678 = n3676 ^ n3667 ^ n3317 ;
  assign n3679 = x95 & n888 ;
  assign n3680 = ( x97 & n878 ) | ( x97 & n3679 ) | ( n878 & n3679 ) ;
  assign n3681 = n3679 | n3680 ;
  assign n3682 = x96 & ~n877 ;
  assign n3683 = ( x96 & n3681 ) | ( x96 & ~n3682 ) | ( n3681 & ~n3682 ) ;
  assign n3684 = n880 & n3668 ;
  assign n3685 = n3683 | n3684 ;
  assign n3686 = n3685 ^ x44 ^ 1'b0 ;
  assign n3687 = ( n2535 & n2946 ) | ( n2535 & n3686 ) | ( n2946 & n3686 ) ;
  assign n3688 = n3686 ^ n2946 ^ n2535 ;
  assign n3689 = x95 & n2560 ;
  assign n3690 = ( x97 & n2567 ) | ( x97 & n3689 ) | ( n2567 & n3689 ) ;
  assign n3691 = n3689 | n3690 ;
  assign n3692 = x96 & ~n2562 ;
  assign n3693 = ( x96 & n3691 ) | ( x96 & ~n3692 ) | ( n3691 & ~n3692 ) ;
  assign n3694 = n2565 & n3668 ;
  assign n3695 = n3693 | n3694 ;
  assign n3696 = n3695 ^ x35 ^ 1'b0 ;
  assign n3697 = ( n2502 & n2545 ) | ( n2502 & n3696 ) | ( n2545 & n3696 ) ;
  assign n3698 = n3696 ^ n2545 ^ n2502 ;
  assign n3699 = x95 & n1058 ;
  assign n3700 = ( x97 & n1065 ) | ( x97 & n3699 ) | ( n1065 & n3699 ) ;
  assign n3701 = n3699 | n3700 ;
  assign n3702 = x96 & ~n1060 ;
  assign n3703 = ( x96 & n3701 ) | ( x96 & ~n3702 ) | ( n3701 & ~n3702 ) ;
  assign n3704 = n1063 & n3668 ;
  assign n3705 = n3703 | n3704 ;
  assign n3706 = n3705 ^ x41 ^ 1'b0 ;
  assign n3707 = n3706 ^ n2916 ^ n2524 ;
  assign n3708 = ( n2524 & n2916 ) | ( n2524 & n3706 ) | ( n2916 & n3706 ) ;
  assign n3709 = x95 & n3025 ;
  assign n3710 = ( x97 & n3015 ) | ( x97 & n3709 ) | ( n3015 & n3709 ) ;
  assign n3711 = n3709 | n3710 ;
  assign n3712 = x96 & ~n3014 ;
  assign n3713 = ( x96 & n3711 ) | ( x96 & ~n3712 ) | ( n3711 & ~n3712 ) ;
  assign n3714 = n3017 & n3668 ;
  assign n3715 = n3713 | n3714 ;
  assign n3716 = n3715 ^ x32 ^ 1'b0 ;
  assign n3717 = n3716 ^ n3337 ^ n2885 ;
  assign n3718 = ( n2885 & n3337 ) | ( n2885 & n3716 ) | ( n3337 & n3716 ) ;
  assign n3719 = x95 & n2156 ;
  assign n3720 = ( x97 & n2163 ) | ( x97 & n3719 ) | ( n2163 & n3719 ) ;
  assign n3721 = n3719 | n3720 ;
  assign n3722 = x96 & ~n2158 ;
  assign n3723 = ( x96 & n3721 ) | ( x96 & ~n3722 ) | ( n3721 & ~n3722 ) ;
  assign n3724 = n2161 & n3668 ;
  assign n3725 = n3723 | n3724 ;
  assign n3726 = n3725 ^ x38 ^ 1'b0 ;
  assign n3727 = n3726 ^ n2936 ^ n2554 ;
  assign n3728 = ( n2554 & n2936 ) | ( n2554 & n3726 ) | ( n2936 & n3726 ) ;
  assign n3729 = x24 ^ x23 ^ 1'b0 ;
  assign n3730 = x26 ^ x25 ^ 1'b0 ;
  assign n3731 = x25 ^ x24 ^ 1'b0 ;
  assign n3732 = n3729 & ~n3730 ;
  assign n3733 = ( ~n3729 & n3730 ) | ( ~n3729 & n3731 ) | ( n3730 & n3731 ) ;
  assign n3734 = ~n3731 & n3733 ;
  assign n3735 = x64 & n3734 ;
  assign n3736 = n3729 & n3730 ;
  assign n3737 = ~n3729 & n3731 ;
  assign n3738 = n139 & n3736 ;
  assign n3739 = x65 & ~n3737 ;
  assign n3740 = x64 & n3729 ;
  assign n3741 = ( x66 & n3732 ) | ( x66 & n3735 ) | ( n3732 & n3735 ) ;
  assign n3742 = n3735 | n3741 ;
  assign n3743 = ( x65 & ~n3739 ) | ( x65 & n3742 ) | ( ~n3739 & n3742 ) ;
  assign n3744 = n3738 | n3743 ;
  assign n3745 = x65 & n3734 ;
  assign n3746 = x64 & n3737 ;
  assign n3747 = ( x67 & n3732 ) | ( x67 & n3745 ) | ( n3732 & n3745 ) ;
  assign n3748 = n3745 | n3747 ;
  assign n3749 = ~x65 & n3732 ;
  assign n3750 = ( n3732 & n3746 ) | ( n3732 & ~n3749 ) | ( n3746 & ~n3749 ) ;
  assign n3751 = x26 & ~n3740 ;
  assign n3752 = ( n190 & n3736 ) | ( n190 & n3746 ) | ( n3736 & n3746 ) ;
  assign n3753 = n3750 | n3752 ;
  assign n3754 = n3753 ^ x26 ^ 1'b0 ;
  assign n3755 = n3754 ^ n3751 ^ 1'b0 ;
  assign n3756 = n3751 & n3754 ;
  assign n3757 = x66 & ~n3737 ;
  assign n3758 = ( x66 & n3748 ) | ( x66 & ~n3757 ) | ( n3748 & ~n3757 ) ;
  assign n3759 = n3744 ^ x26 ^ 1'b0 ;
  assign n3760 = n161 & n3736 ;
  assign n3761 = n3758 | n3760 ;
  assign n3762 = n3756 & n3759 ;
  assign n3763 = n3761 ^ x26 ^ 1'b0 ;
  assign n3764 = n3759 ^ n3756 ^ 1'b0 ;
  assign n3765 = n3763 ^ n3762 ^ n3350 ;
  assign n3766 = ( n3350 & n3762 ) | ( n3350 & n3763 ) | ( n3762 & n3763 ) ;
  assign n3767 = x66 & n3734 ;
  assign n3768 = ( x68 & n3732 ) | ( x68 & n3767 ) | ( n3732 & n3767 ) ;
  assign n3769 = n3767 | n3768 ;
  assign n3770 = x67 & ~n3737 ;
  assign n3771 = ( x67 & n3769 ) | ( x67 & ~n3770 ) | ( n3769 & ~n3770 ) ;
  assign n3772 = n175 & n3736 ;
  assign n3773 = n3771 | n3772 ;
  assign n3774 = n3773 ^ x26 ^ 1'b0 ;
  assign n3775 = n3774 ^ n3766 ^ n3365 ;
  assign n3776 = ( n3365 & n3766 ) | ( n3365 & n3774 ) | ( n3766 & n3774 ) ;
  assign n3777 = x67 & n3734 ;
  assign n3778 = ( x69 & n3732 ) | ( x69 & n3777 ) | ( n3732 & n3777 ) ;
  assign n3779 = n3777 | n3778 ;
  assign n3780 = x68 & ~n3737 ;
  assign n3781 = ( x68 & n3779 ) | ( x68 & ~n3780 ) | ( n3779 & ~n3780 ) ;
  assign n3782 = n172 & n3736 ;
  assign n3783 = n3781 | n3782 ;
  assign n3784 = n3783 ^ x26 ^ 1'b0 ;
  assign n3785 = ( n3374 & n3776 ) | ( n3374 & n3784 ) | ( n3776 & n3784 ) ;
  assign n3786 = n3784 ^ n3776 ^ n3374 ;
  assign n3787 = x68 & n3734 ;
  assign n3788 = ( x70 & n3732 ) | ( x70 & n3787 ) | ( n3732 & n3787 ) ;
  assign n3789 = n3787 | n3788 ;
  assign n3790 = x69 & ~n3737 ;
  assign n3791 = ( x69 & n3789 ) | ( x69 & ~n3790 ) | ( n3789 & ~n3790 ) ;
  assign n3792 = n168 & n3736 ;
  assign n3793 = n3791 | n3792 ;
  assign n3794 = n3793 ^ x26 ^ 1'b0 ;
  assign n3795 = ( n3375 & n3785 ) | ( n3375 & n3794 ) | ( n3785 & n3794 ) ;
  assign n3796 = n3794 ^ n3785 ^ n3375 ;
  assign n3797 = x69 & n3734 ;
  assign n3798 = ( x71 & n3732 ) | ( x71 & n3797 ) | ( n3732 & n3797 ) ;
  assign n3799 = n3797 | n3798 ;
  assign n3800 = x70 & ~n3737 ;
  assign n3801 = ( x70 & n3799 ) | ( x70 & ~n3800 ) | ( n3799 & ~n3800 ) ;
  assign n3802 = n328 & n3736 ;
  assign n3803 = n3801 | n3802 ;
  assign n3804 = n3803 ^ x26 ^ 1'b0 ;
  assign n3805 = ( n3385 & n3795 ) | ( n3385 & n3804 ) | ( n3795 & n3804 ) ;
  assign n3806 = n3804 ^ n3795 ^ n3385 ;
  assign n3807 = x70 & n3734 ;
  assign n3808 = ( x72 & n3732 ) | ( x72 & n3807 ) | ( n3732 & n3807 ) ;
  assign n3809 = n3807 | n3808 ;
  assign n3810 = x71 & ~n3737 ;
  assign n3811 = ( x71 & n3809 ) | ( x71 & ~n3810 ) | ( n3809 & ~n3810 ) ;
  assign n3812 = n349 & n3736 ;
  assign n3813 = n3811 | n3812 ;
  assign n3814 = n3813 ^ x26 ^ 1'b0 ;
  assign n3815 = n3814 ^ n3805 ^ n3396 ;
  assign n3816 = ( n3396 & n3805 ) | ( n3396 & n3814 ) | ( n3805 & n3814 ) ;
  assign n3817 = x71 & n3734 ;
  assign n3818 = ( x73 & n3732 ) | ( x73 & n3817 ) | ( n3732 & n3817 ) ;
  assign n3819 = n3817 | n3818 ;
  assign n3820 = x72 & ~n3737 ;
  assign n3821 = ( x72 & n3819 ) | ( x72 & ~n3820 ) | ( n3819 & ~n3820 ) ;
  assign n3822 = n370 & n3736 ;
  assign n3823 = n3821 | n3822 ;
  assign n3824 = n3823 ^ x26 ^ 1'b0 ;
  assign n3825 = n3824 ^ n3816 ^ n3405 ;
  assign n3826 = ( n3405 & n3816 ) | ( n3405 & n3824 ) | ( n3816 & n3824 ) ;
  assign n3827 = x72 & n3734 ;
  assign n3828 = ( x74 & n3732 ) | ( x74 & n3827 ) | ( n3732 & n3827 ) ;
  assign n3829 = n3827 | n3828 ;
  assign n3830 = x73 & ~n3737 ;
  assign n3831 = ( x73 & n3829 ) | ( x73 & ~n3830 ) | ( n3829 & ~n3830 ) ;
  assign n3832 = n504 & n3736 ;
  assign n3833 = n3831 | n3832 ;
  assign n3834 = n3833 ^ x26 ^ 1'b0 ;
  assign n3835 = n3834 ^ n3826 ^ n3415 ;
  assign n3836 = ( n3415 & n3826 ) | ( n3415 & n3834 ) | ( n3826 & n3834 ) ;
  assign n3837 = x73 & n3734 ;
  assign n3838 = ( x75 & n3732 ) | ( x75 & n3837 ) | ( n3732 & n3837 ) ;
  assign n3839 = n3837 | n3838 ;
  assign n3840 = x74 & ~n3737 ;
  assign n3841 = ( x74 & n3839 ) | ( x74 & ~n3840 ) | ( n3839 & ~n3840 ) ;
  assign n3842 = n525 & n3736 ;
  assign n3843 = n3841 | n3842 ;
  assign n3844 = n3843 ^ x26 ^ 1'b0 ;
  assign n3845 = ( n3425 & n3836 ) | ( n3425 & n3844 ) | ( n3836 & n3844 ) ;
  assign n3846 = n3844 ^ n3836 ^ n3425 ;
  assign n3847 = x74 & n3734 ;
  assign n3848 = ( x76 & n3732 ) | ( x76 & n3847 ) | ( n3732 & n3847 ) ;
  assign n3849 = n3847 | n3848 ;
  assign n3850 = x75 & ~n3737 ;
  assign n3851 = ( x75 & n3849 ) | ( x75 & ~n3850 ) | ( n3849 & ~n3850 ) ;
  assign n3852 = n664 & n3736 ;
  assign n3853 = n3851 | n3852 ;
  assign n3854 = n3853 ^ x26 ^ 1'b0 ;
  assign n3855 = ( n3436 & n3845 ) | ( n3436 & n3854 ) | ( n3845 & n3854 ) ;
  assign n3856 = n3854 ^ n3845 ^ n3436 ;
  assign n3857 = x75 & n3734 ;
  assign n3858 = ( x77 & n3732 ) | ( x77 & n3857 ) | ( n3732 & n3857 ) ;
  assign n3859 = n3857 | n3858 ;
  assign n3860 = x76 & ~n3737 ;
  assign n3861 = ( x76 & n3859 ) | ( x76 & ~n3860 ) | ( n3859 & ~n3860 ) ;
  assign n3862 = n690 & n3736 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = n3863 ^ x26 ^ 1'b0 ;
  assign n3865 = ( n3446 & n3855 ) | ( n3446 & n3864 ) | ( n3855 & n3864 ) ;
  assign n3866 = n3864 ^ n3855 ^ n3446 ;
  assign n3867 = x76 & n3734 ;
  assign n3868 = ( x78 & n3732 ) | ( x78 & n3867 ) | ( n3732 & n3867 ) ;
  assign n3869 = n3867 | n3868 ;
  assign n3870 = x77 & ~n3737 ;
  assign n3871 = ( x77 & n3869 ) | ( x77 & ~n3870 ) | ( n3869 & ~n3870 ) ;
  assign n3872 = n709 & n3736 ;
  assign n3873 = n3871 | n3872 ;
  assign n3874 = n3873 ^ x26 ^ 1'b0 ;
  assign n3875 = ( n3455 & n3865 ) | ( n3455 & n3874 ) | ( n3865 & n3874 ) ;
  assign n3876 = n3874 ^ n3865 ^ n3455 ;
  assign n3877 = x77 & n3734 ;
  assign n3878 = ( x79 & n3732 ) | ( x79 & n3877 ) | ( n3732 & n3877 ) ;
  assign n3879 = n3877 | n3878 ;
  assign n3880 = x78 & ~n3737 ;
  assign n3881 = ( x78 & n3879 ) | ( x78 & ~n3880 ) | ( n3879 & ~n3880 ) ;
  assign n3882 = n1015 & n3736 ;
  assign n3883 = n3881 | n3882 ;
  assign n3884 = n3883 ^ x26 ^ 1'b0 ;
  assign n3885 = n3884 ^ n3875 ^ n3465 ;
  assign n3886 = ( n3465 & n3875 ) | ( n3465 & n3884 ) | ( n3875 & n3884 ) ;
  assign n3887 = x78 & n3734 ;
  assign n3888 = ( x80 & n3732 ) | ( x80 & n3887 ) | ( n3732 & n3887 ) ;
  assign n3889 = n3887 | n3888 ;
  assign n3890 = x79 & ~n3737 ;
  assign n3891 = ( x79 & n3889 ) | ( x79 & ~n3890 ) | ( n3889 & ~n3890 ) ;
  assign n3892 = n1216 & n3736 ;
  assign n3893 = n3891 | n3892 ;
  assign n3894 = n3893 ^ x26 ^ 1'b0 ;
  assign n3895 = ( n3476 & n3886 ) | ( n3476 & n3894 ) | ( n3886 & n3894 ) ;
  assign n3896 = n3894 ^ n3886 ^ n3476 ;
  assign n3897 = x79 & n3734 ;
  assign n3898 = ( x81 & n3732 ) | ( x81 & n3897 ) | ( n3732 & n3897 ) ;
  assign n3899 = n3897 | n3898 ;
  assign n3900 = x80 & ~n3737 ;
  assign n3901 = ( x80 & n3899 ) | ( x80 & ~n3900 ) | ( n3899 & ~n3900 ) ;
  assign n3902 = n1258 & n3736 ;
  assign n3903 = n3901 | n3902 ;
  assign n3904 = n3903 ^ x26 ^ 1'b0 ;
  assign n3905 = ( n3486 & n3895 ) | ( n3486 & n3904 ) | ( n3895 & n3904 ) ;
  assign n3906 = n3904 ^ n3895 ^ n3486 ;
  assign n3907 = x80 & n3734 ;
  assign n3908 = ( x82 & n3732 ) | ( x82 & n3907 ) | ( n3732 & n3907 ) ;
  assign n3909 = n3907 | n3908 ;
  assign n3910 = x81 & ~n3737 ;
  assign n3911 = ( x81 & n3909 ) | ( x81 & ~n3910 ) | ( n3909 & ~n3910 ) ;
  assign n3912 = n1301 & n3736 ;
  assign n3913 = n3911 | n3912 ;
  assign n3914 = n3913 ^ x26 ^ 1'b0 ;
  assign n3915 = n3914 ^ n3905 ^ n3496 ;
  assign n3916 = ( n3496 & n3905 ) | ( n3496 & n3914 ) | ( n3905 & n3914 ) ;
  assign n3917 = x81 & n3734 ;
  assign n3918 = ( x83 & n3732 ) | ( x83 & n3917 ) | ( n3732 & n3917 ) ;
  assign n3919 = n3917 | n3918 ;
  assign n3920 = x82 & ~n3737 ;
  assign n3921 = ( x82 & n3919 ) | ( x82 & ~n3920 ) | ( n3919 & ~n3920 ) ;
  assign n3922 = n1329 & n3736 ;
  assign n3923 = n3921 | n3922 ;
  assign n3924 = n3923 ^ x26 ^ 1'b0 ;
  assign n3925 = ( n3505 & n3916 ) | ( n3505 & n3924 ) | ( n3916 & n3924 ) ;
  assign n3926 = n3924 ^ n3916 ^ n3505 ;
  assign n3927 = x82 & n3734 ;
  assign n3928 = ( x84 & n3732 ) | ( x84 & n3927 ) | ( n3732 & n3927 ) ;
  assign n3929 = n3927 | n3928 ;
  assign n3930 = x83 & ~n3737 ;
  assign n3931 = ( x83 & n3929 ) | ( x83 & ~n3930 ) | ( n3929 & ~n3930 ) ;
  assign n3932 = n1355 & n3736 ;
  assign n3933 = n3931 | n3932 ;
  assign n3934 = n3933 ^ x26 ^ 1'b0 ;
  assign n3935 = ( n3515 & n3925 ) | ( n3515 & n3934 ) | ( n3925 & n3934 ) ;
  assign n3936 = n3934 ^ n3925 ^ n3515 ;
  assign n3937 = x83 & n3734 ;
  assign n3938 = ( x85 & n3732 ) | ( x85 & n3937 ) | ( n3732 & n3937 ) ;
  assign n3939 = n3937 | n3938 ;
  assign n3940 = x84 & ~n3737 ;
  assign n3941 = ( x84 & n3939 ) | ( x84 & ~n3940 ) | ( n3939 & ~n3940 ) ;
  assign n3942 = n1392 & n3736 ;
  assign n3943 = n3941 | n3942 ;
  assign n3944 = n3943 ^ x26 ^ 1'b0 ;
  assign n3945 = ( n3525 & n3935 ) | ( n3525 & n3944 ) | ( n3935 & n3944 ) ;
  assign n3946 = n3944 ^ n3935 ^ n3525 ;
  assign n3947 = x84 & n3734 ;
  assign n3948 = ( x86 & n3732 ) | ( x86 & n3947 ) | ( n3732 & n3947 ) ;
  assign n3949 = n3947 | n3948 ;
  assign n3950 = x85 & ~n3737 ;
  assign n3951 = ( x85 & n3949 ) | ( x85 & ~n3950 ) | ( n3949 & ~n3950 ) ;
  assign n3952 = n1419 & n3736 ;
  assign n3953 = n3951 | n3952 ;
  assign n3954 = n3953 ^ x26 ^ 1'b0 ;
  assign n3955 = n3954 ^ n3945 ^ n3535 ;
  assign n3956 = ( n3535 & n3945 ) | ( n3535 & n3954 ) | ( n3945 & n3954 ) ;
  assign n3957 = x85 & n3734 ;
  assign n3958 = ( x87 & n3732 ) | ( x87 & n3957 ) | ( n3732 & n3957 ) ;
  assign n3959 = n3957 | n3958 ;
  assign n3960 = x86 & ~n3737 ;
  assign n3961 = ( x86 & n3959 ) | ( x86 & ~n3960 ) | ( n3959 & ~n3960 ) ;
  assign n3962 = n1484 & n3736 ;
  assign n3963 = n3961 | n3962 ;
  assign n3964 = n3963 ^ x26 ^ 1'b0 ;
  assign n3965 = n3964 ^ n3956 ^ n3546 ;
  assign n3966 = ( n3546 & n3956 ) | ( n3546 & n3964 ) | ( n3956 & n3964 ) ;
  assign n3967 = x86 & n3734 ;
  assign n3968 = ( x88 & n3732 ) | ( x88 & n3967 ) | ( n3732 & n3967 ) ;
  assign n3969 = n3967 | n3968 ;
  assign n3970 = x87 & ~n3737 ;
  assign n3971 = ( x87 & n3969 ) | ( x87 & ~n3970 ) | ( n3969 & ~n3970 ) ;
  assign n3972 = n1569 & n3736 ;
  assign n3973 = n3971 | n3972 ;
  assign n3974 = n3973 ^ x26 ^ 1'b0 ;
  assign n3975 = n3974 ^ n3966 ^ n3556 ;
  assign n3976 = ( n3556 & n3966 ) | ( n3556 & n3974 ) | ( n3966 & n3974 ) ;
  assign n3977 = x87 & n3734 ;
  assign n3978 = ( x89 & n3732 ) | ( x89 & n3977 ) | ( n3732 & n3977 ) ;
  assign n3979 = n3977 | n3978 ;
  assign n3980 = x88 & ~n3737 ;
  assign n3981 = ( x88 & n3979 ) | ( x88 & ~n3980 ) | ( n3979 & ~n3980 ) ;
  assign n3982 = n1654 & n3736 ;
  assign n3983 = n3981 | n3982 ;
  assign n3984 = n3983 ^ x26 ^ 1'b0 ;
  assign n3985 = ( n3566 & n3976 ) | ( n3566 & n3984 ) | ( n3976 & n3984 ) ;
  assign n3986 = n3984 ^ n3976 ^ n3566 ;
  assign n3987 = x88 & n3734 ;
  assign n3988 = ( x90 & n3732 ) | ( x90 & n3987 ) | ( n3732 & n3987 ) ;
  assign n3989 = n3987 | n3988 ;
  assign n3990 = x89 & ~n3737 ;
  assign n3991 = ( x89 & n3989 ) | ( x89 & ~n3990 ) | ( n3989 & ~n3990 ) ;
  assign n3992 = n1741 & n3736 ;
  assign n3993 = n3991 | n3992 ;
  assign n3994 = n3993 ^ x26 ^ 1'b0 ;
  assign n3995 = n3994 ^ n3985 ^ n3576 ;
  assign n3996 = ( n3576 & n3985 ) | ( n3576 & n3994 ) | ( n3985 & n3994 ) ;
  assign n3997 = x89 & n3734 ;
  assign n3998 = ( x91 & n3732 ) | ( x91 & n3997 ) | ( n3732 & n3997 ) ;
  assign n3999 = n3997 | n3998 ;
  assign n4000 = x90 & ~n3737 ;
  assign n4001 = ( x90 & n3999 ) | ( x90 & ~n4000 ) | ( n3999 & ~n4000 ) ;
  assign n4002 = n2114 & n3736 ;
  assign n4003 = n4001 | n4002 ;
  assign n4004 = n4003 ^ x26 ^ 1'b0 ;
  assign n4005 = n4004 ^ n3996 ^ n3585 ;
  assign n4006 = ( n3585 & n3996 ) | ( n3585 & n4004 ) | ( n3996 & n4004 ) ;
  assign n4007 = x90 & n3734 ;
  assign n4008 = ( x92 & n3732 ) | ( x92 & n4007 ) | ( n3732 & n4007 ) ;
  assign n4009 = n4007 | n4008 ;
  assign n4010 = x91 & ~n3737 ;
  assign n4011 = ( x91 & n4009 ) | ( x91 & ~n4010 ) | ( n4009 & ~n4010 ) ;
  assign n4012 = n2420 & n3736 ;
  assign n4013 = n4011 | n4012 ;
  assign n4014 = n4013 ^ x26 ^ 1'b0 ;
  assign n4015 = ( n3595 & n4006 ) | ( n3595 & n4014 ) | ( n4006 & n4014 ) ;
  assign n4016 = n4014 ^ n4006 ^ n3595 ;
  assign n4017 = x91 & n3734 ;
  assign n4018 = ( x93 & n3732 ) | ( x93 & n4017 ) | ( n3732 & n4017 ) ;
  assign n4019 = n4017 | n4018 ;
  assign n4020 = x92 & ~n3737 ;
  assign n4021 = ( x92 & n4019 ) | ( x92 & ~n4020 ) | ( n4019 & ~n4020 ) ;
  assign n4022 = n2476 & n3736 ;
  assign n4023 = n4021 | n4022 ;
  assign n4024 = n4023 ^ x26 ^ 1'b0 ;
  assign n4025 = n4024 ^ n4015 ^ n3605 ;
  assign n4026 = ( n3605 & n4015 ) | ( n3605 & n4024 ) | ( n4015 & n4024 ) ;
  assign n4027 = x92 & n3734 ;
  assign n4028 = ( x94 & n3732 ) | ( x94 & n4027 ) | ( n3732 & n4027 ) ;
  assign n4029 = n4027 | n4028 ;
  assign n4030 = x93 & ~n3737 ;
  assign n4031 = ( x93 & n4029 ) | ( x93 & ~n4030 ) | ( n4029 & ~n4030 ) ;
  assign n4032 = n2518 & n3736 ;
  assign n4033 = n4031 | n4032 ;
  assign n4034 = n4033 ^ x26 ^ 1'b0 ;
  assign n4035 = ( n3616 & n4026 ) | ( n3616 & n4034 ) | ( n4026 & n4034 ) ;
  assign n4036 = n4034 ^ n4026 ^ n3616 ;
  assign n4037 = x96 & n888 ;
  assign n4038 = ( x98 & n878 ) | ( x98 & n4037 ) | ( n878 & n4037 ) ;
  assign n4039 = n4037 | n4038 ;
  assign n4040 = x93 & n3734 ;
  assign n4041 = x97 & ~n877 ;
  assign n4042 = ( x97 & n4039 ) | ( x97 & ~n4041 ) | ( n4039 & ~n4041 ) ;
  assign n4043 = ( x95 & n3732 ) | ( x95 & n4040 ) | ( n3732 & n4040 ) ;
  assign n4044 = n4040 | n4043 ;
  assign n4045 = x94 & ~n3737 ;
  assign n4046 = ( x94 & n4044 ) | ( x94 & ~n4045 ) | ( n4044 & ~n4045 ) ;
  assign n4047 = n2854 & n3736 ;
  assign n4048 = n4046 | n4047 ;
  assign n4049 = n4048 ^ x26 ^ 1'b0 ;
  assign n4050 = ( n3626 & n4035 ) | ( n3626 & n4049 ) | ( n4035 & n4049 ) ;
  assign n4051 = n4049 ^ n4035 ^ n3626 ;
  assign n4052 = n3659 ^ x98 ^ x97 ;
  assign n4053 = n880 & n4052 ;
  assign n4054 = n4042 | n4053 ;
  assign n4055 = n4054 ^ x44 ^ 1'b0 ;
  assign n4056 = n4055 ^ n3010 ^ n2534 ;
  assign n4057 = ( n2534 & n3010 ) | ( n2534 & n4055 ) | ( n3010 & n4055 ) ;
  assign n4058 = x94 & n3734 ;
  assign n4059 = ( x96 & n3732 ) | ( x96 & n4058 ) | ( n3732 & n4058 ) ;
  assign n4060 = n4058 | n4059 ;
  assign n4061 = x95 & ~n3737 ;
  assign n4062 = ( x95 & n4060 ) | ( x95 & ~n4061 ) | ( n4060 & ~n4061 ) ;
  assign n4063 = n2907 & n3736 ;
  assign n4064 = n4062 | n4063 ;
  assign n4065 = n4064 ^ x26 ^ 1'b0 ;
  assign n4066 = n4065 ^ n4050 ^ n3636 ;
  assign n4067 = ( n3636 & n4050 ) | ( n3636 & n4065 ) | ( n4050 & n4065 ) ;
  assign n4068 = x95 & n3734 ;
  assign n4069 = ( x97 & n3732 ) | ( x97 & n4068 ) | ( n3732 & n4068 ) ;
  assign n4070 = n4068 | n4069 ;
  assign n4071 = x96 & ~n3737 ;
  assign n4072 = ( x96 & n4070 ) | ( x96 & ~n4071 ) | ( n4070 & ~n4071 ) ;
  assign n4073 = n3668 & n3736 ;
  assign n4074 = n4072 | n4073 ;
  assign n4075 = n4074 ^ x26 ^ 1'b0 ;
  assign n4076 = n4075 ^ n4067 ^ n3651 ;
  assign n4077 = ( n3651 & n4067 ) | ( n3651 & n4075 ) | ( n4067 & n4075 ) ;
  assign n4078 = x96 & n3734 ;
  assign n4079 = ( x98 & n3732 ) | ( x98 & n4078 ) | ( n3732 & n4078 ) ;
  assign n4080 = ( x97 & x98 ) | ( x97 & n3659 ) | ( x98 & n3659 ) ;
  assign n4081 = n4078 | n4079 ;
  assign n4082 = x97 & ~n3737 ;
  assign n4083 = ( x97 & n4081 ) | ( x97 & ~n4082 ) | ( n4081 & ~n4082 ) ;
  assign n4084 = n3736 & n4052 ;
  assign n4085 = n4083 | n4084 ;
  assign n4086 = n4085 ^ x26 ^ 1'b0 ;
  assign n4087 = n4086 ^ n4077 ^ n3656 ;
  assign n4088 = ( n3656 & n4077 ) | ( n3656 & n4086 ) | ( n4077 & n4086 ) ;
  assign n4089 = x96 & n1058 ;
  assign n4090 = ( x98 & n1065 ) | ( x98 & n4089 ) | ( n1065 & n4089 ) ;
  assign n4091 = n4089 | n4090 ;
  assign n4092 = x97 & ~n1060 ;
  assign n4093 = ( x97 & n4091 ) | ( x97 & ~n4092 ) | ( n4091 & ~n4092 ) ;
  assign n4094 = n1063 & n4052 ;
  assign n4095 = n4093 | n4094 ;
  assign n4096 = n4095 ^ x41 ^ 1'b0 ;
  assign n4097 = ( n2523 & n2894 ) | ( n2523 & n4096 ) | ( n2894 & n4096 ) ;
  assign n4098 = n4096 ^ n2894 ^ n2523 ;
  assign n4099 = x96 & n3025 ;
  assign n4100 = ( x98 & n3015 ) | ( x98 & n4099 ) | ( n3015 & n4099 ) ;
  assign n4101 = n4099 | n4100 ;
  assign n4102 = x97 & ~n3014 ;
  assign n4103 = ( x97 & n4101 ) | ( x97 & ~n4102 ) | ( n4101 & ~n4102 ) ;
  assign n4104 = n3017 & n4052 ;
  assign n4105 = n4103 | n4104 ;
  assign n4106 = n4105 ^ x32 ^ 1'b0 ;
  assign n4107 = ( n2905 & n3718 ) | ( n2905 & n4106 ) | ( n3718 & n4106 ) ;
  assign n4108 = n4106 ^ n3718 ^ n2905 ;
  assign n4109 = x96 & n2156 ;
  assign n4110 = ( x98 & n2163 ) | ( x98 & n4109 ) | ( n2163 & n4109 ) ;
  assign n4111 = n4109 | n4110 ;
  assign n4112 = x97 & ~n2158 ;
  assign n4113 = ( x97 & n4111 ) | ( x97 & ~n4112 ) | ( n4111 & ~n4112 ) ;
  assign n4114 = n2161 & n4052 ;
  assign n4115 = n4113 | n4114 ;
  assign n4116 = n4115 ^ x38 ^ 1'b0 ;
  assign n4117 = n4116 ^ n2863 ^ n2555 ;
  assign n4118 = ( n2555 & n2863 ) | ( n2555 & n4116 ) | ( n2863 & n4116 ) ;
  assign n4119 = x96 & n3344 ;
  assign n4120 = ( x98 & n3342 ) | ( x98 & n4119 ) | ( n3342 & n4119 ) ;
  assign n4121 = n4119 | n4120 ;
  assign n4122 = x97 & ~n3347 ;
  assign n4123 = ( x97 & n4121 ) | ( x97 & ~n4122 ) | ( n4121 & ~n4122 ) ;
  assign n4124 = n3346 & n4052 ;
  assign n4125 = n4123 | n4124 ;
  assign n4126 = n4125 ^ x29 ^ 1'b0 ;
  assign n4127 = n4126 ^ n3677 ^ n3327 ;
  assign n4128 = ( n3327 & n3677 ) | ( n3327 & n4126 ) | ( n3677 & n4126 ) ;
  assign n4129 = x96 & n2560 ;
  assign n4130 = ( x98 & n2567 ) | ( x98 & n4129 ) | ( n2567 & n4129 ) ;
  assign n4131 = n4129 | n4130 ;
  assign n4132 = x97 & ~n2562 ;
  assign n4133 = ( x97 & n4131 ) | ( x97 & ~n4132 ) | ( n4131 & ~n4132 ) ;
  assign n4134 = n2565 & n4052 ;
  assign n4135 = n4133 | n4134 ;
  assign n4136 = n4135 ^ x35 ^ 1'b0 ;
  assign n4137 = n4136 ^ n2875 ^ n2544 ;
  assign n4138 = ( n2544 & n2875 ) | ( n2544 & n4136 ) | ( n2875 & n4136 ) ;
  assign n4139 = x82 & n133 ;
  assign n4140 = x79 & n208 ;
  assign n4141 = ( x81 & n194 ) | ( x81 & n4140 ) | ( n194 & n4140 ) ;
  assign n4142 = n4140 | n4141 ;
  assign n4143 = x83 & ~n134 ;
  assign n4144 = ( x84 & n142 ) | ( x84 & n4139 ) | ( n142 & n4139 ) ;
  assign n4145 = n4139 | n4144 ;
  assign n4146 = ( x83 & ~n4143 ) | ( x83 & n4145 ) | ( ~n4143 & n4145 ) ;
  assign n4147 = x78 & ~n242 ;
  assign n4148 = x80 & ~n192 ;
  assign n4149 = ( x80 & n4142 ) | ( x80 & ~n4148 ) | ( n4142 & ~n4148 ) ;
  assign n4150 = x77 & n325 ;
  assign n4151 = ( x78 & ~n4147 ) | ( x78 & n4150 ) | ( ~n4147 & n4150 ) ;
  assign n4152 = ( n197 & n1258 ) | ( n197 & n4149 ) | ( n1258 & n4149 ) ;
  assign n4153 = n4149 | n4152 ;
  assign n4154 = n4153 ^ x62 ^ 1'b0 ;
  assign n4155 = n140 & n1355 ;
  assign n4156 = n4146 | n4155 ;
  assign n4157 = n4156 ^ x59 ^ 1'b0 ;
  assign n4158 = ( ~n2967 & n4151 ) | ( ~n2967 & n4154 ) | ( n4151 & n4154 ) ;
  assign n4159 = n4154 ^ n4151 ^ n2967 ;
  assign n4160 = n4159 ^ n4157 ^ n2974 ;
  assign n4161 = ( n2974 & n4157 ) | ( n2974 & ~n4159 ) | ( n4157 & ~n4159 ) ;
  assign n4162 = x85 & n263 ;
  assign n4163 = ( x87 & n264 ) | ( x87 & n4162 ) | ( n264 & n4162 ) ;
  assign n4164 = n4162 | n4163 ;
  assign n4165 = x86 & ~n260 ;
  assign n4166 = ( x86 & n4164 ) | ( x86 & ~n4165 ) | ( n4164 & ~n4165 ) ;
  assign n4167 = n272 & n1484 ;
  assign n4168 = n4166 | n4167 ;
  assign n4169 = n4168 ^ x56 ^ 1'b0 ;
  assign n4170 = ( n2978 & ~n4160 ) | ( n2978 & n4169 ) | ( ~n4160 & n4169 ) ;
  assign n4171 = n4169 ^ n4160 ^ n2978 ;
  assign n4172 = x88 & n408 ;
  assign n4173 = ( x90 & n403 ) | ( x90 & n4172 ) | ( n403 & n4172 ) ;
  assign n4174 = n4172 | n4173 ;
  assign n4175 = x89 & ~n410 ;
  assign n4176 = ( x89 & n4174 ) | ( x89 & ~n4175 ) | ( n4174 & ~n4175 ) ;
  assign n4177 = n402 & n1741 ;
  assign n4178 = n4176 | n4177 ;
  assign n4179 = n4178 ^ x53 ^ 1'b0 ;
  assign n4180 = ( n2988 & ~n4171 ) | ( n2988 & n4179 ) | ( ~n4171 & n4179 ) ;
  assign n4181 = n4179 ^ n4171 ^ n2988 ;
  assign n4182 = x91 & n561 ;
  assign n4183 = ( x93 & n551 ) | ( x93 & n4182 ) | ( n551 & n4182 ) ;
  assign n4184 = n4182 | n4183 ;
  assign n4185 = x92 & ~n550 ;
  assign n4186 = ( x92 & n4184 ) | ( x92 & ~n4185 ) | ( n4184 & ~n4185 ) ;
  assign n4187 = n553 & n2476 ;
  assign n4188 = n4186 | n4187 ;
  assign n4189 = n4188 ^ x50 ^ 1'b0 ;
  assign n4190 = ( n2998 & n4181 ) | ( n2998 & ~n4189 ) | ( n4181 & ~n4189 ) ;
  assign n4191 = n4189 ^ n4181 ^ n2998 ;
  assign n4192 = x94 & n744 ;
  assign n4193 = ( x96 & n730 ) | ( x96 & n4192 ) | ( n730 & n4192 ) ;
  assign n4194 = n4192 | n4193 ;
  assign n4195 = x95 & ~n732 ;
  assign n4196 = ( x95 & n4194 ) | ( x95 & ~n4195 ) | ( n4194 & ~n4195 ) ;
  assign n4197 = n731 & n2907 ;
  assign n4198 = n4196 | n4197 ;
  assign n4199 = n4198 ^ x47 ^ 1'b0 ;
  assign n4200 = n4199 ^ n4191 ^ n3007 ;
  assign n4201 = ( n3007 & n4191 ) | ( n3007 & n4199 ) | ( n4191 & n4199 ) ;
  assign n4202 = x80 & n208 ;
  assign n4203 = ( x82 & n194 ) | ( x82 & n4202 ) | ( n194 & n4202 ) ;
  assign n4204 = x78 & n325 ;
  assign n4205 = n4202 | n4203 ;
  assign n4206 = x79 & ~n242 ;
  assign n4207 = ( x79 & n4204 ) | ( x79 & ~n4206 ) | ( n4204 & ~n4206 ) ;
  assign n4208 = x81 & ~n192 ;
  assign n4209 = ( x81 & n4205 ) | ( x81 & ~n4208 ) | ( n4205 & ~n4208 ) ;
  assign n4210 = ( ~x14 & n2967 ) | ( ~x14 & n4207 ) | ( n2967 & n4207 ) ;
  assign n4211 = n4207 ^ n2967 ^ x14 ;
  assign n4212 = n197 & n1301 ;
  assign n4213 = n4209 | n4212 ;
  assign n4214 = n4213 ^ x62 ^ 1'b0 ;
  assign n4215 = n4214 ^ n4211 ^ n4158 ;
  assign n4216 = ( n4158 & ~n4211 ) | ( n4158 & n4214 ) | ( ~n4211 & n4214 ) ;
  assign n4217 = x83 & n133 ;
  assign n4218 = ( x85 & n142 ) | ( x85 & n4217 ) | ( n142 & n4217 ) ;
  assign n4219 = n4217 | n4218 ;
  assign n4220 = x84 & ~n134 ;
  assign n4221 = ( x84 & n4219 ) | ( x84 & ~n4220 ) | ( n4219 & ~n4220 ) ;
  assign n4222 = n140 & n1392 ;
  assign n4223 = n4221 | n4222 ;
  assign n4224 = n4223 ^ x59 ^ 1'b0 ;
  assign n4225 = n4224 ^ n4215 ^ n4161 ;
  assign n4226 = ( n4161 & ~n4215 ) | ( n4161 & n4224 ) | ( ~n4215 & n4224 ) ;
  assign n4227 = x86 & n263 ;
  assign n4228 = ( x88 & n264 ) | ( x88 & n4227 ) | ( n264 & n4227 ) ;
  assign n4229 = n4227 | n4228 ;
  assign n4230 = x87 & ~n260 ;
  assign n4231 = ( x87 & n4229 ) | ( x87 & ~n4230 ) | ( n4229 & ~n4230 ) ;
  assign n4232 = n272 & n1569 ;
  assign n4233 = n4231 | n4232 ;
  assign n4234 = n4233 ^ x56 ^ 1'b0 ;
  assign n4235 = n4234 ^ n4225 ^ n4170 ;
  assign n4236 = ( n4170 & ~n4225 ) | ( n4170 & n4234 ) | ( ~n4225 & n4234 ) ;
  assign n4237 = x89 & n408 ;
  assign n4238 = ( x91 & n403 ) | ( x91 & n4237 ) | ( n403 & n4237 ) ;
  assign n4239 = n4237 | n4238 ;
  assign n4240 = x90 & ~n410 ;
  assign n4241 = ( x90 & n4239 ) | ( x90 & ~n4240 ) | ( n4239 & ~n4240 ) ;
  assign n4242 = n402 & n2114 ;
  assign n4243 = n4241 | n4242 ;
  assign n4244 = n4243 ^ x53 ^ 1'b0 ;
  assign n4245 = n4244 ^ n4235 ^ n4180 ;
  assign n4246 = ( n4180 & ~n4235 ) | ( n4180 & n4244 ) | ( ~n4235 & n4244 ) ;
  assign n4247 = x92 & n561 ;
  assign n4248 = ( x94 & n551 ) | ( x94 & n4247 ) | ( n551 & n4247 ) ;
  assign n4249 = n4247 | n4248 ;
  assign n4250 = x93 & ~n550 ;
  assign n4251 = ( x93 & n4249 ) | ( x93 & ~n4250 ) | ( n4249 & ~n4250 ) ;
  assign n4252 = n553 & n2518 ;
  assign n4253 = n4251 | n4252 ;
  assign n4254 = n4253 ^ x50 ^ 1'b0 ;
  assign n4255 = ( n4190 & n4245 ) | ( n4190 & ~n4254 ) | ( n4245 & ~n4254 ) ;
  assign n4256 = n4254 ^ n4245 ^ n4190 ;
  assign n4257 = x95 & n744 ;
  assign n4258 = ( x97 & n730 ) | ( x97 & n4257 ) | ( n730 & n4257 ) ;
  assign n4259 = n4257 | n4258 ;
  assign n4260 = x96 & ~n732 ;
  assign n4261 = ( x96 & n4259 ) | ( x96 & ~n4260 ) | ( n4259 & ~n4260 ) ;
  assign n4262 = n731 & n3668 ;
  assign n4263 = n4261 | n4262 ;
  assign n4264 = n4263 ^ x47 ^ 1'b0 ;
  assign n4265 = n4264 ^ n4256 ^ n4201 ;
  assign n4266 = ( n4201 & n4256 ) | ( n4201 & n4264 ) | ( n4256 & n4264 ) ;
  assign n4267 = x97 & n3025 ;
  assign n4268 = ( x99 & n3015 ) | ( x99 & n4267 ) | ( n3015 & n4267 ) ;
  assign n4269 = n4267 | n4268 ;
  assign n4270 = n4080 ^ x99 ^ x98 ;
  assign n4271 = x98 & ~n3014 ;
  assign n4272 = ( x98 & n4269 ) | ( x98 & ~n4271 ) | ( n4269 & ~n4271 ) ;
  assign n4273 = n3017 & n4270 ;
  assign n4274 = n4272 | n4273 ;
  assign n4275 = n4274 ^ x32 ^ 1'b0 ;
  assign n4276 = n4275 ^ n4107 ^ n2927 ;
  assign n4277 = ( n2927 & n4107 ) | ( n2927 & n4275 ) | ( n4107 & n4275 ) ;
  assign n4278 = x97 & n2560 ;
  assign n4279 = ( x99 & n2567 ) | ( x99 & n4278 ) | ( n2567 & n4278 ) ;
  assign n4280 = n4278 | n4279 ;
  assign n4281 = x98 & ~n2562 ;
  assign n4282 = ( x98 & n4280 ) | ( x98 & ~n4281 ) | ( n4280 & ~n4281 ) ;
  assign n4283 = n2565 & n4270 ;
  assign n4284 = n4282 | n4283 ;
  assign n4285 = n4284 ^ x35 ^ 1'b0 ;
  assign n4286 = ( x98 & x99 ) | ( x98 & n4080 ) | ( x99 & n4080 ) ;
  assign n4287 = ( n2874 & n2937 ) | ( n2874 & n4285 ) | ( n2937 & n4285 ) ;
  assign n4288 = n4285 ^ n2937 ^ n2874 ;
  assign n4289 = x97 & n3734 ;
  assign n4290 = ( x99 & n3732 ) | ( x99 & n4289 ) | ( n3732 & n4289 ) ;
  assign n4291 = n4289 | n4290 ;
  assign n4292 = x98 & ~n3737 ;
  assign n4293 = ( x98 & n4291 ) | ( x98 & ~n4292 ) | ( n4291 & ~n4292 ) ;
  assign n4294 = n3736 & n4270 ;
  assign n4295 = n4293 | n4294 ;
  assign n4296 = n4295 ^ x26 ^ 1'b0 ;
  assign n4297 = n4296 ^ n4088 ^ n3666 ;
  assign n4298 = ( n3666 & n4088 ) | ( n3666 & n4296 ) | ( n4088 & n4296 ) ;
  assign n4299 = x97 & n3344 ;
  assign n4300 = ( x99 & n3342 ) | ( x99 & n4299 ) | ( n3342 & n4299 ) ;
  assign n4301 = n4299 | n4300 ;
  assign n4302 = x98 & ~n3347 ;
  assign n4303 = ( x98 & n4301 ) | ( x98 & ~n4302 ) | ( n4301 & ~n4302 ) ;
  assign n4304 = n3346 & n4270 ;
  assign n4305 = n4303 | n4304 ;
  assign n4306 = n4305 ^ x29 ^ 1'b0 ;
  assign n4307 = ( n3338 & n4128 ) | ( n3338 & n4306 ) | ( n4128 & n4306 ) ;
  assign n4308 = n4306 ^ n4128 ^ n3338 ;
  assign n4309 = x97 & n2156 ;
  assign n4310 = ( x99 & n2163 ) | ( x99 & n4309 ) | ( n2163 & n4309 ) ;
  assign n4311 = n4309 | n4310 ;
  assign n4312 = x98 & ~n2158 ;
  assign n4313 = ( x98 & n4311 ) | ( x98 & ~n4312 ) | ( n4311 & ~n4312 ) ;
  assign n4314 = n2161 & n4270 ;
  assign n4315 = n4313 | n4314 ;
  assign n4316 = n4315 ^ x38 ^ 1'b0 ;
  assign n4317 = ( n2864 & n2917 ) | ( n2864 & n4316 ) | ( n2917 & n4316 ) ;
  assign n4318 = n4316 ^ n2917 ^ n2864 ;
  assign n4319 = x97 & n888 ;
  assign n4320 = ( x99 & n878 ) | ( x99 & n4319 ) | ( n878 & n4319 ) ;
  assign n4321 = n4319 | n4320 ;
  assign n4322 = x98 & ~n877 ;
  assign n4323 = ( x98 & n4321 ) | ( x98 & ~n4322 ) | ( n4321 & ~n4322 ) ;
  assign n4324 = n880 & n4270 ;
  assign n4325 = n4323 | n4324 ;
  assign n4326 = n4325 ^ x44 ^ 1'b0 ;
  assign n4327 = ( n3009 & n4200 ) | ( n3009 & n4326 ) | ( n4200 & n4326 ) ;
  assign n4328 = n4326 ^ n4200 ^ n3009 ;
  assign n4329 = x98 & n2156 ;
  assign n4330 = ( x100 & n2163 ) | ( x100 & n4329 ) | ( n2163 & n4329 ) ;
  assign n4331 = x99 & ~n2158 ;
  assign n4332 = n4329 | n4330 ;
  assign n4333 = ( x99 & ~n4331 ) | ( x99 & n4332 ) | ( ~n4331 & n4332 ) ;
  assign n4334 = n4286 ^ x100 ^ x99 ;
  assign n4335 = n2161 & n4334 ;
  assign n4336 = n4333 | n4335 ;
  assign n4337 = n4336 ^ x38 ^ 1'b0 ;
  assign n4338 = n4337 ^ n4317 ^ n3707 ;
  assign n4339 = ( n3707 & n4317 ) | ( n3707 & n4337 ) | ( n4317 & n4337 ) ;
  assign n4340 = x98 & n3734 ;
  assign n4341 = ( x100 & n3732 ) | ( x100 & n4340 ) | ( n3732 & n4340 ) ;
  assign n4342 = n4340 | n4341 ;
  assign n4343 = x99 & ~n3737 ;
  assign n4344 = ( x99 & n4342 ) | ( x99 & ~n4343 ) | ( n4342 & ~n4343 ) ;
  assign n4345 = n3736 & n4334 ;
  assign n4346 = n4344 | n4345 ;
  assign n4347 = n4346 ^ x26 ^ 1'b0 ;
  assign n4348 = n4347 ^ n4298 ^ n3678 ;
  assign n4349 = ( n3678 & n4298 ) | ( n3678 & n4347 ) | ( n4298 & n4347 ) ;
  assign n4350 = x98 & n3344 ;
  assign n4351 = ( x100 & n3342 ) | ( x100 & n4350 ) | ( n3342 & n4350 ) ;
  assign n4352 = n4350 | n4351 ;
  assign n4353 = x99 & ~n3347 ;
  assign n4354 = ( x99 & n4352 ) | ( x99 & ~n4353 ) | ( n4352 & ~n4353 ) ;
  assign n4355 = n3346 & n4334 ;
  assign n4356 = n4354 | n4355 ;
  assign n4357 = n4356 ^ x29 ^ 1'b0 ;
  assign n4358 = n4357 ^ n4307 ^ n3717 ;
  assign n4359 = ( n3717 & n4307 ) | ( n3717 & n4357 ) | ( n4307 & n4357 ) ;
  assign n4360 = x98 & n888 ;
  assign n4361 = ( x100 & n878 ) | ( x100 & n4360 ) | ( n878 & n4360 ) ;
  assign n4362 = n4360 | n4361 ;
  assign n4363 = x99 & ~n877 ;
  assign n4364 = ( x99 & n4362 ) | ( x99 & ~n4363 ) | ( n4362 & ~n4363 ) ;
  assign n4365 = n880 & n4334 ;
  assign n4366 = n4364 | n4365 ;
  assign n4367 = n4366 ^ x44 ^ 1'b0 ;
  assign n4368 = n4367 ^ n4327 ^ n4265 ;
  assign n4369 = ( n4265 & n4327 ) | ( n4265 & n4367 ) | ( n4327 & n4367 ) ;
  assign n4370 = x98 & n2560 ;
  assign n4371 = ( x100 & n2567 ) | ( x100 & n4370 ) | ( n2567 & n4370 ) ;
  assign n4372 = n4370 | n4371 ;
  assign n4373 = x99 & ~n2562 ;
  assign n4374 = ( x99 & n4372 ) | ( x99 & ~n4373 ) | ( n4372 & ~n4373 ) ;
  assign n4375 = n2565 & n4334 ;
  assign n4376 = n4374 | n4375 ;
  assign n4377 = n4376 ^ x35 ^ 1'b0 ;
  assign n4378 = n4377 ^ n4287 ^ n3727 ;
  assign n4379 = ( n3727 & n4287 ) | ( n3727 & n4377 ) | ( n4287 & n4377 ) ;
  assign n4380 = x98 & n3025 ;
  assign n4381 = ( x100 & n3015 ) | ( x100 & n4380 ) | ( n3015 & n4380 ) ;
  assign n4382 = n4380 | n4381 ;
  assign n4383 = x99 & ~n3014 ;
  assign n4384 = ( x99 & n4382 ) | ( x99 & ~n4383 ) | ( n4382 & ~n4383 ) ;
  assign n4385 = ( n3017 & n4334 ) | ( n3017 & n4384 ) | ( n4334 & n4384 ) ;
  assign n4386 = n4384 | n4385 ;
  assign n4387 = n4386 ^ x32 ^ 1'b0 ;
  assign n4388 = ( n2926 & n3698 ) | ( n2926 & n4387 ) | ( n3698 & n4387 ) ;
  assign n4389 = n4387 ^ n3698 ^ n2926 ;
  assign n4390 = x80 & ~n242 ;
  assign n4391 = x84 & n133 ;
  assign n4392 = ( x86 & n142 ) | ( x86 & n4391 ) | ( n142 & n4391 ) ;
  assign n4393 = n4391 | n4392 ;
  assign n4394 = x81 & n208 ;
  assign n4395 = x79 & n325 ;
  assign n4396 = ( x80 & ~n4390 ) | ( x80 & n4395 ) | ( ~n4390 & n4395 ) ;
  assign n4397 = ( x83 & n194 ) | ( x83 & n4394 ) | ( n194 & n4394 ) ;
  assign n4398 = n4394 | n4397 ;
  assign n4399 = x82 & ~n192 ;
  assign n4400 = ( x82 & n4398 ) | ( x82 & ~n4399 ) | ( n4398 & ~n4399 ) ;
  assign n4401 = ( n197 & n1329 ) | ( n197 & n4400 ) | ( n1329 & n4400 ) ;
  assign n4402 = n4400 | n4401 ;
  assign n4403 = x85 & ~n134 ;
  assign n4404 = n4402 ^ x62 ^ 1'b0 ;
  assign n4405 = ( x85 & n4393 ) | ( x85 & ~n4403 ) | ( n4393 & ~n4403 ) ;
  assign n4406 = n140 & n1419 ;
  assign n4407 = n4405 | n4406 ;
  assign n4408 = n4404 ^ n4396 ^ n4210 ;
  assign n4409 = ( n4210 & ~n4396 ) | ( n4210 & n4404 ) | ( ~n4396 & n4404 ) ;
  assign n4410 = n4407 ^ x59 ^ 1'b0 ;
  assign n4411 = n4410 ^ n4408 ^ n4216 ;
  assign n4412 = ( n4216 & ~n4408 ) | ( n4216 & n4410 ) | ( ~n4408 & n4410 ) ;
  assign n4413 = x87 & n263 ;
  assign n4414 = ( x89 & n264 ) | ( x89 & n4413 ) | ( n264 & n4413 ) ;
  assign n4415 = n4413 | n4414 ;
  assign n4416 = x88 & ~n260 ;
  assign n4417 = ( x88 & n4415 ) | ( x88 & ~n4416 ) | ( n4415 & ~n4416 ) ;
  assign n4418 = n272 & n1654 ;
  assign n4419 = n4417 | n4418 ;
  assign n4420 = n4419 ^ x56 ^ 1'b0 ;
  assign n4421 = ( n4226 & ~n4411 ) | ( n4226 & n4420 ) | ( ~n4411 & n4420 ) ;
  assign n4422 = n4420 ^ n4411 ^ n4226 ;
  assign n4423 = x90 & n408 ;
  assign n4424 = ( x92 & n403 ) | ( x92 & n4423 ) | ( n403 & n4423 ) ;
  assign n4425 = n4423 | n4424 ;
  assign n4426 = x91 & ~n410 ;
  assign n4427 = ( x91 & n4425 ) | ( x91 & ~n4426 ) | ( n4425 & ~n4426 ) ;
  assign n4428 = n402 & n2420 ;
  assign n4429 = n4427 | n4428 ;
  assign n4430 = n4429 ^ x53 ^ 1'b0 ;
  assign n4431 = n4430 ^ n4422 ^ n4236 ;
  assign n4432 = ( n4236 & ~n4422 ) | ( n4236 & n4430 ) | ( ~n4422 & n4430 ) ;
  assign n4433 = x93 & n561 ;
  assign n4434 = ( x95 & n551 ) | ( x95 & n4433 ) | ( n551 & n4433 ) ;
  assign n4435 = n4433 | n4434 ;
  assign n4436 = x94 & ~n550 ;
  assign n4437 = ( x94 & n4435 ) | ( x94 & ~n4436 ) | ( n4435 & ~n4436 ) ;
  assign n4438 = n553 & n2854 ;
  assign n4439 = n4437 | n4438 ;
  assign n4440 = n4439 ^ x50 ^ 1'b0 ;
  assign n4441 = ( n4246 & ~n4431 ) | ( n4246 & n4440 ) | ( ~n4431 & n4440 ) ;
  assign n4442 = n4440 ^ n4431 ^ n4246 ;
  assign n4443 = ( x99 & x100 ) | ( x99 & n4286 ) | ( x100 & n4286 ) ;
  assign n4444 = x96 & n744 ;
  assign n4445 = ( x98 & n730 ) | ( x98 & n4444 ) | ( n730 & n4444 ) ;
  assign n4446 = n4444 | n4445 ;
  assign n4447 = x97 & ~n732 ;
  assign n4448 = ( x97 & n4446 ) | ( x97 & ~n4447 ) | ( n4446 & ~n4447 ) ;
  assign n4449 = n731 & n4052 ;
  assign n4450 = n4448 | n4449 ;
  assign n4451 = n4450 ^ x47 ^ 1'b0 ;
  assign n4452 = ( n4255 & n4442 ) | ( n4255 & ~n4451 ) | ( n4442 & ~n4451 ) ;
  assign n4453 = n4451 ^ n4442 ^ n4255 ;
  assign n4454 = x92 & ~n410 ;
  assign n4455 = x91 & n408 ;
  assign n4456 = ( x93 & n403 ) | ( x93 & n4455 ) | ( n403 & n4455 ) ;
  assign n4457 = n4455 | n4456 ;
  assign n4458 = ( x92 & ~n4454 ) | ( x92 & n4457 ) | ( ~n4454 & n4457 ) ;
  assign n4459 = x97 & n1058 ;
  assign n4460 = ( x99 & n1065 ) | ( x99 & n4459 ) | ( n1065 & n4459 ) ;
  assign n4461 = n4459 | n4460 ;
  assign n4462 = x98 & ~n1060 ;
  assign n4463 = ( x98 & n4461 ) | ( x98 & ~n4462 ) | ( n4461 & ~n4462 ) ;
  assign n4464 = n1063 & n4270 ;
  assign n4465 = n4463 | n4464 ;
  assign n4466 = n4465 ^ x41 ^ 1'b0 ;
  assign n4467 = n402 & n2476 ;
  assign n4468 = n4458 | n4467 ;
  assign n4469 = n4468 ^ x53 ^ 1'b0 ;
  assign n4470 = ( n2895 & n2947 ) | ( n2895 & n4466 ) | ( n2947 & n4466 ) ;
  assign n4471 = n4466 ^ n2947 ^ n2895 ;
  assign n4472 = x98 & n1058 ;
  assign n4473 = ( x100 & n1065 ) | ( x100 & n4472 ) | ( n1065 & n4472 ) ;
  assign n4474 = n4472 | n4473 ;
  assign n4475 = x99 & ~n1060 ;
  assign n4476 = ( x99 & n4474 ) | ( x99 & ~n4475 ) | ( n4474 & ~n4475 ) ;
  assign n4477 = n1063 & n4334 ;
  assign n4478 = n4476 | n4477 ;
  assign n4479 = n4478 ^ x41 ^ 1'b0 ;
  assign n4480 = n4479 ^ n4470 ^ n3688 ;
  assign n4481 = ( n3688 & n4470 ) | ( n3688 & n4479 ) | ( n4470 & n4479 ) ;
  assign n4482 = x94 & n561 ;
  assign n4483 = ( x96 & n551 ) | ( x96 & n4482 ) | ( n551 & n4482 ) ;
  assign n4484 = n4482 | n4483 ;
  assign n4485 = x95 & ~n550 ;
  assign n4486 = ( x95 & n4484 ) | ( x95 & ~n4485 ) | ( n4484 & ~n4485 ) ;
  assign n4487 = n553 & n2907 ;
  assign n4488 = n4486 | n4487 ;
  assign n4489 = n4488 ^ x50 ^ 1'b0 ;
  assign n4490 = x81 & ~n242 ;
  assign n4491 = x82 & n208 ;
  assign n4492 = x83 & ~n192 ;
  assign n4493 = ( x84 & n194 ) | ( x84 & n4491 ) | ( n194 & n4491 ) ;
  assign n4494 = n4491 | n4493 ;
  assign n4495 = x85 & n133 ;
  assign n4496 = ( x83 & ~n4492 ) | ( x83 & n4494 ) | ( ~n4492 & n4494 ) ;
  assign n4497 = ( x87 & n142 ) | ( x87 & n4495 ) | ( n142 & n4495 ) ;
  assign n4498 = n4495 | n4497 ;
  assign n4499 = x86 & ~n134 ;
  assign n4500 = ( x86 & n4498 ) | ( x86 & ~n4499 ) | ( n4498 & ~n4499 ) ;
  assign n4501 = x80 & n325 ;
  assign n4502 = ( x81 & ~n4490 ) | ( x81 & n4501 ) | ( ~n4490 & n4501 ) ;
  assign n4503 = n197 & n1355 ;
  assign n4504 = n4496 | n4503 ;
  assign n4505 = n140 & n1484 ;
  assign n4506 = n4504 ^ x62 ^ 1'b0 ;
  assign n4507 = n4500 | n4505 ;
  assign n4508 = n4506 ^ n4502 ^ n4396 ;
  assign n4509 = ( n4396 & ~n4502 ) | ( n4396 & n4506 ) | ( ~n4502 & n4506 ) ;
  assign n4510 = n4507 ^ x59 ^ 1'b0 ;
  assign n4511 = ( n4409 & ~n4508 ) | ( n4409 & n4510 ) | ( ~n4508 & n4510 ) ;
  assign n4512 = n4510 ^ n4508 ^ n4409 ;
  assign n4513 = x88 & n263 ;
  assign n4514 = ( x90 & n264 ) | ( x90 & n4513 ) | ( n264 & n4513 ) ;
  assign n4515 = n4513 | n4514 ;
  assign n4516 = x89 & ~n260 ;
  assign n4517 = ( x89 & n4515 ) | ( x89 & ~n4516 ) | ( n4515 & ~n4516 ) ;
  assign n4518 = n272 & n1741 ;
  assign n4519 = n4517 | n4518 ;
  assign n4520 = n4519 ^ x56 ^ 1'b0 ;
  assign n4521 = ( n4412 & ~n4512 ) | ( n4412 & n4520 ) | ( ~n4512 & n4520 ) ;
  assign n4522 = n4520 ^ n4512 ^ n4412 ;
  assign n4523 = n4522 ^ n4469 ^ n4421 ;
  assign n4524 = ( n4432 & n4489 ) | ( n4432 & ~n4523 ) | ( n4489 & ~n4523 ) ;
  assign n4525 = n4523 ^ n4489 ^ n4432 ;
  assign n4526 = x97 & n744 ;
  assign n4527 = ( x99 & n730 ) | ( x99 & n4526 ) | ( n730 & n4526 ) ;
  assign n4528 = n4526 | n4527 ;
  assign n4529 = x95 & n561 ;
  assign n4530 = ( n4421 & n4469 ) | ( n4421 & ~n4522 ) | ( n4469 & ~n4522 ) ;
  assign n4531 = x98 & ~n732 ;
  assign n4532 = ( x98 & n4528 ) | ( x98 & ~n4531 ) | ( n4528 & ~n4531 ) ;
  assign n4533 = ( x97 & n551 ) | ( x97 & n4529 ) | ( n551 & n4529 ) ;
  assign n4534 = n731 & n4270 ;
  assign n4535 = n4532 | n4534 ;
  assign n4536 = n4529 | n4533 ;
  assign n4537 = n4535 ^ x47 ^ 1'b0 ;
  assign n4538 = ( n4441 & ~n4525 ) | ( n4441 & n4537 ) | ( ~n4525 & n4537 ) ;
  assign n4539 = n4537 ^ n4525 ^ n4441 ;
  assign n4540 = x81 & n325 ;
  assign n4541 = x82 & ~n242 ;
  assign n4542 = ( x82 & n4540 ) | ( x82 & ~n4541 ) | ( n4540 & ~n4541 ) ;
  assign n4543 = x83 & n208 ;
  assign n4544 = ( x85 & n194 ) | ( x85 & n4543 ) | ( n194 & n4543 ) ;
  assign n4545 = n4543 | n4544 ;
  assign n4546 = x84 & ~n192 ;
  assign n4547 = ( x84 & n4545 ) | ( x84 & ~n4546 ) | ( n4545 & ~n4546 ) ;
  assign n4548 = n197 & n1392 ;
  assign n4549 = n4547 | n4548 ;
  assign n4550 = n4549 ^ x62 ^ 1'b0 ;
  assign n4551 = ( ~x17 & n4502 ) | ( ~x17 & n4542 ) | ( n4502 & n4542 ) ;
  assign n4552 = n4542 ^ n4502 ^ x17 ;
  assign n4553 = ( n4509 & n4550 ) | ( n4509 & ~n4552 ) | ( n4550 & ~n4552 ) ;
  assign n4554 = n4552 ^ n4550 ^ n4509 ;
  assign n4555 = x86 & n133 ;
  assign n4556 = ( x88 & n142 ) | ( x88 & n4555 ) | ( n142 & n4555 ) ;
  assign n4557 = n4555 | n4556 ;
  assign n4558 = x87 & ~n134 ;
  assign n4559 = ( x87 & n4557 ) | ( x87 & ~n4558 ) | ( n4557 & ~n4558 ) ;
  assign n4560 = n140 & n1569 ;
  assign n4561 = n4559 | n4560 ;
  assign n4562 = n4561 ^ x59 ^ 1'b0 ;
  assign n4563 = ( n4511 & ~n4554 ) | ( n4511 & n4562 ) | ( ~n4554 & n4562 ) ;
  assign n4564 = n4562 ^ n4554 ^ n4511 ;
  assign n4565 = x89 & n263 ;
  assign n4566 = ( x91 & n264 ) | ( x91 & n4565 ) | ( n264 & n4565 ) ;
  assign n4567 = n4565 | n4566 ;
  assign n4568 = x90 & ~n260 ;
  assign n4569 = ( x90 & n4567 ) | ( x90 & ~n4568 ) | ( n4567 & ~n4568 ) ;
  assign n4570 = n272 & n2114 ;
  assign n4571 = n4569 | n4570 ;
  assign n4572 = n4571 ^ x56 ^ 1'b0 ;
  assign n4573 = n4572 ^ n4564 ^ n4521 ;
  assign n4574 = ( n4521 & ~n4564 ) | ( n4521 & n4572 ) | ( ~n4564 & n4572 ) ;
  assign n4575 = x92 & n408 ;
  assign n4576 = x96 & ~n550 ;
  assign n4577 = ( x96 & n4536 ) | ( x96 & ~n4576 ) | ( n4536 & ~n4576 ) ;
  assign n4578 = ( x94 & n403 ) | ( x94 & n4575 ) | ( n403 & n4575 ) ;
  assign n4579 = n4575 | n4578 ;
  assign n4580 = x93 & ~n410 ;
  assign n4581 = ( x93 & n4579 ) | ( x93 & ~n4580 ) | ( n4579 & ~n4580 ) ;
  assign n4582 = n402 & n2518 ;
  assign n4583 = n4581 | n4582 ;
  assign n4584 = n4583 ^ x53 ^ 1'b0 ;
  assign n4585 = n553 & n3668 ;
  assign n4586 = n4577 | n4585 ;
  assign n4587 = n4584 ^ n4573 ^ n4530 ;
  assign n4588 = ( n4530 & ~n4573 ) | ( n4530 & n4584 ) | ( ~n4573 & n4584 ) ;
  assign n4589 = x98 & n744 ;
  assign n4590 = ( x100 & n730 ) | ( x100 & n4589 ) | ( n730 & n4589 ) ;
  assign n4591 = n4589 | n4590 ;
  assign n4592 = x99 & ~n732 ;
  assign n4593 = ( x99 & n4591 ) | ( x99 & ~n4592 ) | ( n4591 & ~n4592 ) ;
  assign n4594 = n731 & n4334 ;
  assign n4595 = n4593 | n4594 ;
  assign n4596 = n4595 ^ x47 ^ 1'b0 ;
  assign n4597 = n4586 ^ x50 ^ 1'b0 ;
  assign n4598 = n4597 ^ n4587 ^ n4524 ;
  assign n4599 = ( n4524 & ~n4587 ) | ( n4524 & n4597 ) | ( ~n4587 & n4597 ) ;
  assign n4600 = n4598 ^ n4596 ^ n4538 ;
  assign n4601 = ( n4538 & n4596 ) | ( n4538 & ~n4598 ) | ( n4596 & ~n4598 ) ;
  assign n4602 = x22 ^ x21 ^ 1'b0 ;
  assign n4603 = x21 ^ x20 ^ 1'b0 ;
  assign n4604 = x23 ^ x22 ^ 1'b0 ;
  assign n4605 = n4602 & ~n4603 ;
  assign n4606 = n4603 & ~n4604 ;
  assign n4607 = ~x65 & n4606 ;
  assign n4608 = n4603 & n4604 ;
  assign n4609 = x64 & n4605 ;
  assign n4610 = ( n4606 & ~n4607 ) | ( n4606 & n4609 ) | ( ~n4607 & n4609 ) ;
  assign n4611 = ( n190 & n4608 ) | ( n190 & n4609 ) | ( n4608 & n4609 ) ;
  assign n4612 = n139 & n4608 ;
  assign n4613 = n4610 | n4611 ;
  assign n4614 = x65 & ~n4605 ;
  assign n4615 = ( n4602 & ~n4603 ) | ( n4602 & n4604 ) | ( ~n4603 & n4604 ) ;
  assign n4616 = ~n4602 & n4615 ;
  assign n4617 = x64 & n4616 ;
  assign n4618 = ( x66 & n4606 ) | ( x66 & n4617 ) | ( n4606 & n4617 ) ;
  assign n4619 = n4617 | n4618 ;
  assign n4620 = x64 & n4603 ;
  assign n4621 = ( x65 & ~n4614 ) | ( x65 & n4619 ) | ( ~n4614 & n4619 ) ;
  assign n4622 = x23 & ~n4620 ;
  assign n4623 = n4612 | n4621 ;
  assign n4624 = n4623 ^ x23 ^ 1'b0 ;
  assign n4625 = n4613 ^ x23 ^ 1'b0 ;
  assign n4626 = n4622 & n4625 ;
  assign n4627 = n4626 ^ n4624 ^ 1'b0 ;
  assign n4628 = n4624 & n4626 ;
  assign n4629 = n4625 ^ n4622 ^ 1'b0 ;
  assign n4630 = x65 & n4616 ;
  assign n4631 = ( x67 & n4606 ) | ( x67 & n4630 ) | ( n4606 & n4630 ) ;
  assign n4632 = n4630 | n4631 ;
  assign n4633 = x66 & ~n4605 ;
  assign n4634 = ( x66 & n4632 ) | ( x66 & ~n4633 ) | ( n4632 & ~n4633 ) ;
  assign n4635 = n161 & n4608 ;
  assign n4636 = n4634 | n4635 ;
  assign n4637 = n4636 ^ x23 ^ 1'b0 ;
  assign n4638 = ( n3740 & n4628 ) | ( n3740 & n4637 ) | ( n4628 & n4637 ) ;
  assign n4639 = n4637 ^ n4628 ^ n3740 ;
  assign n4640 = x66 & n4616 ;
  assign n4641 = ( x68 & n4606 ) | ( x68 & n4640 ) | ( n4606 & n4640 ) ;
  assign n4642 = n4640 | n4641 ;
  assign n4643 = x67 & ~n4605 ;
  assign n4644 = ( x67 & n4642 ) | ( x67 & ~n4643 ) | ( n4642 & ~n4643 ) ;
  assign n4645 = n175 & n4608 ;
  assign n4646 = n4644 | n4645 ;
  assign n4647 = n4646 ^ x23 ^ 1'b0 ;
  assign n4648 = n4647 ^ n4638 ^ n3755 ;
  assign n4649 = ( n3755 & n4638 ) | ( n3755 & n4647 ) | ( n4638 & n4647 ) ;
  assign n4650 = x67 & n4616 ;
  assign n4651 = ( x69 & n4606 ) | ( x69 & n4650 ) | ( n4606 & n4650 ) ;
  assign n4652 = n4650 | n4651 ;
  assign n4653 = x68 & ~n4605 ;
  assign n4654 = ( x68 & n4652 ) | ( x68 & ~n4653 ) | ( n4652 & ~n4653 ) ;
  assign n4655 = n172 & n4608 ;
  assign n4656 = n4654 | n4655 ;
  assign n4657 = n4656 ^ x23 ^ 1'b0 ;
  assign n4658 = n4657 ^ n4649 ^ n3764 ;
  assign n4659 = ( n3764 & n4649 ) | ( n3764 & n4657 ) | ( n4649 & n4657 ) ;
  assign n4660 = x68 & n4616 ;
  assign n4661 = ( x70 & n4606 ) | ( x70 & n4660 ) | ( n4606 & n4660 ) ;
  assign n4662 = n4660 | n4661 ;
  assign n4663 = x69 & ~n4605 ;
  assign n4664 = ( x69 & n4662 ) | ( x69 & ~n4663 ) | ( n4662 & ~n4663 ) ;
  assign n4665 = n168 & n4608 ;
  assign n4666 = n4664 | n4665 ;
  assign n4667 = n4666 ^ x23 ^ 1'b0 ;
  assign n4668 = n4667 ^ n4659 ^ n3765 ;
  assign n4669 = ( n3765 & n4659 ) | ( n3765 & n4667 ) | ( n4659 & n4667 ) ;
  assign n4670 = x69 & n4616 ;
  assign n4671 = ( x71 & n4606 ) | ( x71 & n4670 ) | ( n4606 & n4670 ) ;
  assign n4672 = n4670 | n4671 ;
  assign n4673 = x70 & ~n4605 ;
  assign n4674 = ( x70 & n4672 ) | ( x70 & ~n4673 ) | ( n4672 & ~n4673 ) ;
  assign n4675 = n328 & n4608 ;
  assign n4676 = n4674 | n4675 ;
  assign n4677 = n4676 ^ x23 ^ 1'b0 ;
  assign n4678 = n4677 ^ n4669 ^ n3775 ;
  assign n4679 = ( n3775 & n4669 ) | ( n3775 & n4677 ) | ( n4669 & n4677 ) ;
  assign n4680 = x70 & n4616 ;
  assign n4681 = ( x72 & n4606 ) | ( x72 & n4680 ) | ( n4606 & n4680 ) ;
  assign n4682 = n4680 | n4681 ;
  assign n4683 = x71 & ~n4605 ;
  assign n4684 = ( x71 & n4682 ) | ( x71 & ~n4683 ) | ( n4682 & ~n4683 ) ;
  assign n4685 = n349 & n4608 ;
  assign n4686 = n4684 | n4685 ;
  assign n4687 = n4686 ^ x23 ^ 1'b0 ;
  assign n4688 = ( n3786 & n4679 ) | ( n3786 & n4687 ) | ( n4679 & n4687 ) ;
  assign n4689 = n4687 ^ n4679 ^ n3786 ;
  assign n4690 = x71 & n4616 ;
  assign n4691 = ( x73 & n4606 ) | ( x73 & n4690 ) | ( n4606 & n4690 ) ;
  assign n4692 = n4690 | n4691 ;
  assign n4693 = x72 & ~n4605 ;
  assign n4694 = ( x72 & n4692 ) | ( x72 & ~n4693 ) | ( n4692 & ~n4693 ) ;
  assign n4695 = n370 & n4608 ;
  assign n4696 = n4694 | n4695 ;
  assign n4697 = n4696 ^ x23 ^ 1'b0 ;
  assign n4698 = ( n3796 & n4688 ) | ( n3796 & n4697 ) | ( n4688 & n4697 ) ;
  assign n4699 = n4697 ^ n4688 ^ n3796 ;
  assign n4700 = x72 & n4616 ;
  assign n4701 = ( x74 & n4606 ) | ( x74 & n4700 ) | ( n4606 & n4700 ) ;
  assign n4702 = n4700 | n4701 ;
  assign n4703 = x73 & ~n4605 ;
  assign n4704 = ( x73 & n4702 ) | ( x73 & ~n4703 ) | ( n4702 & ~n4703 ) ;
  assign n4705 = n504 & n4608 ;
  assign n4706 = n4704 | n4705 ;
  assign n4707 = n4706 ^ x23 ^ 1'b0 ;
  assign n4708 = n4707 ^ n4698 ^ n3806 ;
  assign n4709 = ( n3806 & n4698 ) | ( n3806 & n4707 ) | ( n4698 & n4707 ) ;
  assign n4710 = x73 & n4616 ;
  assign n4711 = ( x75 & n4606 ) | ( x75 & n4710 ) | ( n4606 & n4710 ) ;
  assign n4712 = n4710 | n4711 ;
  assign n4713 = x74 & ~n4605 ;
  assign n4714 = ( x74 & n4712 ) | ( x74 & ~n4713 ) | ( n4712 & ~n4713 ) ;
  assign n4715 = n525 & n4608 ;
  assign n4716 = n4714 | n4715 ;
  assign n4717 = n4716 ^ x23 ^ 1'b0 ;
  assign n4718 = n4717 ^ n4709 ^ n3815 ;
  assign n4719 = ( n3815 & n4709 ) | ( n3815 & n4717 ) | ( n4709 & n4717 ) ;
  assign n4720 = x74 & n4616 ;
  assign n4721 = ( x76 & n4606 ) | ( x76 & n4720 ) | ( n4606 & n4720 ) ;
  assign n4722 = n4720 | n4721 ;
  assign n4723 = x75 & ~n4605 ;
  assign n4724 = ( x75 & n4722 ) | ( x75 & ~n4723 ) | ( n4722 & ~n4723 ) ;
  assign n4725 = n664 & n4608 ;
  assign n4726 = n4724 | n4725 ;
  assign n4727 = n4726 ^ x23 ^ 1'b0 ;
  assign n4728 = ( n3825 & n4719 ) | ( n3825 & n4727 ) | ( n4719 & n4727 ) ;
  assign n4729 = n4727 ^ n4719 ^ n3825 ;
  assign n4730 = x75 & n4616 ;
  assign n4731 = ( x77 & n4606 ) | ( x77 & n4730 ) | ( n4606 & n4730 ) ;
  assign n4732 = n4730 | n4731 ;
  assign n4733 = x76 & ~n4605 ;
  assign n4734 = ( x76 & n4732 ) | ( x76 & ~n4733 ) | ( n4732 & ~n4733 ) ;
  assign n4735 = n690 & n4608 ;
  assign n4736 = n4734 | n4735 ;
  assign n4737 = n4736 ^ x23 ^ 1'b0 ;
  assign n4738 = n4737 ^ n4728 ^ n3835 ;
  assign n4739 = ( n3835 & n4728 ) | ( n3835 & n4737 ) | ( n4728 & n4737 ) ;
  assign n4740 = x79 & n4616 ;
  assign n4741 = ( x81 & n4606 ) | ( x81 & n4740 ) | ( n4606 & n4740 ) ;
  assign n4742 = n4740 | n4741 ;
  assign n4743 = n1015 & n4608 ;
  assign n4744 = x77 & n4616 ;
  assign n4745 = ( x79 & n4606 ) | ( x79 & n4744 ) | ( n4606 & n4744 ) ;
  assign n4746 = n4744 | n4745 ;
  assign n4747 = x78 & ~n4605 ;
  assign n4748 = ( x78 & n4746 ) | ( x78 & ~n4747 ) | ( n4746 & ~n4747 ) ;
  assign n4749 = x76 & n4616 ;
  assign n4750 = n4743 | n4748 ;
  assign n4751 = ( x78 & n4606 ) | ( x78 & n4749 ) | ( n4606 & n4749 ) ;
  assign n4752 = n4749 | n4751 ;
  assign n4753 = x77 & ~n4605 ;
  assign n4754 = ( x77 & n4752 ) | ( x77 & ~n4753 ) | ( n4752 & ~n4753 ) ;
  assign n4755 = n709 & n4608 ;
  assign n4756 = n4754 | n4755 ;
  assign n4757 = x80 & ~n4605 ;
  assign n4758 = ( x80 & n4742 ) | ( x80 & ~n4757 ) | ( n4742 & ~n4757 ) ;
  assign n4759 = n1258 & n4608 ;
  assign n4760 = n4756 ^ x23 ^ 1'b0 ;
  assign n4761 = n4758 | n4759 ;
  assign n4762 = ( n3846 & n4739 ) | ( n3846 & n4760 ) | ( n4739 & n4760 ) ;
  assign n4763 = n4760 ^ n4739 ^ n3846 ;
  assign n4764 = x78 & n4616 ;
  assign n4765 = ( x80 & n4606 ) | ( x80 & n4764 ) | ( n4606 & n4764 ) ;
  assign n4766 = n4764 | n4765 ;
  assign n4767 = n4761 ^ x23 ^ 1'b0 ;
  assign n4768 = n4750 ^ x23 ^ 1'b0 ;
  assign n4769 = x79 & ~n4605 ;
  assign n4770 = ( x79 & n4766 ) | ( x79 & ~n4769 ) | ( n4766 & ~n4769 ) ;
  assign n4771 = n1216 & n4608 ;
  assign n4772 = n4770 | n4771 ;
  assign n4773 = n4772 ^ x23 ^ 1'b0 ;
  assign n4774 = n4768 ^ n4762 ^ n3856 ;
  assign n4775 = ( n3856 & n4762 ) | ( n3856 & n4768 ) | ( n4762 & n4768 ) ;
  assign n4776 = ( n3866 & n4773 ) | ( n3866 & n4775 ) | ( n4773 & n4775 ) ;
  assign n4777 = n4776 ^ n4767 ^ n3876 ;
  assign n4778 = ( n3876 & n4767 ) | ( n3876 & n4776 ) | ( n4767 & n4776 ) ;
  assign n4779 = n4775 ^ n4773 ^ n3866 ;
  assign n4780 = x13 ^ x12 ^ 1'b0 ;
  assign n4781 = x12 ^ x11 ^ 1'b0 ;
  assign n4782 = x19 ^ x18 ^ 1'b0 ;
  assign n4783 = x14 ^ x13 ^ 1'b0 ;
  assign n4784 = x20 ^ x19 ^ 1'b0 ;
  assign n4785 = x18 ^ x17 ^ 1'b0 ;
  assign n4786 = n4782 & ~n4785 ;
  assign n4787 = n4784 & n4785 ;
  assign n4788 = ( n4782 & n4784 ) | ( n4782 & ~n4785 ) | ( n4784 & ~n4785 ) ;
  assign n4789 = x64 & n4786 ;
  assign n4790 = ~n4782 & n4788 ;
  assign n4791 = ( n190 & n4787 ) | ( n190 & n4789 ) | ( n4787 & n4789 ) ;
  assign n4792 = ~n4784 & n4785 ;
  assign n4793 = x65 & n4790 ;
  assign n4794 = ~x65 & n4792 ;
  assign n4795 = ( n4789 & n4792 ) | ( n4789 & ~n4794 ) | ( n4792 & ~n4794 ) ;
  assign n4796 = n4791 | n4795 ;
  assign n4797 = ( x67 & n4792 ) | ( x67 & n4793 ) | ( n4792 & n4793 ) ;
  assign n4798 = n4793 | n4797 ;
  assign n4799 = x66 & ~n4786 ;
  assign n4800 = ( x66 & n4798 ) | ( x66 & ~n4799 ) | ( n4798 & ~n4799 ) ;
  assign n4801 = n161 & n4787 ;
  assign n4802 = n4800 | n4801 ;
  assign n4803 = x64 & n4785 ;
  assign n4804 = x20 & ~n4803 ;
  assign n4805 = x64 & n4790 ;
  assign n4806 = ( x66 & n4792 ) | ( x66 & n4805 ) | ( n4792 & n4805 ) ;
  assign n4807 = n4805 | n4806 ;
  assign n4808 = x65 & ~n4786 ;
  assign n4809 = ( x65 & n4807 ) | ( x65 & ~n4808 ) | ( n4807 & ~n4808 ) ;
  assign n4810 = n139 & n4787 ;
  assign n4811 = n4809 | n4810 ;
  assign n4812 = n4802 ^ x20 ^ 1'b0 ;
  assign n4813 = n4796 ^ x20 ^ 1'b0 ;
  assign n4814 = n4804 & n4813 ;
  assign n4815 = n4811 ^ x20 ^ 1'b0 ;
  assign n4816 = n4813 ^ n4804 ^ 1'b0 ;
  assign n4817 = n4814 & n4815 ;
  assign n4818 = n4815 ^ n4814 ^ 1'b0 ;
  assign n4819 = n4817 ^ n4812 ^ n4620 ;
  assign n4820 = ( n4620 & n4812 ) | ( n4620 & n4817 ) | ( n4812 & n4817 ) ;
  assign n4821 = x66 & n4790 ;
  assign n4822 = ( x68 & n4792 ) | ( x68 & n4821 ) | ( n4792 & n4821 ) ;
  assign n4823 = n4821 | n4822 ;
  assign n4824 = x67 & ~n4786 ;
  assign n4825 = ( x67 & n4823 ) | ( x67 & ~n4824 ) | ( n4823 & ~n4824 ) ;
  assign n4826 = n175 & n4787 ;
  assign n4827 = n4825 | n4826 ;
  assign n4828 = n4827 ^ x20 ^ 1'b0 ;
  assign n4829 = n4828 ^ n4820 ^ n4629 ;
  assign n4830 = ( n4629 & n4820 ) | ( n4629 & n4828 ) | ( n4820 & n4828 ) ;
  assign n4831 = x67 & n4790 ;
  assign n4832 = ( x69 & n4792 ) | ( x69 & n4831 ) | ( n4792 & n4831 ) ;
  assign n4833 = n4831 | n4832 ;
  assign n4834 = x68 & ~n4786 ;
  assign n4835 = ( x68 & n4833 ) | ( x68 & ~n4834 ) | ( n4833 & ~n4834 ) ;
  assign n4836 = n172 & n4787 ;
  assign n4837 = n4835 | n4836 ;
  assign n4838 = n4837 ^ x20 ^ 1'b0 ;
  assign n4839 = n4838 ^ n4830 ^ n4627 ;
  assign n4840 = ( n4627 & n4830 ) | ( n4627 & n4838 ) | ( n4830 & n4838 ) ;
  assign n4841 = x68 & n4790 ;
  assign n4842 = ( x70 & n4792 ) | ( x70 & n4841 ) | ( n4792 & n4841 ) ;
  assign n4843 = n4841 | n4842 ;
  assign n4844 = x69 & ~n4786 ;
  assign n4845 = ( x69 & n4843 ) | ( x69 & ~n4844 ) | ( n4843 & ~n4844 ) ;
  assign n4846 = n168 & n4787 ;
  assign n4847 = n4845 | n4846 ;
  assign n4848 = n4847 ^ x20 ^ 1'b0 ;
  assign n4849 = n4848 ^ n4840 ^ n4639 ;
  assign n4850 = ( n4639 & n4840 ) | ( n4639 & n4848 ) | ( n4840 & n4848 ) ;
  assign n4851 = x69 & n4790 ;
  assign n4852 = ( x71 & n4792 ) | ( x71 & n4851 ) | ( n4792 & n4851 ) ;
  assign n4853 = n4851 | n4852 ;
  assign n4854 = x70 & ~n4786 ;
  assign n4855 = ( x70 & n4853 ) | ( x70 & ~n4854 ) | ( n4853 & ~n4854 ) ;
  assign n4856 = n328 & n4787 ;
  assign n4857 = n4855 | n4856 ;
  assign n4858 = n4857 ^ x20 ^ 1'b0 ;
  assign n4859 = ( n4648 & n4850 ) | ( n4648 & n4858 ) | ( n4850 & n4858 ) ;
  assign n4860 = n4858 ^ n4850 ^ n4648 ;
  assign n4861 = x70 & n4790 ;
  assign n4862 = ( x72 & n4792 ) | ( x72 & n4861 ) | ( n4792 & n4861 ) ;
  assign n4863 = n4861 | n4862 ;
  assign n4864 = x71 & ~n4786 ;
  assign n4865 = ( x71 & n4863 ) | ( x71 & ~n4864 ) | ( n4863 & ~n4864 ) ;
  assign n4866 = n349 & n4787 ;
  assign n4867 = n4865 | n4866 ;
  assign n4868 = n4867 ^ x20 ^ 1'b0 ;
  assign n4869 = n4868 ^ n4859 ^ n4658 ;
  assign n4870 = ( n4658 & n4859 ) | ( n4658 & n4868 ) | ( n4859 & n4868 ) ;
  assign n4871 = x71 & n4790 ;
  assign n4872 = ( x73 & n4792 ) | ( x73 & n4871 ) | ( n4792 & n4871 ) ;
  assign n4873 = n4871 | n4872 ;
  assign n4874 = x72 & ~n4786 ;
  assign n4875 = ( x72 & n4873 ) | ( x72 & ~n4874 ) | ( n4873 & ~n4874 ) ;
  assign n4876 = n370 & n4787 ;
  assign n4877 = n4875 | n4876 ;
  assign n4878 = n4877 ^ x20 ^ 1'b0 ;
  assign n4879 = n4878 ^ n4870 ^ n4668 ;
  assign n4880 = ( n4668 & n4870 ) | ( n4668 & n4878 ) | ( n4870 & n4878 ) ;
  assign n4881 = x72 & n4790 ;
  assign n4882 = ( x74 & n4792 ) | ( x74 & n4881 ) | ( n4792 & n4881 ) ;
  assign n4883 = n4881 | n4882 ;
  assign n4884 = x73 & ~n4786 ;
  assign n4885 = ( x73 & n4883 ) | ( x73 & ~n4884 ) | ( n4883 & ~n4884 ) ;
  assign n4886 = n504 & n4787 ;
  assign n4887 = n4885 | n4886 ;
  assign n4888 = n4887 ^ x20 ^ 1'b0 ;
  assign n4889 = n4888 ^ n4880 ^ n4678 ;
  assign n4890 = ( n4678 & n4880 ) | ( n4678 & n4888 ) | ( n4880 & n4888 ) ;
  assign n4891 = x73 & n4790 ;
  assign n4892 = ( x75 & n4792 ) | ( x75 & n4891 ) | ( n4792 & n4891 ) ;
  assign n4893 = n4891 | n4892 ;
  assign n4894 = x74 & ~n4786 ;
  assign n4895 = ( x74 & n4893 ) | ( x74 & ~n4894 ) | ( n4893 & ~n4894 ) ;
  assign n4896 = n525 & n4787 ;
  assign n4897 = n4895 | n4896 ;
  assign n4898 = n4897 ^ x20 ^ 1'b0 ;
  assign n4899 = n4898 ^ n4890 ^ n4689 ;
  assign n4900 = ( n4689 & n4890 ) | ( n4689 & n4898 ) | ( n4890 & n4898 ) ;
  assign n4901 = x74 & n4790 ;
  assign n4902 = ( x76 & n4792 ) | ( x76 & n4901 ) | ( n4792 & n4901 ) ;
  assign n4903 = n4901 | n4902 ;
  assign n4904 = x75 & ~n4786 ;
  assign n4905 = ( x75 & n4903 ) | ( x75 & ~n4904 ) | ( n4903 & ~n4904 ) ;
  assign n4906 = n664 & n4787 ;
  assign n4907 = n4905 | n4906 ;
  assign n4908 = n4907 ^ x20 ^ 1'b0 ;
  assign n4909 = ( n4699 & n4900 ) | ( n4699 & n4908 ) | ( n4900 & n4908 ) ;
  assign n4910 = n4908 ^ n4900 ^ n4699 ;
  assign n4911 = x75 & n4790 ;
  assign n4912 = ( x77 & n4792 ) | ( x77 & n4911 ) | ( n4792 & n4911 ) ;
  assign n4913 = n4911 | n4912 ;
  assign n4914 = x76 & ~n4786 ;
  assign n4915 = ( x76 & n4913 ) | ( x76 & ~n4914 ) | ( n4913 & ~n4914 ) ;
  assign n4916 = n690 & n4787 ;
  assign n4917 = n4915 | n4916 ;
  assign n4918 = n4917 ^ x20 ^ 1'b0 ;
  assign n4919 = n4918 ^ n4909 ^ n4708 ;
  assign n4920 = ( n4708 & n4909 ) | ( n4708 & n4918 ) | ( n4909 & n4918 ) ;
  assign n4921 = x76 & n4790 ;
  assign n4922 = ( x78 & n4792 ) | ( x78 & n4921 ) | ( n4792 & n4921 ) ;
  assign n4923 = n4921 | n4922 ;
  assign n4924 = x77 & ~n4786 ;
  assign n4925 = ( x77 & n4923 ) | ( x77 & ~n4924 ) | ( n4923 & ~n4924 ) ;
  assign n4926 = n709 & n4787 ;
  assign n4927 = n4925 | n4926 ;
  assign n4928 = n4927 ^ x20 ^ 1'b0 ;
  assign n4929 = ( n4718 & n4920 ) | ( n4718 & n4928 ) | ( n4920 & n4928 ) ;
  assign n4930 = n4928 ^ n4920 ^ n4718 ;
  assign n4931 = x77 & n4790 ;
  assign n4932 = ( x79 & n4792 ) | ( x79 & n4931 ) | ( n4792 & n4931 ) ;
  assign n4933 = n4931 | n4932 ;
  assign n4934 = x78 & ~n4786 ;
  assign n4935 = ( x78 & n4933 ) | ( x78 & ~n4934 ) | ( n4933 & ~n4934 ) ;
  assign n4936 = n1015 & n4787 ;
  assign n4937 = n4935 | n4936 ;
  assign n4938 = n4937 ^ x20 ^ 1'b0 ;
  assign n4939 = ( n4729 & n4929 ) | ( n4729 & n4938 ) | ( n4929 & n4938 ) ;
  assign n4940 = n4938 ^ n4929 ^ n4729 ;
  assign n4941 = x78 & n4790 ;
  assign n4942 = ( x80 & n4792 ) | ( x80 & n4941 ) | ( n4792 & n4941 ) ;
  assign n4943 = n4941 | n4942 ;
  assign n4944 = x79 & ~n4786 ;
  assign n4945 = ( x79 & n4943 ) | ( x79 & ~n4944 ) | ( n4943 & ~n4944 ) ;
  assign n4946 = n1216 & n4787 ;
  assign n4947 = n4945 | n4946 ;
  assign n4948 = n4947 ^ x20 ^ 1'b0 ;
  assign n4949 = n4948 ^ n4939 ^ n4738 ;
  assign n4950 = ( n4738 & n4939 ) | ( n4738 & n4948 ) | ( n4939 & n4948 ) ;
  assign n4951 = x79 & n4790 ;
  assign n4952 = x80 & ~n4786 ;
  assign n4953 = x81 & ~n4786 ;
  assign n4954 = ( x81 & n4792 ) | ( x81 & n4951 ) | ( n4792 & n4951 ) ;
  assign n4955 = n4951 | n4954 ;
  assign n4956 = n1258 & n4787 ;
  assign n4957 = ( x80 & ~n4952 ) | ( x80 & n4955 ) | ( ~n4952 & n4955 ) ;
  assign n4958 = x80 & n4790 ;
  assign n4959 = n4956 | n4957 ;
  assign n4960 = ( x82 & n4792 ) | ( x82 & n4958 ) | ( n4792 & n4958 ) ;
  assign n4961 = n4958 | n4960 ;
  assign n4962 = ( x81 & ~n4953 ) | ( x81 & n4961 ) | ( ~n4953 & n4961 ) ;
  assign n4963 = n4959 ^ x20 ^ 1'b0 ;
  assign n4964 = n1301 & n4787 ;
  assign n4965 = n4962 | n4964 ;
  assign n4966 = n4965 ^ x20 ^ 1'b0 ;
  assign n4967 = ( n4763 & n4950 ) | ( n4763 & n4963 ) | ( n4950 & n4963 ) ;
  assign n4968 = n4967 ^ n4966 ^ n4774 ;
  assign n4969 = ( n4774 & n4966 ) | ( n4774 & n4967 ) | ( n4966 & n4967 ) ;
  assign n4970 = n1329 & n4787 ;
  assign n4971 = ( n4780 & ~n4781 ) | ( n4780 & n4783 ) | ( ~n4781 & n4783 ) ;
  assign n4972 = ~n4780 & n4971 ;
  assign n4973 = n4963 ^ n4950 ^ n4763 ;
  assign n4974 = x81 & n4790 ;
  assign n4975 = ( x83 & n4792 ) | ( x83 & n4974 ) | ( n4792 & n4974 ) ;
  assign n4976 = n4974 | n4975 ;
  assign n4977 = x82 & ~n4786 ;
  assign n4978 = ( x82 & n4976 ) | ( x82 & ~n4977 ) | ( n4976 & ~n4977 ) ;
  assign n4979 = x82 & n4790 ;
  assign n4980 = n4780 & ~n4781 ;
  assign n4981 = n4970 | n4978 ;
  assign n4982 = n4981 ^ x20 ^ 1'b0 ;
  assign n4983 = n4982 ^ n4969 ^ n4779 ;
  assign n4984 = ( n4779 & n4969 ) | ( n4779 & n4982 ) | ( n4969 & n4982 ) ;
  assign n4985 = n4781 & ~n4783 ;
  assign n4986 = ( x84 & n4792 ) | ( x84 & n4979 ) | ( n4792 & n4979 ) ;
  assign n4987 = n4781 & n4783 ;
  assign n4988 = n4979 | n4986 ;
  assign n4989 = x83 & ~n4786 ;
  assign n4990 = ( x83 & n4988 ) | ( x83 & ~n4989 ) | ( n4988 & ~n4989 ) ;
  assign n4991 = n1355 & n4787 ;
  assign n4992 = n4990 | n4991 ;
  assign n4993 = n4992 ^ x20 ^ 1'b0 ;
  assign n4994 = n4993 ^ n4984 ^ n4777 ;
  assign n4995 = x64 & n4781 ;
  assign n4996 = ( n4777 & n4984 ) | ( n4777 & n4993 ) | ( n4984 & n4993 ) ;
  assign n4997 = x67 & n4972 ;
  assign n4998 = ( x69 & n4985 ) | ( x69 & n4997 ) | ( n4985 & n4997 ) ;
  assign n4999 = n4997 | n4998 ;
  assign n5000 = x68 & ~n4980 ;
  assign n5001 = ( x68 & n4999 ) | ( x68 & ~n5000 ) | ( n4999 & ~n5000 ) ;
  assign n5002 = n172 & n4987 ;
  assign n5003 = n5001 | n5002 ;
  assign n5004 = n5003 ^ x14 ^ 1'b0 ;
  assign n5005 = x17 ^ x16 ^ 1'b0 ;
  assign n5006 = x15 ^ x14 ^ 1'b0 ;
  assign n5007 = x16 ^ x15 ^ 1'b0 ;
  assign n5008 = ~n5006 & n5007 ;
  assign n5009 = x64 & n5008 ;
  assign n5010 = ( n5005 & ~n5006 ) | ( n5005 & n5007 ) | ( ~n5006 & n5007 ) ;
  assign n5011 = ~n5007 & n5010 ;
  assign n5012 = ~n5005 & n5006 ;
  assign n5013 = ~x65 & n5012 ;
  assign n5014 = x64 & n5011 ;
  assign n5015 = ( x66 & n5012 ) | ( x66 & n5014 ) | ( n5012 & n5014 ) ;
  assign n5016 = n5014 | n5015 ;
  assign n5017 = ( n5009 & n5012 ) | ( n5009 & ~n5013 ) | ( n5012 & ~n5013 ) ;
  assign n5018 = x65 & ~n5008 ;
  assign n5019 = ( x65 & n5016 ) | ( x65 & ~n5018 ) | ( n5016 & ~n5018 ) ;
  assign n5020 = n5005 & n5006 ;
  assign n5021 = x64 & n5006 ;
  assign n5022 = ( n190 & n5009 ) | ( n190 & n5020 ) | ( n5009 & n5020 ) ;
  assign n5023 = n139 & n5020 ;
  assign n5024 = n5019 | n5023 ;
  assign n5025 = n5017 | n5022 ;
  assign n5026 = x17 & ~n5021 ;
  assign n5027 = n5025 ^ x17 ^ 1'b0 ;
  assign n5028 = x65 & n5011 ;
  assign n5029 = ( x67 & n5012 ) | ( x67 & n5028 ) | ( n5012 & n5028 ) ;
  assign n5030 = n5028 | n5029 ;
  assign n5031 = n5026 & n5027 ;
  assign n5032 = n5024 ^ x17 ^ 1'b0 ;
  assign n5033 = n5027 ^ n5026 ^ 1'b0 ;
  assign n5034 = n5031 & n5032 ;
  assign n5035 = n5032 ^ n5031 ^ 1'b0 ;
  assign n5036 = x66 & ~n5008 ;
  assign n5037 = ( x66 & n5030 ) | ( x66 & ~n5036 ) | ( n5030 & ~n5036 ) ;
  assign n5038 = n161 & n5020 ;
  assign n5039 = n5037 | n5038 ;
  assign n5040 = n5039 ^ x17 ^ 1'b0 ;
  assign n5041 = ( n4803 & n5034 ) | ( n4803 & n5040 ) | ( n5034 & n5040 ) ;
  assign n5042 = n5040 ^ n5034 ^ n4803 ;
  assign n5043 = x66 & n5011 ;
  assign n5044 = ( x68 & n5012 ) | ( x68 & n5043 ) | ( n5012 & n5043 ) ;
  assign n5045 = n5043 | n5044 ;
  assign n5046 = x67 & ~n5008 ;
  assign n5047 = ( x67 & n5045 ) | ( x67 & ~n5046 ) | ( n5045 & ~n5046 ) ;
  assign n5048 = n175 & n5020 ;
  assign n5049 = n5047 | n5048 ;
  assign n5050 = n5049 ^ x17 ^ 1'b0 ;
  assign n5051 = n5050 ^ n5041 ^ n4816 ;
  assign n5052 = ( n4816 & n5041 ) | ( n4816 & n5050 ) | ( n5041 & n5050 ) ;
  assign n5053 = x67 & n5011 ;
  assign n5054 = ( x69 & n5012 ) | ( x69 & n5053 ) | ( n5012 & n5053 ) ;
  assign n5055 = n5053 | n5054 ;
  assign n5056 = x68 & ~n5008 ;
  assign n5057 = ( x68 & n5055 ) | ( x68 & ~n5056 ) | ( n5055 & ~n5056 ) ;
  assign n5058 = n172 & n5020 ;
  assign n5059 = n5057 | n5058 ;
  assign n5060 = n5059 ^ x17 ^ 1'b0 ;
  assign n5061 = ( n4818 & n5052 ) | ( n4818 & n5060 ) | ( n5052 & n5060 ) ;
  assign n5062 = n5060 ^ n5052 ^ n4818 ;
  assign n5063 = x68 & n5011 ;
  assign n5064 = ( x70 & n5012 ) | ( x70 & n5063 ) | ( n5012 & n5063 ) ;
  assign n5065 = n5063 | n5064 ;
  assign n5066 = x69 & ~n5008 ;
  assign n5067 = ( x69 & n5065 ) | ( x69 & ~n5066 ) | ( n5065 & ~n5066 ) ;
  assign n5068 = n168 & n5020 ;
  assign n5069 = n5067 | n5068 ;
  assign n5070 = n5069 ^ x17 ^ 1'b0 ;
  assign n5071 = n5070 ^ n5061 ^ n4819 ;
  assign n5072 = ( n4819 & n5061 ) | ( n4819 & n5070 ) | ( n5061 & n5070 ) ;
  assign n5073 = x69 & n5011 ;
  assign n5074 = ( x71 & n5012 ) | ( x71 & n5073 ) | ( n5012 & n5073 ) ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = x70 & ~n5008 ;
  assign n5077 = ( x70 & n5075 ) | ( x70 & ~n5076 ) | ( n5075 & ~n5076 ) ;
  assign n5078 = n328 & n5020 ;
  assign n5079 = n5077 | n5078 ;
  assign n5080 = n5079 ^ x17 ^ 1'b0 ;
  assign n5081 = n5080 ^ n5072 ^ n4829 ;
  assign n5082 = ( n4829 & n5072 ) | ( n4829 & n5080 ) | ( n5072 & n5080 ) ;
  assign n5083 = x70 & n5011 ;
  assign n5084 = ( x72 & n5012 ) | ( x72 & n5083 ) | ( n5012 & n5083 ) ;
  assign n5085 = n5083 | n5084 ;
  assign n5086 = x71 & ~n5008 ;
  assign n5087 = ( x71 & n5085 ) | ( x71 & ~n5086 ) | ( n5085 & ~n5086 ) ;
  assign n5088 = n349 & n5020 ;
  assign n5089 = n5087 | n5088 ;
  assign n5090 = n5089 ^ x17 ^ 1'b0 ;
  assign n5091 = ( n4839 & n5082 ) | ( n4839 & n5090 ) | ( n5082 & n5090 ) ;
  assign n5092 = n5090 ^ n5082 ^ n4839 ;
  assign n5093 = x71 & n5011 ;
  assign n5094 = ( x73 & n5012 ) | ( x73 & n5093 ) | ( n5012 & n5093 ) ;
  assign n5095 = n5093 | n5094 ;
  assign n5096 = x72 & ~n5008 ;
  assign n5097 = ( x72 & n5095 ) | ( x72 & ~n5096 ) | ( n5095 & ~n5096 ) ;
  assign n5098 = n370 & n5020 ;
  assign n5099 = n5097 | n5098 ;
  assign n5100 = n5099 ^ x17 ^ 1'b0 ;
  assign n5101 = n5100 ^ n5091 ^ n4849 ;
  assign n5102 = ( n4849 & n5091 ) | ( n4849 & n5100 ) | ( n5091 & n5100 ) ;
  assign n5103 = x72 & n5011 ;
  assign n5104 = ( x74 & n5012 ) | ( x74 & n5103 ) | ( n5012 & n5103 ) ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = x73 & ~n5008 ;
  assign n5107 = ( x73 & n5105 ) | ( x73 & ~n5106 ) | ( n5105 & ~n5106 ) ;
  assign n5108 = n504 & n5020 ;
  assign n5109 = n5107 | n5108 ;
  assign n5110 = n5109 ^ x17 ^ 1'b0 ;
  assign n5111 = ( n4860 & n5102 ) | ( n4860 & n5110 ) | ( n5102 & n5110 ) ;
  assign n5112 = n5110 ^ n5102 ^ n4860 ;
  assign n5113 = x73 & n5011 ;
  assign n5114 = ( x75 & n5012 ) | ( x75 & n5113 ) | ( n5012 & n5113 ) ;
  assign n5115 = n5113 | n5114 ;
  assign n5116 = x74 & ~n5008 ;
  assign n5117 = ( x74 & n5115 ) | ( x74 & ~n5116 ) | ( n5115 & ~n5116 ) ;
  assign n5118 = n525 & n5020 ;
  assign n5119 = n5117 | n5118 ;
  assign n5120 = n5119 ^ x17 ^ 1'b0 ;
  assign n5121 = ( n4869 & n5111 ) | ( n4869 & n5120 ) | ( n5111 & n5120 ) ;
  assign n5122 = n5120 ^ n5111 ^ n4869 ;
  assign n5123 = x74 & n5011 ;
  assign n5124 = ( x76 & n5012 ) | ( x76 & n5123 ) | ( n5012 & n5123 ) ;
  assign n5125 = n5123 | n5124 ;
  assign n5126 = x75 & ~n5008 ;
  assign n5127 = ( x75 & n5125 ) | ( x75 & ~n5126 ) | ( n5125 & ~n5126 ) ;
  assign n5128 = n664 & n5020 ;
  assign n5129 = n5127 | n5128 ;
  assign n5130 = n5129 ^ x17 ^ 1'b0 ;
  assign n5131 = n5130 ^ n5121 ^ n4879 ;
  assign n5132 = ( n4879 & n5121 ) | ( n4879 & n5130 ) | ( n5121 & n5130 ) ;
  assign n5133 = x75 & n5011 ;
  assign n5134 = ( x77 & n5012 ) | ( x77 & n5133 ) | ( n5012 & n5133 ) ;
  assign n5135 = n5133 | n5134 ;
  assign n5136 = x76 & ~n5008 ;
  assign n5137 = ( x76 & n5135 ) | ( x76 & ~n5136 ) | ( n5135 & ~n5136 ) ;
  assign n5138 = n690 & n5020 ;
  assign n5139 = n5137 | n5138 ;
  assign n5140 = n5139 ^ x17 ^ 1'b0 ;
  assign n5141 = ( n4889 & n5132 ) | ( n4889 & n5140 ) | ( n5132 & n5140 ) ;
  assign n5142 = n5140 ^ n5132 ^ n4889 ;
  assign n5143 = x76 & n5011 ;
  assign n5144 = ( x78 & n5012 ) | ( x78 & n5143 ) | ( n5012 & n5143 ) ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = x77 & ~n5008 ;
  assign n5147 = ( x77 & n5145 ) | ( x77 & ~n5146 ) | ( n5145 & ~n5146 ) ;
  assign n5148 = n709 & n5020 ;
  assign n5149 = n5147 | n5148 ;
  assign n5150 = n5149 ^ x17 ^ 1'b0 ;
  assign n5151 = n5150 ^ n5141 ^ n4899 ;
  assign n5152 = ( n4899 & n5141 ) | ( n4899 & n5150 ) | ( n5141 & n5150 ) ;
  assign n5153 = x77 & n5011 ;
  assign n5154 = ( x79 & n5012 ) | ( x79 & n5153 ) | ( n5012 & n5153 ) ;
  assign n5155 = n5153 | n5154 ;
  assign n5156 = x78 & ~n5008 ;
  assign n5157 = ( x78 & n5155 ) | ( x78 & ~n5156 ) | ( n5155 & ~n5156 ) ;
  assign n5158 = n1015 & n5020 ;
  assign n5159 = n5157 | n5158 ;
  assign n5160 = n5159 ^ x17 ^ 1'b0 ;
  assign n5161 = ( n4910 & n5152 ) | ( n4910 & n5160 ) | ( n5152 & n5160 ) ;
  assign n5162 = n5160 ^ n5152 ^ n4910 ;
  assign n5163 = x78 & n5011 ;
  assign n5164 = ( x80 & n5012 ) | ( x80 & n5163 ) | ( n5012 & n5163 ) ;
  assign n5165 = n5163 | n5164 ;
  assign n5166 = x79 & ~n5008 ;
  assign n5167 = ( x79 & n5165 ) | ( x79 & ~n5166 ) | ( n5165 & ~n5166 ) ;
  assign n5168 = n1216 & n5020 ;
  assign n5169 = n5167 | n5168 ;
  assign n5170 = n5169 ^ x17 ^ 1'b0 ;
  assign n5171 = n5170 ^ n5161 ^ n4919 ;
  assign n5172 = ( n4919 & n5161 ) | ( n4919 & n5170 ) | ( n5161 & n5170 ) ;
  assign n5173 = x79 & n5011 ;
  assign n5174 = ( x81 & n5012 ) | ( x81 & n5173 ) | ( n5012 & n5173 ) ;
  assign n5175 = n5173 | n5174 ;
  assign n5176 = x80 & ~n5008 ;
  assign n5177 = ( x80 & n5175 ) | ( x80 & ~n5176 ) | ( n5175 & ~n5176 ) ;
  assign n5178 = n1258 & n5020 ;
  assign n5179 = n5177 | n5178 ;
  assign n5180 = n5179 ^ x17 ^ 1'b0 ;
  assign n5181 = ( n4930 & n5172 ) | ( n4930 & n5180 ) | ( n5172 & n5180 ) ;
  assign n5182 = n5180 ^ n5172 ^ n4930 ;
  assign n5183 = x80 & n5011 ;
  assign n5184 = ( x82 & n5012 ) | ( x82 & n5183 ) | ( n5012 & n5183 ) ;
  assign n5185 = n5183 | n5184 ;
  assign n5186 = x81 & ~n5008 ;
  assign n5187 = ( x81 & n5185 ) | ( x81 & ~n5186 ) | ( n5185 & ~n5186 ) ;
  assign n5188 = n1301 & n5020 ;
  assign n5189 = n5187 | n5188 ;
  assign n5190 = n5189 ^ x17 ^ 1'b0 ;
  assign n5191 = n5190 ^ n5181 ^ n4940 ;
  assign n5192 = ( n4940 & n5181 ) | ( n4940 & n5190 ) | ( n5181 & n5190 ) ;
  assign n5193 = x81 & n5011 ;
  assign n5194 = ( x83 & n5012 ) | ( x83 & n5193 ) | ( n5012 & n5193 ) ;
  assign n5195 = n5193 | n5194 ;
  assign n5196 = x82 & ~n5008 ;
  assign n5197 = ( x82 & n5195 ) | ( x82 & ~n5196 ) | ( n5195 & ~n5196 ) ;
  assign n5198 = n1329 & n5020 ;
  assign n5199 = n5197 | n5198 ;
  assign n5200 = n5199 ^ x17 ^ 1'b0 ;
  assign n5201 = n5200 ^ n5192 ^ n4949 ;
  assign n5202 = ( n4949 & n5192 ) | ( n4949 & n5200 ) | ( n5192 & n5200 ) ;
  assign n5203 = x82 & n5011 ;
  assign n5204 = ( x84 & n5012 ) | ( x84 & n5203 ) | ( n5012 & n5203 ) ;
  assign n5205 = n5203 | n5204 ;
  assign n5206 = x83 & ~n5008 ;
  assign n5207 = ( x83 & n5205 ) | ( x83 & ~n5206 ) | ( n5205 & ~n5206 ) ;
  assign n5208 = n1355 & n5020 ;
  assign n5209 = n5207 | n5208 ;
  assign n5210 = n5209 ^ x17 ^ 1'b0 ;
  assign n5211 = n5210 ^ n5202 ^ n4973 ;
  assign n5212 = ( n4973 & n5202 ) | ( n4973 & n5210 ) | ( n5202 & n5210 ) ;
  assign n5213 = x83 & n5011 ;
  assign n5214 = ( x85 & n5012 ) | ( x85 & n5213 ) | ( n5012 & n5213 ) ;
  assign n5215 = n5213 | n5214 ;
  assign n5216 = x84 & ~n5008 ;
  assign n5217 = ( x84 & n5215 ) | ( x84 & ~n5216 ) | ( n5215 & ~n5216 ) ;
  assign n5218 = n1392 & n5020 ;
  assign n5219 = n5217 | n5218 ;
  assign n5220 = n5219 ^ x17 ^ 1'b0 ;
  assign n5221 = ( n4968 & n5212 ) | ( n4968 & n5220 ) | ( n5212 & n5220 ) ;
  assign n5222 = n5220 ^ n5212 ^ n4968 ;
  assign n5223 = x84 & n5011 ;
  assign n5224 = ( x86 & n5012 ) | ( x86 & n5223 ) | ( n5012 & n5223 ) ;
  assign n5225 = n5223 | n5224 ;
  assign n5226 = x85 & ~n5008 ;
  assign n5227 = ( x85 & n5225 ) | ( x85 & ~n5226 ) | ( n5225 & ~n5226 ) ;
  assign n5228 = n1419 & n5020 ;
  assign n5229 = n5227 | n5228 ;
  assign n5230 = n5229 ^ x17 ^ 1'b0 ;
  assign n5231 = ( n4983 & n5221 ) | ( n4983 & n5230 ) | ( n5221 & n5230 ) ;
  assign n5232 = n5230 ^ n5221 ^ n4983 ;
  assign n5233 = x85 & n5011 ;
  assign n5234 = ( x87 & n5012 ) | ( x87 & n5233 ) | ( n5012 & n5233 ) ;
  assign n5235 = n5233 | n5234 ;
  assign n5236 = x86 & ~n5008 ;
  assign n5237 = ( x86 & n5235 ) | ( x86 & ~n5236 ) | ( n5235 & ~n5236 ) ;
  assign n5238 = n1484 & n5020 ;
  assign n5239 = n5237 | n5238 ;
  assign n5240 = n5239 ^ x17 ^ 1'b0 ;
  assign n5241 = n5240 ^ n5231 ^ n4994 ;
  assign n5242 = ( n4994 & n5231 ) | ( n4994 & n5240 ) | ( n5231 & n5240 ) ;
  assign n5243 = x64 & n4972 ;
  assign n5244 = ~x65 & n4985 ;
  assign n5245 = x64 & n4980 ;
  assign n5246 = ( n4985 & ~n5244 ) | ( n4985 & n5245 ) | ( ~n5244 & n5245 ) ;
  assign n5247 = ( x66 & n4985 ) | ( x66 & n5243 ) | ( n4985 & n5243 ) ;
  assign n5248 = x65 & ~n4980 ;
  assign n5249 = n5243 | n5247 ;
  assign n5250 = ( x65 & ~n5248 ) | ( x65 & n5249 ) | ( ~n5248 & n5249 ) ;
  assign n5251 = n139 & n4987 ;
  assign n5252 = n5250 | n5251 ;
  assign n5253 = x14 & ~n4995 ;
  assign n5254 = n5252 ^ x14 ^ 1'b0 ;
  assign n5255 = ( n190 & n4987 ) | ( n190 & n5245 ) | ( n4987 & n5245 ) ;
  assign n5256 = n5246 | n5255 ;
  assign n5257 = n5256 ^ x14 ^ 1'b0 ;
  assign n5258 = n5253 & n5257 ;
  assign n5259 = n5254 & n5258 ;
  assign n5260 = n5257 ^ n5253 ^ 1'b0 ;
  assign n5261 = x65 & n4972 ;
  assign n5262 = n5258 ^ n5254 ^ 1'b0 ;
  assign n5263 = ( x67 & n4985 ) | ( x67 & n5261 ) | ( n4985 & n5261 ) ;
  assign n5264 = n5261 | n5263 ;
  assign n5265 = x66 & ~n4980 ;
  assign n5266 = ( x66 & n5264 ) | ( x66 & ~n5265 ) | ( n5264 & ~n5265 ) ;
  assign n5267 = n161 & n4987 ;
  assign n5268 = n5266 | n5267 ;
  assign n5269 = n5268 ^ x14 ^ 1'b0 ;
  assign n5270 = ( n5021 & n5259 ) | ( n5021 & n5269 ) | ( n5259 & n5269 ) ;
  assign n5271 = n5269 ^ n5259 ^ n5021 ;
  assign n5272 = x66 & n4972 ;
  assign n5273 = ( x68 & n4985 ) | ( x68 & n5272 ) | ( n4985 & n5272 ) ;
  assign n5274 = n5272 | n5273 ;
  assign n5275 = x67 & ~n4980 ;
  assign n5276 = ( x67 & n5274 ) | ( x67 & ~n5275 ) | ( n5274 & ~n5275 ) ;
  assign n5277 = n175 & n4987 ;
  assign n5278 = n5276 | n5277 ;
  assign n5279 = n5278 ^ x14 ^ 1'b0 ;
  assign n5280 = ( n5033 & n5270 ) | ( n5033 & n5279 ) | ( n5270 & n5279 ) ;
  assign n5281 = n5279 ^ n5270 ^ n5033 ;
  assign n5282 = x70 & n4972 ;
  assign n5283 = ( x72 & n4985 ) | ( x72 & n5282 ) | ( n4985 & n5282 ) ;
  assign n5284 = n5282 | n5283 ;
  assign n5285 = x71 & ~n4980 ;
  assign n5286 = ( x71 & n5284 ) | ( x71 & ~n5285 ) | ( n5284 & ~n5285 ) ;
  assign n5287 = n349 & n4987 ;
  assign n5288 = n5286 | n5287 ;
  assign n5289 = ( n5004 & n5035 ) | ( n5004 & n5280 ) | ( n5035 & n5280 ) ;
  assign n5290 = n5280 ^ n5035 ^ n5004 ;
  assign n5291 = n5288 ^ x14 ^ 1'b0 ;
  assign n5292 = x68 & n4972 ;
  assign n5293 = ( x70 & n4985 ) | ( x70 & n5292 ) | ( n4985 & n5292 ) ;
  assign n5294 = n5292 | n5293 ;
  assign n5295 = x69 & ~n4980 ;
  assign n5296 = ( x69 & n5294 ) | ( x69 & ~n5295 ) | ( n5294 & ~n5295 ) ;
  assign n5297 = n168 & n4987 ;
  assign n5298 = n5296 | n5297 ;
  assign n5299 = n5298 ^ x14 ^ 1'b0 ;
  assign n5300 = n5299 ^ n5289 ^ n5042 ;
  assign n5301 = ( n5042 & n5289 ) | ( n5042 & n5299 ) | ( n5289 & n5299 ) ;
  assign n5302 = x69 & n4972 ;
  assign n5303 = ( x71 & n4985 ) | ( x71 & n5302 ) | ( n4985 & n5302 ) ;
  assign n5304 = n5302 | n5303 ;
  assign n5305 = x70 & ~n4980 ;
  assign n5306 = ( x70 & n5304 ) | ( x70 & ~n5305 ) | ( n5304 & ~n5305 ) ;
  assign n5307 = n328 & n4987 ;
  assign n5308 = n5306 | n5307 ;
  assign n5309 = n5308 ^ x14 ^ 1'b0 ;
  assign n5310 = n5309 ^ n5301 ^ n5051 ;
  assign n5311 = ( n5051 & n5301 ) | ( n5051 & n5309 ) | ( n5301 & n5309 ) ;
  assign n5312 = n5311 ^ n5291 ^ n5062 ;
  assign n5313 = ( n5062 & n5291 ) | ( n5062 & n5311 ) | ( n5291 & n5311 ) ;
  assign n5314 = x71 & n4972 ;
  assign n5315 = ( x73 & n4985 ) | ( x73 & n5314 ) | ( n4985 & n5314 ) ;
  assign n5316 = n5314 | n5315 ;
  assign n5317 = x72 & ~n4980 ;
  assign n5318 = ( x72 & n5316 ) | ( x72 & ~n5317 ) | ( n5316 & ~n5317 ) ;
  assign n5319 = n370 & n4987 ;
  assign n5320 = n5318 | n5319 ;
  assign n5321 = n5320 ^ x14 ^ 1'b0 ;
  assign n5322 = ( n5071 & n5313 ) | ( n5071 & n5321 ) | ( n5313 & n5321 ) ;
  assign n5323 = n5321 ^ n5313 ^ n5071 ;
  assign n5324 = x72 & n4972 ;
  assign n5325 = ( x74 & n4985 ) | ( x74 & n5324 ) | ( n4985 & n5324 ) ;
  assign n5326 = n5324 | n5325 ;
  assign n5327 = x73 & ~n4980 ;
  assign n5328 = ( x73 & n5326 ) | ( x73 & ~n5327 ) | ( n5326 & ~n5327 ) ;
  assign n5329 = n504 & n4987 ;
  assign n5330 = n5328 | n5329 ;
  assign n5331 = n5330 ^ x14 ^ 1'b0 ;
  assign n5332 = ( n5081 & n5322 ) | ( n5081 & n5331 ) | ( n5322 & n5331 ) ;
  assign n5333 = n5331 ^ n5322 ^ n5081 ;
  assign n5334 = x73 & n4972 ;
  assign n5335 = ( x75 & n4985 ) | ( x75 & n5334 ) | ( n4985 & n5334 ) ;
  assign n5336 = n5334 | n5335 ;
  assign n5337 = x74 & ~n4980 ;
  assign n5338 = ( x74 & n5336 ) | ( x74 & ~n5337 ) | ( n5336 & ~n5337 ) ;
  assign n5339 = n525 & n4987 ;
  assign n5340 = n5338 | n5339 ;
  assign n5341 = n5340 ^ x14 ^ 1'b0 ;
  assign n5342 = n5341 ^ n5332 ^ n5092 ;
  assign n5343 = ( n5092 & n5332 ) | ( n5092 & n5341 ) | ( n5332 & n5341 ) ;
  assign n5344 = x74 & n4972 ;
  assign n5345 = ( x76 & n4985 ) | ( x76 & n5344 ) | ( n4985 & n5344 ) ;
  assign n5346 = n5344 | n5345 ;
  assign n5347 = x75 & ~n4980 ;
  assign n5348 = ( x75 & n5346 ) | ( x75 & ~n5347 ) | ( n5346 & ~n5347 ) ;
  assign n5349 = n664 & n4987 ;
  assign n5350 = n5348 | n5349 ;
  assign n5351 = n5350 ^ x14 ^ 1'b0 ;
  assign n5352 = ( n5101 & n5343 ) | ( n5101 & n5351 ) | ( n5343 & n5351 ) ;
  assign n5353 = n5351 ^ n5343 ^ n5101 ;
  assign n5354 = x75 & n4972 ;
  assign n5355 = ( x77 & n4985 ) | ( x77 & n5354 ) | ( n4985 & n5354 ) ;
  assign n5356 = n5354 | n5355 ;
  assign n5357 = x76 & ~n4980 ;
  assign n5358 = ( x76 & n5356 ) | ( x76 & ~n5357 ) | ( n5356 & ~n5357 ) ;
  assign n5359 = n690 & n4987 ;
  assign n5360 = n5358 | n5359 ;
  assign n5361 = n5360 ^ x14 ^ 1'b0 ;
  assign n5362 = n5361 ^ n5352 ^ n5112 ;
  assign n5363 = ( n5112 & n5352 ) | ( n5112 & n5361 ) | ( n5352 & n5361 ) ;
  assign n5364 = x76 & n4972 ;
  assign n5365 = ( x78 & n4985 ) | ( x78 & n5364 ) | ( n4985 & n5364 ) ;
  assign n5366 = n5364 | n5365 ;
  assign n5367 = x77 & ~n4980 ;
  assign n5368 = ( x77 & n5366 ) | ( x77 & ~n5367 ) | ( n5366 & ~n5367 ) ;
  assign n5369 = n709 & n4987 ;
  assign n5370 = n5368 | n5369 ;
  assign n5371 = n5370 ^ x14 ^ 1'b0 ;
  assign n5372 = n5371 ^ n5363 ^ n5122 ;
  assign n5373 = ( n5122 & n5363 ) | ( n5122 & n5371 ) | ( n5363 & n5371 ) ;
  assign n5374 = x77 & n4972 ;
  assign n5375 = ( x79 & n4985 ) | ( x79 & n5374 ) | ( n4985 & n5374 ) ;
  assign n5376 = n5374 | n5375 ;
  assign n5377 = x78 & ~n4980 ;
  assign n5378 = ( x78 & n5376 ) | ( x78 & ~n5377 ) | ( n5376 & ~n5377 ) ;
  assign n5379 = n1015 & n4987 ;
  assign n5380 = n5378 | n5379 ;
  assign n5381 = n5380 ^ x14 ^ 1'b0 ;
  assign n5382 = ( n5131 & n5373 ) | ( n5131 & n5381 ) | ( n5373 & n5381 ) ;
  assign n5383 = n5381 ^ n5373 ^ n5131 ;
  assign n5384 = x78 & n4972 ;
  assign n5385 = ( x80 & n4985 ) | ( x80 & n5384 ) | ( n4985 & n5384 ) ;
  assign n5386 = n5384 | n5385 ;
  assign n5387 = x79 & ~n4980 ;
  assign n5388 = ( x79 & n5386 ) | ( x79 & ~n5387 ) | ( n5386 & ~n5387 ) ;
  assign n5389 = n1216 & n4987 ;
  assign n5390 = n5388 | n5389 ;
  assign n5391 = n5390 ^ x14 ^ 1'b0 ;
  assign n5392 = ( n5142 & n5382 ) | ( n5142 & n5391 ) | ( n5382 & n5391 ) ;
  assign n5393 = n5391 ^ n5382 ^ n5142 ;
  assign n5394 = x79 & n4972 ;
  assign n5395 = ( x81 & n4985 ) | ( x81 & n5394 ) | ( n4985 & n5394 ) ;
  assign n5396 = n5394 | n5395 ;
  assign n5397 = x80 & ~n4980 ;
  assign n5398 = ( x80 & n5396 ) | ( x80 & ~n5397 ) | ( n5396 & ~n5397 ) ;
  assign n5399 = n1258 & n4987 ;
  assign n5400 = n5398 | n5399 ;
  assign n5401 = n5400 ^ x14 ^ 1'b0 ;
  assign n5402 = ( n5151 & n5392 ) | ( n5151 & n5401 ) | ( n5392 & n5401 ) ;
  assign n5403 = n5401 ^ n5392 ^ n5151 ;
  assign n5404 = x80 & n4972 ;
  assign n5405 = ( x82 & n4985 ) | ( x82 & n5404 ) | ( n4985 & n5404 ) ;
  assign n5406 = n5404 | n5405 ;
  assign n5407 = x81 & ~n4980 ;
  assign n5408 = ( x81 & n5406 ) | ( x81 & ~n5407 ) | ( n5406 & ~n5407 ) ;
  assign n5409 = n1301 & n4987 ;
  assign n5410 = n5408 | n5409 ;
  assign n5411 = n5410 ^ x14 ^ 1'b0 ;
  assign n5412 = n5411 ^ n5402 ^ n5162 ;
  assign n5413 = ( n5162 & n5402 ) | ( n5162 & n5411 ) | ( n5402 & n5411 ) ;
  assign n5414 = x81 & n4972 ;
  assign n5415 = ( x83 & n4985 ) | ( x83 & n5414 ) | ( n4985 & n5414 ) ;
  assign n5416 = n5414 | n5415 ;
  assign n5417 = x82 & ~n4980 ;
  assign n5418 = ( x82 & n5416 ) | ( x82 & ~n5417 ) | ( n5416 & ~n5417 ) ;
  assign n5419 = n1329 & n4987 ;
  assign n5420 = n5418 | n5419 ;
  assign n5421 = n5420 ^ x14 ^ 1'b0 ;
  assign n5422 = n5421 ^ n5413 ^ n5171 ;
  assign n5423 = ( n5171 & n5413 ) | ( n5171 & n5421 ) | ( n5413 & n5421 ) ;
  assign n5424 = x82 & n4972 ;
  assign n5425 = ( x84 & n4985 ) | ( x84 & n5424 ) | ( n4985 & n5424 ) ;
  assign n5426 = n5424 | n5425 ;
  assign n5427 = x83 & ~n4980 ;
  assign n5428 = ( x83 & n5426 ) | ( x83 & ~n5427 ) | ( n5426 & ~n5427 ) ;
  assign n5429 = n1355 & n4987 ;
  assign n5430 = n5428 | n5429 ;
  assign n5431 = n5430 ^ x14 ^ 1'b0 ;
  assign n5432 = n5431 ^ n5423 ^ n5182 ;
  assign n5433 = ( n5182 & n5423 ) | ( n5182 & n5431 ) | ( n5423 & n5431 ) ;
  assign n5434 = x83 & n4972 ;
  assign n5435 = ( x85 & n4985 ) | ( x85 & n5434 ) | ( n4985 & n5434 ) ;
  assign n5436 = n5434 | n5435 ;
  assign n5437 = x84 & ~n4980 ;
  assign n5438 = ( x84 & n5436 ) | ( x84 & ~n5437 ) | ( n5436 & ~n5437 ) ;
  assign n5439 = n1392 & n4987 ;
  assign n5440 = n5438 | n5439 ;
  assign n5441 = n5440 ^ x14 ^ 1'b0 ;
  assign n5442 = ( n5191 & n5433 ) | ( n5191 & n5441 ) | ( n5433 & n5441 ) ;
  assign n5443 = n5441 ^ n5433 ^ n5191 ;
  assign n5444 = x84 & n4972 ;
  assign n5445 = ( x86 & n4985 ) | ( x86 & n5444 ) | ( n4985 & n5444 ) ;
  assign n5446 = n5444 | n5445 ;
  assign n5447 = x85 & ~n4980 ;
  assign n5448 = ( x85 & n5446 ) | ( x85 & ~n5447 ) | ( n5446 & ~n5447 ) ;
  assign n5449 = n1419 & n4987 ;
  assign n5450 = n5448 | n5449 ;
  assign n5451 = n5450 ^ x14 ^ 1'b0 ;
  assign n5452 = ( n5201 & n5442 ) | ( n5201 & n5451 ) | ( n5442 & n5451 ) ;
  assign n5453 = n5451 ^ n5442 ^ n5201 ;
  assign n5454 = x85 & n4972 ;
  assign n5455 = ( x87 & n4985 ) | ( x87 & n5454 ) | ( n4985 & n5454 ) ;
  assign n5456 = n5454 | n5455 ;
  assign n5457 = x86 & ~n4980 ;
  assign n5458 = ( x86 & n5456 ) | ( x86 & ~n5457 ) | ( n5456 & ~n5457 ) ;
  assign n5459 = n1484 & n4987 ;
  assign n5460 = n5458 | n5459 ;
  assign n5461 = n5460 ^ x14 ^ 1'b0 ;
  assign n5462 = n5461 ^ n5452 ^ n5211 ;
  assign n5463 = ( n5211 & n5452 ) | ( n5211 & n5461 ) | ( n5452 & n5461 ) ;
  assign n5464 = x86 & n4972 ;
  assign n5465 = ( x88 & n4985 ) | ( x88 & n5464 ) | ( n4985 & n5464 ) ;
  assign n5466 = n5464 | n5465 ;
  assign n5467 = x87 & ~n4980 ;
  assign n5468 = ( x87 & n5466 ) | ( x87 & ~n5467 ) | ( n5466 & ~n5467 ) ;
  assign n5469 = n1569 & n4987 ;
  assign n5470 = n5468 | n5469 ;
  assign n5471 = n5470 ^ x14 ^ 1'b0 ;
  assign n5472 = ( n5222 & n5463 ) | ( n5222 & n5471 ) | ( n5463 & n5471 ) ;
  assign n5473 = n5471 ^ n5463 ^ n5222 ;
  assign n5474 = x87 & n4972 ;
  assign n5475 = ( x89 & n4985 ) | ( x89 & n5474 ) | ( n4985 & n5474 ) ;
  assign n5476 = n5474 | n5475 ;
  assign n5477 = x88 & ~n4980 ;
  assign n5478 = ( x88 & n5476 ) | ( x88 & ~n5477 ) | ( n5476 & ~n5477 ) ;
  assign n5479 = n1654 & n4987 ;
  assign n5480 = n5478 | n5479 ;
  assign n5481 = n5480 ^ x14 ^ 1'b0 ;
  assign n5482 = n5481 ^ n5472 ^ n5232 ;
  assign n5483 = ( n5232 & n5472 ) | ( n5232 & n5481 ) | ( n5472 & n5481 ) ;
  assign n5484 = x88 & n4972 ;
  assign n5485 = ( x90 & n4985 ) | ( x90 & n5484 ) | ( n4985 & n5484 ) ;
  assign n5486 = n5484 | n5485 ;
  assign n5487 = x89 & ~n4980 ;
  assign n5488 = ( x89 & n5486 ) | ( x89 & ~n5487 ) | ( n5486 & ~n5487 ) ;
  assign n5489 = n1741 & n4987 ;
  assign n5490 = n5488 | n5489 ;
  assign n5491 = n5490 ^ x14 ^ 1'b0 ;
  assign n5492 = n5491 ^ n5483 ^ n5241 ;
  assign n5493 = ( n5241 & n5483 ) | ( n5241 & n5491 ) | ( n5483 & n5491 ) ;
  assign n5494 = x9 ^ x8 ^ 1'b0 ;
  assign n5495 = x11 ^ x10 ^ 1'b0 ;
  assign n5496 = x10 ^ x9 ^ 1'b0 ;
  assign n5497 = n5494 & ~n5495 ;
  assign n5498 = ( ~n5494 & n5495 ) | ( ~n5494 & n5496 ) | ( n5495 & n5496 ) ;
  assign n5499 = ~n5496 & n5498 ;
  assign n5500 = x64 & n5499 ;
  assign n5501 = n5494 & n5495 ;
  assign n5502 = ~n5494 & n5496 ;
  assign n5503 = n139 & n5501 ;
  assign n5504 = x65 & ~n5502 ;
  assign n5505 = x64 & n5494 ;
  assign n5506 = ( x66 & n5497 ) | ( x66 & n5500 ) | ( n5497 & n5500 ) ;
  assign n5507 = n5500 | n5506 ;
  assign n5508 = ( x65 & ~n5504 ) | ( x65 & n5507 ) | ( ~n5504 & n5507 ) ;
  assign n5509 = n5503 | n5508 ;
  assign n5510 = x65 & n5499 ;
  assign n5511 = x64 & n5502 ;
  assign n5512 = ( x67 & n5497 ) | ( x67 & n5510 ) | ( n5497 & n5510 ) ;
  assign n5513 = n5510 | n5512 ;
  assign n5514 = ~x65 & n5497 ;
  assign n5515 = ( n5497 & n5511 ) | ( n5497 & ~n5514 ) | ( n5511 & ~n5514 ) ;
  assign n5516 = x11 & ~n5505 ;
  assign n5517 = ( n190 & n5501 ) | ( n190 & n5511 ) | ( n5501 & n5511 ) ;
  assign n5518 = n5515 | n5517 ;
  assign n5519 = n5518 ^ x11 ^ 1'b0 ;
  assign n5520 = n5519 ^ n5516 ^ 1'b0 ;
  assign n5521 = n5516 & n5519 ;
  assign n5522 = x66 & ~n5502 ;
  assign n5523 = ( x66 & n5513 ) | ( x66 & ~n5522 ) | ( n5513 & ~n5522 ) ;
  assign n5524 = n5509 ^ x11 ^ 1'b0 ;
  assign n5525 = n161 & n5501 ;
  assign n5526 = n5523 | n5525 ;
  assign n5527 = n5521 & n5524 ;
  assign n5528 = n5526 ^ x11 ^ 1'b0 ;
  assign n5529 = n5524 ^ n5521 ^ 1'b0 ;
  assign n5530 = n5528 ^ n5527 ^ n4995 ;
  assign n5531 = ( n4995 & n5527 ) | ( n4995 & n5528 ) | ( n5527 & n5528 ) ;
  assign n5532 = x66 & n5499 ;
  assign n5533 = ( x68 & n5497 ) | ( x68 & n5532 ) | ( n5497 & n5532 ) ;
  assign n5534 = n5532 | n5533 ;
  assign n5535 = x67 & ~n5502 ;
  assign n5536 = ( x67 & n5534 ) | ( x67 & ~n5535 ) | ( n5534 & ~n5535 ) ;
  assign n5537 = n175 & n5501 ;
  assign n5538 = n5536 | n5537 ;
  assign n5539 = n5538 ^ x11 ^ 1'b0 ;
  assign n5540 = n5539 ^ n5531 ^ n5260 ;
  assign n5541 = ( n5260 & n5531 ) | ( n5260 & n5539 ) | ( n5531 & n5539 ) ;
  assign n5542 = x67 & n5499 ;
  assign n5543 = ( x69 & n5497 ) | ( x69 & n5542 ) | ( n5497 & n5542 ) ;
  assign n5544 = n5542 | n5543 ;
  assign n5545 = x68 & ~n5502 ;
  assign n5546 = ( x68 & n5544 ) | ( x68 & ~n5545 ) | ( n5544 & ~n5545 ) ;
  assign n5547 = n172 & n5501 ;
  assign n5548 = n5546 | n5547 ;
  assign n5549 = n5548 ^ x11 ^ 1'b0 ;
  assign n5550 = ( n5262 & n5541 ) | ( n5262 & n5549 ) | ( n5541 & n5549 ) ;
  assign n5551 = n5549 ^ n5541 ^ n5262 ;
  assign n5552 = x68 & n5499 ;
  assign n5553 = ( x70 & n5497 ) | ( x70 & n5552 ) | ( n5497 & n5552 ) ;
  assign n5554 = n5552 | n5553 ;
  assign n5555 = x69 & ~n5502 ;
  assign n5556 = ( x69 & n5554 ) | ( x69 & ~n5555 ) | ( n5554 & ~n5555 ) ;
  assign n5557 = n168 & n5501 ;
  assign n5558 = n5556 | n5557 ;
  assign n5559 = n5558 ^ x11 ^ 1'b0 ;
  assign n5560 = n5559 ^ n5550 ^ n5271 ;
  assign n5561 = ( n5271 & n5550 ) | ( n5271 & n5559 ) | ( n5550 & n5559 ) ;
  assign n5562 = x69 & n5499 ;
  assign n5563 = ( x71 & n5497 ) | ( x71 & n5562 ) | ( n5497 & n5562 ) ;
  assign n5564 = n5562 | n5563 ;
  assign n5565 = x70 & ~n5502 ;
  assign n5566 = ( x70 & n5564 ) | ( x70 & ~n5565 ) | ( n5564 & ~n5565 ) ;
  assign n5567 = n328 & n5501 ;
  assign n5568 = n5566 | n5567 ;
  assign n5569 = n5568 ^ x11 ^ 1'b0 ;
  assign n5570 = ( n5281 & n5561 ) | ( n5281 & n5569 ) | ( n5561 & n5569 ) ;
  assign n5571 = n5569 ^ n5561 ^ n5281 ;
  assign n5572 = x70 & n5499 ;
  assign n5573 = ( x72 & n5497 ) | ( x72 & n5572 ) | ( n5497 & n5572 ) ;
  assign n5574 = n5572 | n5573 ;
  assign n5575 = x71 & ~n5502 ;
  assign n5576 = ( x71 & n5574 ) | ( x71 & ~n5575 ) | ( n5574 & ~n5575 ) ;
  assign n5577 = n349 & n5501 ;
  assign n5578 = n5576 | n5577 ;
  assign n5579 = n5578 ^ x11 ^ 1'b0 ;
  assign n5580 = n5579 ^ n5570 ^ n5290 ;
  assign n5581 = ( n5290 & n5570 ) | ( n5290 & n5579 ) | ( n5570 & n5579 ) ;
  assign n5582 = x71 & n5499 ;
  assign n5583 = ( x73 & n5497 ) | ( x73 & n5582 ) | ( n5497 & n5582 ) ;
  assign n5584 = n5582 | n5583 ;
  assign n5585 = x72 & ~n5502 ;
  assign n5586 = ( x72 & n5584 ) | ( x72 & ~n5585 ) | ( n5584 & ~n5585 ) ;
  assign n5587 = n370 & n5501 ;
  assign n5588 = n5586 | n5587 ;
  assign n5589 = n5588 ^ x11 ^ 1'b0 ;
  assign n5590 = n5589 ^ n5581 ^ n5300 ;
  assign n5591 = ( n5300 & n5581 ) | ( n5300 & n5589 ) | ( n5581 & n5589 ) ;
  assign n5592 = x72 & n5499 ;
  assign n5593 = ( x74 & n5497 ) | ( x74 & n5592 ) | ( n5497 & n5592 ) ;
  assign n5594 = n5592 | n5593 ;
  assign n5595 = x73 & ~n5502 ;
  assign n5596 = ( x73 & n5594 ) | ( x73 & ~n5595 ) | ( n5594 & ~n5595 ) ;
  assign n5597 = n504 & n5501 ;
  assign n5598 = n5596 | n5597 ;
  assign n5599 = n5598 ^ x11 ^ 1'b0 ;
  assign n5600 = n5599 ^ n5591 ^ n5310 ;
  assign n5601 = ( n5310 & n5591 ) | ( n5310 & n5599 ) | ( n5591 & n5599 ) ;
  assign n5602 = x73 & n5499 ;
  assign n5603 = ( x75 & n5497 ) | ( x75 & n5602 ) | ( n5497 & n5602 ) ;
  assign n5604 = n5602 | n5603 ;
  assign n5605 = x74 & ~n5502 ;
  assign n5606 = ( x74 & n5604 ) | ( x74 & ~n5605 ) | ( n5604 & ~n5605 ) ;
  assign n5607 = n525 & n5501 ;
  assign n5608 = n5606 | n5607 ;
  assign n5609 = n5608 ^ x11 ^ 1'b0 ;
  assign n5610 = n5609 ^ n5601 ^ n5312 ;
  assign n5611 = ( n5312 & n5601 ) | ( n5312 & n5609 ) | ( n5601 & n5609 ) ;
  assign n5612 = x74 & n5499 ;
  assign n5613 = ( x76 & n5497 ) | ( x76 & n5612 ) | ( n5497 & n5612 ) ;
  assign n5614 = n5612 | n5613 ;
  assign n5615 = x75 & ~n5502 ;
  assign n5616 = ( x75 & n5614 ) | ( x75 & ~n5615 ) | ( n5614 & ~n5615 ) ;
  assign n5617 = n664 & n5501 ;
  assign n5618 = n5616 | n5617 ;
  assign n5619 = n5618 ^ x11 ^ 1'b0 ;
  assign n5620 = ( n5323 & n5611 ) | ( n5323 & n5619 ) | ( n5611 & n5619 ) ;
  assign n5621 = n5619 ^ n5611 ^ n5323 ;
  assign n5622 = x75 & n5499 ;
  assign n5623 = ( x77 & n5497 ) | ( x77 & n5622 ) | ( n5497 & n5622 ) ;
  assign n5624 = n5622 | n5623 ;
  assign n5625 = x76 & ~n5502 ;
  assign n5626 = ( x76 & n5624 ) | ( x76 & ~n5625 ) | ( n5624 & ~n5625 ) ;
  assign n5627 = n690 & n5501 ;
  assign n5628 = n5626 | n5627 ;
  assign n5629 = n5628 ^ x11 ^ 1'b0 ;
  assign n5630 = n5629 ^ n5620 ^ n5333 ;
  assign n5631 = ( n5333 & n5620 ) | ( n5333 & n5629 ) | ( n5620 & n5629 ) ;
  assign n5632 = x76 & n5499 ;
  assign n5633 = ( x78 & n5497 ) | ( x78 & n5632 ) | ( n5497 & n5632 ) ;
  assign n5634 = n5632 | n5633 ;
  assign n5635 = x77 & ~n5502 ;
  assign n5636 = ( x77 & n5634 ) | ( x77 & ~n5635 ) | ( n5634 & ~n5635 ) ;
  assign n5637 = n709 & n5501 ;
  assign n5638 = n5636 | n5637 ;
  assign n5639 = n5638 ^ x11 ^ 1'b0 ;
  assign n5640 = ( n5342 & n5631 ) | ( n5342 & n5639 ) | ( n5631 & n5639 ) ;
  assign n5641 = n5639 ^ n5631 ^ n5342 ;
  assign n5642 = x77 & n5499 ;
  assign n5643 = ( x79 & n5497 ) | ( x79 & n5642 ) | ( n5497 & n5642 ) ;
  assign n5644 = n5642 | n5643 ;
  assign n5645 = x78 & ~n5502 ;
  assign n5646 = ( x78 & n5644 ) | ( x78 & ~n5645 ) | ( n5644 & ~n5645 ) ;
  assign n5647 = n1015 & n5501 ;
  assign n5648 = n5646 | n5647 ;
  assign n5649 = n5648 ^ x11 ^ 1'b0 ;
  assign n5650 = ( n5353 & n5640 ) | ( n5353 & n5649 ) | ( n5640 & n5649 ) ;
  assign n5651 = n5649 ^ n5640 ^ n5353 ;
  assign n5652 = x78 & n5499 ;
  assign n5653 = ( x80 & n5497 ) | ( x80 & n5652 ) | ( n5497 & n5652 ) ;
  assign n5654 = n5652 | n5653 ;
  assign n5655 = x79 & ~n5502 ;
  assign n5656 = ( x79 & n5654 ) | ( x79 & ~n5655 ) | ( n5654 & ~n5655 ) ;
  assign n5657 = n1216 & n5501 ;
  assign n5658 = n5656 | n5657 ;
  assign n5659 = n5658 ^ x11 ^ 1'b0 ;
  assign n5660 = ( n5362 & n5650 ) | ( n5362 & n5659 ) | ( n5650 & n5659 ) ;
  assign n5661 = n5659 ^ n5650 ^ n5362 ;
  assign n5662 = x80 & ~n5502 ;
  assign n5663 = x79 & n5499 ;
  assign n5664 = ( x81 & n5497 ) | ( x81 & n5663 ) | ( n5497 & n5663 ) ;
  assign n5665 = n5663 | n5664 ;
  assign n5666 = ( x80 & ~n5662 ) | ( x80 & n5665 ) | ( ~n5662 & n5665 ) ;
  assign n5667 = n1258 & n5501 ;
  assign n5668 = n5666 | n5667 ;
  assign n5669 = x80 & n5499 ;
  assign n5670 = n5668 ^ x11 ^ 1'b0 ;
  assign n5671 = ( n5372 & n5660 ) | ( n5372 & n5670 ) | ( n5660 & n5670 ) ;
  assign n5672 = n5670 ^ n5660 ^ n5372 ;
  assign n5673 = x99 & n1058 ;
  assign n5674 = ( x82 & n5497 ) | ( x82 & n5669 ) | ( n5497 & n5669 ) ;
  assign n5675 = n5669 | n5674 ;
  assign n5676 = x81 & ~n5502 ;
  assign n5677 = ( x81 & n5675 ) | ( x81 & ~n5676 ) | ( n5675 & ~n5676 ) ;
  assign n5678 = ( x101 & n1065 ) | ( x101 & n5673 ) | ( n1065 & n5673 ) ;
  assign n5679 = n5673 | n5678 ;
  assign n5680 = n1301 & n5501 ;
  assign n5681 = n5677 | n5680 ;
  assign n5682 = x100 & ~n1060 ;
  assign n5683 = n5681 ^ x11 ^ 1'b0 ;
  assign n5684 = ( x100 & n5679 ) | ( x100 & ~n5682 ) | ( n5679 & ~n5682 ) ;
  assign n5685 = n5683 ^ n5671 ^ n5383 ;
  assign n5686 = ( n5383 & n5671 ) | ( n5383 & n5683 ) | ( n5671 & n5683 ) ;
  assign n5687 = n4443 ^ x101 ^ x100 ;
  assign n5688 = n1063 & n5687 ;
  assign n5689 = n5684 | n5688 ;
  assign n5690 = n5689 ^ x41 ^ 1'b0 ;
  assign n5691 = n5690 ^ n4056 ^ n3687 ;
  assign n5692 = ( n3687 & n4056 ) | ( n3687 & n5690 ) | ( n4056 & n5690 ) ;
  assign n5693 = x81 & n5499 ;
  assign n5694 = ( x83 & n5497 ) | ( x83 & n5693 ) | ( n5497 & n5693 ) ;
  assign n5695 = n5693 | n5694 ;
  assign n5696 = x82 & ~n5502 ;
  assign n5697 = ( x82 & n5695 ) | ( x82 & ~n5696 ) | ( n5695 & ~n5696 ) ;
  assign n5698 = n1329 & n5501 ;
  assign n5699 = n5697 | n5698 ;
  assign n5700 = n5699 ^ x11 ^ 1'b0 ;
  assign n5701 = n5700 ^ n5686 ^ n5393 ;
  assign n5702 = ( x100 & x101 ) | ( x100 & n4443 ) | ( x101 & n4443 ) ;
  assign n5703 = ( n5393 & n5686 ) | ( n5393 & n5700 ) | ( n5686 & n5700 ) ;
  assign n5704 = x99 & n888 ;
  assign n5705 = ( x101 & n878 ) | ( x101 & n5704 ) | ( n878 & n5704 ) ;
  assign n5706 = n5704 | n5705 ;
  assign n5707 = x100 & ~n877 ;
  assign n5708 = ( x100 & n5706 ) | ( x100 & ~n5707 ) | ( n5706 & ~n5707 ) ;
  assign n5709 = n880 & n5687 ;
  assign n5710 = n5708 | n5709 ;
  assign n5711 = n5710 ^ x44 ^ 1'b0 ;
  assign n5712 = ( n4266 & n4453 ) | ( n4266 & n5711 ) | ( n4453 & n5711 ) ;
  assign n5713 = n5711 ^ n4453 ^ n4266 ;
  assign n5714 = x6 ^ x5 ^ 1'b0 ;
  assign n5715 = x8 ^ x7 ^ 1'b0 ;
  assign n5716 = x7 ^ x6 ^ 1'b0 ;
  assign n5717 = ( ~n5714 & n5715 ) | ( ~n5714 & n5716 ) | ( n5715 & n5716 ) ;
  assign n5718 = ~n5716 & n5717 ;
  assign n5719 = x65 & n5718 ;
  assign n5720 = n5714 & ~n5715 ;
  assign n5721 = x64 & n5718 ;
  assign n5722 = ( x67 & n5719 ) | ( x67 & n5720 ) | ( n5719 & n5720 ) ;
  assign n5723 = ( x66 & n5720 ) | ( x66 & n5721 ) | ( n5720 & n5721 ) ;
  assign n5724 = n5721 | n5723 ;
  assign n5725 = n5719 | n5722 ;
  assign n5726 = n5714 & n5715 ;
  assign n5727 = ~n5714 & n5716 ;
  assign n5728 = x66 & ~n5727 ;
  assign n5729 = ( x66 & n5725 ) | ( x66 & ~n5728 ) | ( n5725 & ~n5728 ) ;
  assign n5730 = x65 & ~n5727 ;
  assign n5731 = ( x65 & n5724 ) | ( x65 & ~n5730 ) | ( n5724 & ~n5730 ) ;
  assign n5732 = n161 & n5726 ;
  assign n5733 = n139 & n5726 ;
  assign n5734 = n5731 | n5733 ;
  assign n5735 = n5729 | n5732 ;
  assign n5736 = x64 & n5727 ;
  assign n5737 = ( n190 & n5726 ) | ( n190 & n5736 ) | ( n5726 & n5736 ) ;
  assign n5738 = ~x65 & n5720 ;
  assign n5739 = ( n5720 & n5736 ) | ( n5720 & ~n5738 ) | ( n5736 & ~n5738 ) ;
  assign n5740 = n5737 | n5739 ;
  assign n5741 = n5740 ^ x8 ^ 1'b0 ;
  assign n5742 = x64 & n5714 ;
  assign n5743 = n5735 ^ x8 ^ 1'b0 ;
  assign n5744 = x8 & ~n5742 ;
  assign n5745 = n5741 & n5744 ;
  assign n5746 = n5734 ^ x8 ^ 1'b0 ;
  assign n5747 = n5744 ^ n5741 ^ 1'b0 ;
  assign n5748 = n5745 & n5746 ;
  assign n5749 = n5746 ^ n5745 ^ 1'b0 ;
  assign n5750 = n5748 ^ n5743 ^ n5505 ;
  assign n5751 = ( n5505 & n5743 ) | ( n5505 & n5748 ) | ( n5743 & n5748 ) ;
  assign n5752 = x66 & n5718 ;
  assign n5753 = ( x68 & n5720 ) | ( x68 & n5752 ) | ( n5720 & n5752 ) ;
  assign n5754 = n5752 | n5753 ;
  assign n5755 = x67 & ~n5727 ;
  assign n5756 = ( x67 & n5754 ) | ( x67 & ~n5755 ) | ( n5754 & ~n5755 ) ;
  assign n5757 = n175 & n5726 ;
  assign n5758 = n5756 | n5757 ;
  assign n5759 = n5758 ^ x8 ^ 1'b0 ;
  assign n5760 = ( n5520 & n5751 ) | ( n5520 & n5759 ) | ( n5751 & n5759 ) ;
  assign n5761 = n5759 ^ n5751 ^ n5520 ;
  assign n5762 = x67 & n5718 ;
  assign n5763 = ( x69 & n5720 ) | ( x69 & n5762 ) | ( n5720 & n5762 ) ;
  assign n5764 = n5762 | n5763 ;
  assign n5765 = x68 & ~n5727 ;
  assign n5766 = ( x68 & n5764 ) | ( x68 & ~n5765 ) | ( n5764 & ~n5765 ) ;
  assign n5767 = n172 & n5726 ;
  assign n5768 = n5766 | n5767 ;
  assign n5769 = n5768 ^ x8 ^ 1'b0 ;
  assign n5770 = ( n5529 & n5760 ) | ( n5529 & n5769 ) | ( n5760 & n5769 ) ;
  assign n5771 = n5769 ^ n5760 ^ n5529 ;
  assign n5772 = x68 & n5718 ;
  assign n5773 = ( x70 & n5720 ) | ( x70 & n5772 ) | ( n5720 & n5772 ) ;
  assign n5774 = n5772 | n5773 ;
  assign n5775 = x69 & ~n5727 ;
  assign n5776 = ( x69 & n5774 ) | ( x69 & ~n5775 ) | ( n5774 & ~n5775 ) ;
  assign n5777 = n168 & n5726 ;
  assign n5778 = n5776 | n5777 ;
  assign n5779 = n5778 ^ x8 ^ 1'b0 ;
  assign n5780 = ( n5530 & n5770 ) | ( n5530 & n5779 ) | ( n5770 & n5779 ) ;
  assign n5781 = n5779 ^ n5770 ^ n5530 ;
  assign n5782 = x69 & n5718 ;
  assign n5783 = ( x71 & n5720 ) | ( x71 & n5782 ) | ( n5720 & n5782 ) ;
  assign n5784 = n5782 | n5783 ;
  assign n5785 = x70 & ~n5727 ;
  assign n5786 = ( x70 & n5784 ) | ( x70 & ~n5785 ) | ( n5784 & ~n5785 ) ;
  assign n5787 = n328 & n5726 ;
  assign n5788 = n5786 | n5787 ;
  assign n5789 = n5788 ^ x8 ^ 1'b0 ;
  assign n5790 = n5789 ^ n5780 ^ n5540 ;
  assign n5791 = ( n5540 & n5780 ) | ( n5540 & n5789 ) | ( n5780 & n5789 ) ;
  assign n5792 = x70 & n5718 ;
  assign n5793 = ( x72 & n5720 ) | ( x72 & n5792 ) | ( n5720 & n5792 ) ;
  assign n5794 = n5792 | n5793 ;
  assign n5795 = x71 & ~n5727 ;
  assign n5796 = ( x71 & n5794 ) | ( x71 & ~n5795 ) | ( n5794 & ~n5795 ) ;
  assign n5797 = n349 & n5726 ;
  assign n5798 = n5796 | n5797 ;
  assign n5799 = n5798 ^ x8 ^ 1'b0 ;
  assign n5800 = n5799 ^ n5791 ^ n5551 ;
  assign n5801 = ( n5551 & n5791 ) | ( n5551 & n5799 ) | ( n5791 & n5799 ) ;
  assign n5802 = x71 & n5718 ;
  assign n5803 = ( x73 & n5720 ) | ( x73 & n5802 ) | ( n5720 & n5802 ) ;
  assign n5804 = n5802 | n5803 ;
  assign n5805 = x72 & ~n5727 ;
  assign n5806 = ( x72 & n5804 ) | ( x72 & ~n5805 ) | ( n5804 & ~n5805 ) ;
  assign n5807 = n370 & n5726 ;
  assign n5808 = n5806 | n5807 ;
  assign n5809 = n5808 ^ x8 ^ 1'b0 ;
  assign n5810 = n5809 ^ n5801 ^ n5560 ;
  assign n5811 = ( n5560 & n5801 ) | ( n5560 & n5809 ) | ( n5801 & n5809 ) ;
  assign n5812 = x72 & n5718 ;
  assign n5813 = ( x74 & n5720 ) | ( x74 & n5812 ) | ( n5720 & n5812 ) ;
  assign n5814 = n5812 | n5813 ;
  assign n5815 = x73 & ~n5727 ;
  assign n5816 = ( x73 & n5814 ) | ( x73 & ~n5815 ) | ( n5814 & ~n5815 ) ;
  assign n5817 = n504 & n5726 ;
  assign n5818 = n5816 | n5817 ;
  assign n5819 = n5818 ^ x8 ^ 1'b0 ;
  assign n5820 = n5819 ^ n5811 ^ n5571 ;
  assign n5821 = ( n5571 & n5811 ) | ( n5571 & n5819 ) | ( n5811 & n5819 ) ;
  assign n5822 = x73 & n5718 ;
  assign n5823 = ( x75 & n5720 ) | ( x75 & n5822 ) | ( n5720 & n5822 ) ;
  assign n5824 = n5822 | n5823 ;
  assign n5825 = x74 & ~n5727 ;
  assign n5826 = ( x74 & n5824 ) | ( x74 & ~n5825 ) | ( n5824 & ~n5825 ) ;
  assign n5827 = n525 & n5726 ;
  assign n5828 = n5826 | n5827 ;
  assign n5829 = n5828 ^ x8 ^ 1'b0 ;
  assign n5830 = n5829 ^ n5821 ^ n5580 ;
  assign n5831 = ( n5580 & n5821 ) | ( n5580 & n5829 ) | ( n5821 & n5829 ) ;
  assign n5832 = x74 & n5718 ;
  assign n5833 = ( x76 & n5720 ) | ( x76 & n5832 ) | ( n5720 & n5832 ) ;
  assign n5834 = n5832 | n5833 ;
  assign n5835 = x75 & ~n5727 ;
  assign n5836 = ( x75 & n5834 ) | ( x75 & ~n5835 ) | ( n5834 & ~n5835 ) ;
  assign n5837 = n664 & n5726 ;
  assign n5838 = n5836 | n5837 ;
  assign n5839 = n5838 ^ x8 ^ 1'b0 ;
  assign n5840 = n5839 ^ n5831 ^ n5590 ;
  assign n5841 = ( n5590 & n5831 ) | ( n5590 & n5839 ) | ( n5831 & n5839 ) ;
  assign n5842 = x75 & n5718 ;
  assign n5843 = ( x77 & n5720 ) | ( x77 & n5842 ) | ( n5720 & n5842 ) ;
  assign n5844 = n5842 | n5843 ;
  assign n5845 = x76 & ~n5727 ;
  assign n5846 = ( x76 & n5844 ) | ( x76 & ~n5845 ) | ( n5844 & ~n5845 ) ;
  assign n5847 = n690 & n5726 ;
  assign n5848 = n5846 | n5847 ;
  assign n5849 = n5848 ^ x8 ^ 1'b0 ;
  assign n5850 = n5849 ^ n5841 ^ n5600 ;
  assign n5851 = ( n5600 & n5841 ) | ( n5600 & n5849 ) | ( n5841 & n5849 ) ;
  assign n5852 = x76 & n5718 ;
  assign n5853 = ( x78 & n5720 ) | ( x78 & n5852 ) | ( n5720 & n5852 ) ;
  assign n5854 = n5852 | n5853 ;
  assign n5855 = x77 & ~n5727 ;
  assign n5856 = ( x77 & n5854 ) | ( x77 & ~n5855 ) | ( n5854 & ~n5855 ) ;
  assign n5857 = n709 & n5726 ;
  assign n5858 = n5856 | n5857 ;
  assign n5859 = n5858 ^ x8 ^ 1'b0 ;
  assign n5860 = n5859 ^ n5851 ^ n5610 ;
  assign n5861 = ( n5610 & n5851 ) | ( n5610 & n5859 ) | ( n5851 & n5859 ) ;
  assign n5862 = x77 & n5718 ;
  assign n5863 = ( x79 & n5720 ) | ( x79 & n5862 ) | ( n5720 & n5862 ) ;
  assign n5864 = n5862 | n5863 ;
  assign n5865 = x78 & ~n5727 ;
  assign n5866 = ( x78 & n5864 ) | ( x78 & ~n5865 ) | ( n5864 & ~n5865 ) ;
  assign n5867 = n1015 & n5726 ;
  assign n5868 = n5866 | n5867 ;
  assign n5869 = n5868 ^ x8 ^ 1'b0 ;
  assign n5870 = ( n5621 & n5861 ) | ( n5621 & n5869 ) | ( n5861 & n5869 ) ;
  assign n5871 = n5869 ^ n5861 ^ n5621 ;
  assign n5872 = x78 & n5718 ;
  assign n5873 = ( x80 & n5720 ) | ( x80 & n5872 ) | ( n5720 & n5872 ) ;
  assign n5874 = n5872 | n5873 ;
  assign n5875 = x79 & ~n5727 ;
  assign n5876 = ( x79 & n5874 ) | ( x79 & ~n5875 ) | ( n5874 & ~n5875 ) ;
  assign n5877 = n1216 & n5726 ;
  assign n5878 = n5876 | n5877 ;
  assign n5879 = n5878 ^ x8 ^ 1'b0 ;
  assign n5880 = ( n5630 & n5870 ) | ( n5630 & n5879 ) | ( n5870 & n5879 ) ;
  assign n5881 = n5879 ^ n5870 ^ n5630 ;
  assign n5882 = x79 & n5718 ;
  assign n5883 = ( x81 & n5720 ) | ( x81 & n5882 ) | ( n5720 & n5882 ) ;
  assign n5884 = n5882 | n5883 ;
  assign n5885 = x80 & ~n5727 ;
  assign n5886 = ( x80 & n5884 ) | ( x80 & ~n5885 ) | ( n5884 & ~n5885 ) ;
  assign n5887 = n1258 & n5726 ;
  assign n5888 = n5886 | n5887 ;
  assign n5889 = n5888 ^ x8 ^ 1'b0 ;
  assign n5890 = n5889 ^ n5880 ^ n5641 ;
  assign n5891 = ( n5641 & n5880 ) | ( n5641 & n5889 ) | ( n5880 & n5889 ) ;
  assign n5892 = x80 & n5718 ;
  assign n5893 = ( x82 & n5720 ) | ( x82 & n5892 ) | ( n5720 & n5892 ) ;
  assign n5894 = n5892 | n5893 ;
  assign n5895 = x81 & ~n5727 ;
  assign n5896 = ( x81 & n5894 ) | ( x81 & ~n5895 ) | ( n5894 & ~n5895 ) ;
  assign n5897 = n1301 & n5726 ;
  assign n5898 = n5896 | n5897 ;
  assign n5899 = n5898 ^ x8 ^ 1'b0 ;
  assign n5900 = ( n5651 & n5891 ) | ( n5651 & n5899 ) | ( n5891 & n5899 ) ;
  assign n5901 = n5899 ^ n5891 ^ n5651 ;
  assign n5902 = x81 & n5718 ;
  assign n5903 = x82 & n5718 ;
  assign n5904 = ( x84 & n5720 ) | ( x84 & n5903 ) | ( n5720 & n5903 ) ;
  assign n5905 = n5903 | n5904 ;
  assign n5906 = ( x83 & n5720 ) | ( x83 & n5902 ) | ( n5720 & n5902 ) ;
  assign n5907 = n5902 | n5906 ;
  assign n5908 = x82 & ~n5727 ;
  assign n5909 = ( x82 & n5907 ) | ( x82 & ~n5908 ) | ( n5907 & ~n5908 ) ;
  assign n5910 = n1329 & n5726 ;
  assign n5911 = n5909 | n5910 ;
  assign n5912 = n5911 ^ x8 ^ 1'b0 ;
  assign n5913 = n5912 ^ n5900 ^ n5661 ;
  assign n5914 = ( n5661 & n5900 ) | ( n5661 & n5912 ) | ( n5900 & n5912 ) ;
  assign n5915 = x83 & ~n5727 ;
  assign n5916 = ( x83 & n5905 ) | ( x83 & ~n5915 ) | ( n5905 & ~n5915 ) ;
  assign n5917 = n1355 & n5726 ;
  assign n5918 = n5916 | n5917 ;
  assign n5919 = n5918 ^ x8 ^ 1'b0 ;
  assign n5920 = ( n5672 & n5914 ) | ( n5672 & n5919 ) | ( n5914 & n5919 ) ;
  assign n5921 = n5919 ^ n5914 ^ n5672 ;
  assign n5922 = x83 & n5718 ;
  assign n5923 = ( x85 & n5720 ) | ( x85 & n5922 ) | ( n5720 & n5922 ) ;
  assign n5924 = n5922 | n5923 ;
  assign n5925 = x84 & ~n5727 ;
  assign n5926 = x84 & n5718 ;
  assign n5927 = ( x84 & n5924 ) | ( x84 & ~n5925 ) | ( n5924 & ~n5925 ) ;
  assign n5928 = n1392 & n5726 ;
  assign n5929 = n5927 | n5928 ;
  assign n5930 = ( x86 & n5720 ) | ( x86 & n5926 ) | ( n5720 & n5926 ) ;
  assign n5931 = n5926 | n5930 ;
  assign n5932 = x85 & ~n5727 ;
  assign n5933 = ( x85 & n5931 ) | ( x85 & ~n5932 ) | ( n5931 & ~n5932 ) ;
  assign n5934 = n5929 ^ x8 ^ 1'b0 ;
  assign n5935 = ( n5685 & n5920 ) | ( n5685 & n5934 ) | ( n5920 & n5934 ) ;
  assign n5936 = n5934 ^ n5920 ^ n5685 ;
  assign n5937 = x100 & n1058 ;
  assign n5938 = ( x102 & n1065 ) | ( x102 & n5937 ) | ( n1065 & n5937 ) ;
  assign n5939 = n5937 | n5938 ;
  assign n5940 = x101 & ~n1060 ;
  assign n5941 = ( x101 & n5939 ) | ( x101 & ~n5940 ) | ( n5939 & ~n5940 ) ;
  assign n5942 = n1419 & n5726 ;
  assign n5943 = n5933 | n5942 ;
  assign n5944 = n5943 ^ x8 ^ 1'b0 ;
  assign n5945 = ( n5701 & n5935 ) | ( n5701 & n5944 ) | ( n5935 & n5944 ) ;
  assign n5946 = n5944 ^ n5935 ^ n5701 ;
  assign n5947 = n5702 ^ x102 ^ x101 ;
  assign n5948 = n1063 & n5947 ;
  assign n5949 = n5941 | n5948 ;
  assign n5950 = n5949 ^ x41 ^ 1'b0 ;
  assign n5951 = ( n4057 & n4328 ) | ( n4057 & n5950 ) | ( n4328 & n5950 ) ;
  assign n5952 = ( x101 & x102 ) | ( x101 & n5702 ) | ( x102 & n5702 ) ;
  assign n5953 = n5950 ^ n4328 ^ n4057 ;
  assign n5954 = x100 & n888 ;
  assign n5955 = ( x102 & n878 ) | ( x102 & n5954 ) | ( n878 & n5954 ) ;
  assign n5956 = n5954 | n5955 ;
  assign n5957 = x101 & ~n877 ;
  assign n5958 = ( x101 & n5956 ) | ( x101 & ~n5957 ) | ( n5956 & ~n5957 ) ;
  assign n5959 = n880 & n5947 ;
  assign n5960 = n5958 | n5959 ;
  assign n5961 = n5960 ^ x44 ^ 1'b0 ;
  assign n5962 = ( n4452 & n4539 ) | ( n4452 & ~n5961 ) | ( n4539 & ~n5961 ) ;
  assign n5963 = n5961 ^ n4539 ^ n4452 ;
  assign n5964 = x3 ^ x2 ^ 1'b0 ;
  assign n5965 = x64 & n5964 ;
  assign n5966 = x4 ^ x3 ^ 1'b0 ;
  assign n5967 = x5 ^ x4 ^ 1'b0 ;
  assign n5968 = n5964 & n5967 ;
  assign n5969 = n5964 & ~n5967 ;
  assign n5970 = ~n5964 & n5966 ;
  assign n5971 = x64 & n5970 ;
  assign n5972 = ( n190 & n5968 ) | ( n190 & n5971 ) | ( n5968 & n5971 ) ;
  assign n5973 = ~x65 & n5969 ;
  assign n5974 = ( n5969 & n5971 ) | ( n5969 & ~n5973 ) | ( n5971 & ~n5973 ) ;
  assign n5975 = x65 & ~n5970 ;
  assign n5976 = n5972 | n5974 ;
  assign n5977 = n5976 ^ x5 ^ 1'b0 ;
  assign n5978 = ( ~n5964 & n5966 ) | ( ~n5964 & n5967 ) | ( n5966 & n5967 ) ;
  assign n5979 = ~n5966 & n5978 ;
  assign n5980 = x64 & n5979 ;
  assign n5981 = ( x66 & n5969 ) | ( x66 & n5980 ) | ( n5969 & n5980 ) ;
  assign n5982 = n5980 | n5981 ;
  assign n5983 = x5 & ~n5965 ;
  assign n5984 = n5977 & n5983 ;
  assign n5985 = ( x65 & ~n5975 ) | ( x65 & n5982 ) | ( ~n5975 & n5982 ) ;
  assign n5986 = ~n139 & n5968 ;
  assign n5987 = ( n5968 & n5985 ) | ( n5968 & ~n5986 ) | ( n5985 & ~n5986 ) ;
  assign n5988 = x65 & n5979 ;
  assign n5989 = n5987 ^ x5 ^ 1'b0 ;
  assign n5990 = n5983 ^ n5977 ^ 1'b0 ;
  assign n5991 = n5989 ^ n5984 ^ 1'b0 ;
  assign n5992 = n5984 & n5989 ;
  assign n5993 = ( x67 & n5969 ) | ( x67 & n5988 ) | ( n5969 & n5988 ) ;
  assign n5994 = n5988 | n5993 ;
  assign n5995 = x66 & ~n5970 ;
  assign n5996 = ( x66 & n5994 ) | ( x66 & ~n5995 ) | ( n5994 & ~n5995 ) ;
  assign n5997 = n161 & n5968 ;
  assign n5998 = n5996 | n5997 ;
  assign n5999 = n5998 ^ x5 ^ 1'b0 ;
  assign n6000 = n5999 ^ n5992 ^ n5742 ;
  assign n6001 = ( n5742 & n5992 ) | ( n5742 & n5999 ) | ( n5992 & n5999 ) ;
  assign n6002 = x66 & n5979 ;
  assign n6003 = ( x68 & n5969 ) | ( x68 & n6002 ) | ( n5969 & n6002 ) ;
  assign n6004 = n6002 | n6003 ;
  assign n6005 = x67 & ~n5970 ;
  assign n6006 = ( x67 & n6004 ) | ( x67 & ~n6005 ) | ( n6004 & ~n6005 ) ;
  assign n6007 = n175 & n5968 ;
  assign n6008 = n6006 | n6007 ;
  assign n6009 = n6008 ^ x5 ^ 1'b0 ;
  assign n6010 = n6009 ^ n6001 ^ n5747 ;
  assign n6011 = ( n5747 & n6001 ) | ( n5747 & n6009 ) | ( n6001 & n6009 ) ;
  assign n6012 = x67 & n5979 ;
  assign n6013 = ( x69 & n5969 ) | ( x69 & n6012 ) | ( n5969 & n6012 ) ;
  assign n6014 = n6012 | n6013 ;
  assign n6015 = x68 & ~n5970 ;
  assign n6016 = ( x68 & n6014 ) | ( x68 & ~n6015 ) | ( n6014 & ~n6015 ) ;
  assign n6017 = n172 & n5968 ;
  assign n6018 = n6016 | n6017 ;
  assign n6019 = n6018 ^ x5 ^ 1'b0 ;
  assign n6020 = ( n5749 & n6011 ) | ( n5749 & n6019 ) | ( n6011 & n6019 ) ;
  assign n6021 = n6019 ^ n6011 ^ n5749 ;
  assign n6022 = x68 & n5979 ;
  assign n6023 = ( x70 & n5969 ) | ( x70 & n6022 ) | ( n5969 & n6022 ) ;
  assign n6024 = n6022 | n6023 ;
  assign n6025 = x69 & ~n5970 ;
  assign n6026 = ( x69 & n6024 ) | ( x69 & ~n6025 ) | ( n6024 & ~n6025 ) ;
  assign n6027 = n168 & n5968 ;
  assign n6028 = n6026 | n6027 ;
  assign n6029 = n6028 ^ x5 ^ 1'b0 ;
  assign n6030 = n6029 ^ n6020 ^ n5750 ;
  assign n6031 = ( n5750 & n6020 ) | ( n5750 & n6029 ) | ( n6020 & n6029 ) ;
  assign n6032 = x69 & n5979 ;
  assign n6033 = ( x71 & n5969 ) | ( x71 & n6032 ) | ( n5969 & n6032 ) ;
  assign n6034 = n6032 | n6033 ;
  assign n6035 = x70 & ~n5970 ;
  assign n6036 = ( x70 & n6034 ) | ( x70 & ~n6035 ) | ( n6034 & ~n6035 ) ;
  assign n6037 = n328 & n5968 ;
  assign n6038 = n6036 | n6037 ;
  assign n6039 = n6038 ^ x5 ^ 1'b0 ;
  assign n6040 = ( n5761 & n6031 ) | ( n5761 & n6039 ) | ( n6031 & n6039 ) ;
  assign n6041 = n6039 ^ n6031 ^ n5761 ;
  assign n6042 = x70 & n5979 ;
  assign n6043 = ( x72 & n5969 ) | ( x72 & n6042 ) | ( n5969 & n6042 ) ;
  assign n6044 = n6042 | n6043 ;
  assign n6045 = x71 & ~n5970 ;
  assign n6046 = ( x71 & n6044 ) | ( x71 & ~n6045 ) | ( n6044 & ~n6045 ) ;
  assign n6047 = n349 & n5968 ;
  assign n6048 = n6046 | n6047 ;
  assign n6049 = n6048 ^ x5 ^ 1'b0 ;
  assign n6050 = ( n5771 & n6040 ) | ( n5771 & n6049 ) | ( n6040 & n6049 ) ;
  assign n6051 = n6049 ^ n6040 ^ n5771 ;
  assign n6052 = x71 & n5979 ;
  assign n6053 = ( x73 & n5969 ) | ( x73 & n6052 ) | ( n5969 & n6052 ) ;
  assign n6054 = n6052 | n6053 ;
  assign n6055 = x72 & ~n5970 ;
  assign n6056 = ( x72 & n6054 ) | ( x72 & ~n6055 ) | ( n6054 & ~n6055 ) ;
  assign n6057 = n370 & n5968 ;
  assign n6058 = n6056 | n6057 ;
  assign n6059 = n6058 ^ x5 ^ 1'b0 ;
  assign n6060 = ( n5781 & n6050 ) | ( n5781 & n6059 ) | ( n6050 & n6059 ) ;
  assign n6061 = n6059 ^ n6050 ^ n5781 ;
  assign n6062 = x72 & n5979 ;
  assign n6063 = ( x74 & n5969 ) | ( x74 & n6062 ) | ( n5969 & n6062 ) ;
  assign n6064 = n6062 | n6063 ;
  assign n6065 = x73 & ~n5970 ;
  assign n6066 = ( x73 & n6064 ) | ( x73 & ~n6065 ) | ( n6064 & ~n6065 ) ;
  assign n6067 = n504 & n5968 ;
  assign n6068 = n6066 | n6067 ;
  assign n6069 = n6068 ^ x5 ^ 1'b0 ;
  assign n6070 = n6069 ^ n6060 ^ n5790 ;
  assign n6071 = ( n5790 & n6060 ) | ( n5790 & n6069 ) | ( n6060 & n6069 ) ;
  assign n6072 = x73 & n5979 ;
  assign n6073 = ( x75 & n5969 ) | ( x75 & n6072 ) | ( n5969 & n6072 ) ;
  assign n6074 = n6072 | n6073 ;
  assign n6075 = x74 & ~n5970 ;
  assign n6076 = ( x74 & n6074 ) | ( x74 & ~n6075 ) | ( n6074 & ~n6075 ) ;
  assign n6077 = n525 & n5968 ;
  assign n6078 = n6076 | n6077 ;
  assign n6079 = n6078 ^ x5 ^ 1'b0 ;
  assign n6080 = ( n5800 & n6071 ) | ( n5800 & n6079 ) | ( n6071 & n6079 ) ;
  assign n6081 = n6079 ^ n6071 ^ n5800 ;
  assign n6082 = x74 & n5979 ;
  assign n6083 = ( x76 & n5969 ) | ( x76 & n6082 ) | ( n5969 & n6082 ) ;
  assign n6084 = n6082 | n6083 ;
  assign n6085 = x75 & ~n5970 ;
  assign n6086 = ( x75 & n6084 ) | ( x75 & ~n6085 ) | ( n6084 & ~n6085 ) ;
  assign n6087 = n664 & n5968 ;
  assign n6088 = n6086 | n6087 ;
  assign n6089 = n6088 ^ x5 ^ 1'b0 ;
  assign n6090 = ( n5810 & n6080 ) | ( n5810 & n6089 ) | ( n6080 & n6089 ) ;
  assign n6091 = n6089 ^ n6080 ^ n5810 ;
  assign n6092 = x75 & n5979 ;
  assign n6093 = ( x77 & n5969 ) | ( x77 & n6092 ) | ( n5969 & n6092 ) ;
  assign n6094 = n6092 | n6093 ;
  assign n6095 = x76 & ~n5970 ;
  assign n6096 = ( x76 & n6094 ) | ( x76 & ~n6095 ) | ( n6094 & ~n6095 ) ;
  assign n6097 = n690 & n5968 ;
  assign n6098 = n6096 | n6097 ;
  assign n6099 = n6098 ^ x5 ^ 1'b0 ;
  assign n6100 = ( n5820 & n6090 ) | ( n5820 & n6099 ) | ( n6090 & n6099 ) ;
  assign n6101 = n6099 ^ n6090 ^ n5820 ;
  assign n6102 = x2 ^ x1 ^ 1'b0 ;
  assign n6103 = ( ~x0 & x1 ) | ( ~x0 & x2 ) | ( x1 & x2 ) ;
  assign n6104 = ~x1 & n6103 ;
  assign n6105 = x0 & ~n6102 ;
  assign n6106 = x70 & n6104 ;
  assign n6107 = ~x0 & x1 ;
  assign n6108 = x0 & n6102 ;
  assign n6109 = ( x72 & n6105 ) | ( x72 & n6106 ) | ( n6105 & n6106 ) ;
  assign n6110 = n6106 | n6109 ;
  assign n6111 = x71 & ~n6107 ;
  assign n6112 = ( x71 & n6110 ) | ( x71 & ~n6111 ) | ( n6110 & ~n6111 ) ;
  assign n6113 = n349 & ~n6108 ;
  assign n6114 = ( n349 & n6112 ) | ( n349 & ~n6113 ) | ( n6112 & ~n6113 ) ;
  assign n6115 = x65 & n6104 ;
  assign n6116 = ( x67 & n6105 ) | ( x67 & n6115 ) | ( n6105 & n6115 ) ;
  assign n6117 = n6115 | n6116 ;
  assign n6118 = x66 & ~n6107 ;
  assign n6119 = ( x66 & n6117 ) | ( x66 & ~n6118 ) | ( n6117 & ~n6118 ) ;
  assign n6120 = n161 & ~n6108 ;
  assign n6121 = ( n161 & n6119 ) | ( n161 & ~n6120 ) | ( n6119 & ~n6120 ) ;
  assign n6122 = x68 & n6104 ;
  assign n6123 = ( x70 & n6105 ) | ( x70 & n6122 ) | ( n6105 & n6122 ) ;
  assign n6124 = n6122 | n6123 ;
  assign n6125 = x69 & ~n6107 ;
  assign n6126 = ( x69 & n6124 ) | ( x69 & ~n6125 ) | ( n6124 & ~n6125 ) ;
  assign n6127 = n168 & ~n6108 ;
  assign n6128 = ( n168 & n6126 ) | ( n168 & ~n6127 ) | ( n6126 & ~n6127 ) ;
  assign n6129 = x69 & n6104 ;
  assign n6130 = ( x71 & n6105 ) | ( x71 & n6129 ) | ( n6105 & n6129 ) ;
  assign n6131 = n6129 | n6130 ;
  assign n6132 = x70 & ~n6107 ;
  assign n6133 = ( x70 & n6131 ) | ( x70 & ~n6132 ) | ( n6131 & ~n6132 ) ;
  assign n6134 = n328 & ~n6108 ;
  assign n6135 = ( n328 & n6133 ) | ( n328 & ~n6134 ) | ( n6133 & ~n6134 ) ;
  assign n6136 = x67 & n6104 ;
  assign n6137 = ( x69 & n6105 ) | ( x69 & n6136 ) | ( n6105 & n6136 ) ;
  assign n6138 = n6136 | n6137 ;
  assign n6139 = x68 & ~n6107 ;
  assign n6140 = ( x68 & n6138 ) | ( x68 & ~n6139 ) | ( n6138 & ~n6139 ) ;
  assign n6141 = n172 & ~n6108 ;
  assign n6142 = ( n172 & n6140 ) | ( n172 & ~n6141 ) | ( n6140 & ~n6141 ) ;
  assign n6143 = ~x65 & n6105 ;
  assign n6144 = x64 & n6104 ;
  assign n6145 = n139 & ~n6108 ;
  assign n6146 = ( n139 & n6144 ) | ( n139 & ~n6145 ) | ( n6144 & ~n6145 ) ;
  assign n6147 = x66 & n6105 ;
  assign n6148 = x65 & n6107 ;
  assign n6149 = ( ~n6144 & n6147 ) | ( ~n6144 & n6148 ) | ( n6147 & n6148 ) ;
  assign n6150 = x67 & ~n6107 ;
  assign n6151 = x64 & n6107 ;
  assign n6152 = ( n6105 & ~n6143 ) | ( n6105 & n6151 ) | ( ~n6143 & n6151 ) ;
  assign n6153 = n6121 ^ x2 ^ 1'b0 ;
  assign n6154 = ( n190 & n6108 ) | ( n190 & n6151 ) | ( n6108 & n6151 ) ;
  assign n6155 = x66 & n6104 ;
  assign n6156 = n6152 | n6154 ;
  assign n6157 = ( x68 & n6105 ) | ( x68 & n6155 ) | ( n6105 & n6155 ) ;
  assign n6158 = n6135 ^ x2 ^ 1'b0 ;
  assign n6159 = n6156 ^ x2 ^ 1'b0 ;
  assign n6160 = n6155 | n6157 ;
  assign n6161 = ( x67 & ~n6150 ) | ( x67 & n6160 ) | ( ~n6150 & n6160 ) ;
  assign n6162 = n175 & ~n6108 ;
  assign n6163 = n6128 ^ x2 ^ 1'b0 ;
  assign n6164 = n6146 | n6149 ;
  assign n6165 = n6164 ^ x2 ^ 1'b0 ;
  assign n6166 = n6114 ^ x2 ^ 1'b0 ;
  assign n6167 = n6142 ^ x2 ^ 1'b0 ;
  assign n6168 = ( n175 & n6161 ) | ( n175 & ~n6162 ) | ( n6161 & ~n6162 ) ;
  assign n6169 = n6168 ^ x2 ^ 1'b0 ;
  assign n6170 = x0 & x64 ;
  assign n6171 = x2 & ~n6170 ;
  assign n6172 = n6171 ^ n6159 ^ 1'b0 ;
  assign n6173 = n6159 & n6171 ;
  assign n6174 = n6165 & n6173 ;
  assign n6175 = n6174 ^ n6153 ^ n5965 ;
  assign n6176 = ( n5965 & n6153 ) | ( n5965 & n6174 ) | ( n6153 & n6174 ) ;
  assign n6177 = ( n5990 & n6169 ) | ( n5990 & n6176 ) | ( n6169 & n6176 ) ;
  assign n6178 = n6177 ^ n6167 ^ n5991 ;
  assign n6179 = n6176 ^ n6169 ^ n5990 ;
  assign n6180 = ( n5991 & n6167 ) | ( n5991 & n6177 ) | ( n6167 & n6177 ) ;
  assign n6181 = ( n6000 & n6163 ) | ( n6000 & n6180 ) | ( n6163 & n6180 ) ;
  assign n6182 = n6181 ^ n6158 ^ n6010 ;
  assign n6183 = n6180 ^ n6163 ^ n6000 ;
  assign n6184 = ( n6010 & n6158 ) | ( n6010 & n6181 ) | ( n6158 & n6181 ) ;
  assign n6185 = ( n6021 & n6166 ) | ( n6021 & n6184 ) | ( n6166 & n6184 ) ;
  assign n6186 = n6184 ^ n6166 ^ n6021 ;
  assign n6187 = x73 & n6104 ;
  assign n6188 = n6173 ^ n6165 ^ 1'b0 ;
  assign n6189 = ( x75 & n6105 ) | ( x75 & n6187 ) | ( n6105 & n6187 ) ;
  assign n6190 = n6187 | n6189 ;
  assign n6191 = x74 & ~n6107 ;
  assign n6192 = ( x74 & n6190 ) | ( x74 & ~n6191 ) | ( n6190 & ~n6191 ) ;
  assign n6193 = n525 & ~n6108 ;
  assign n6194 = ( n525 & n6192 ) | ( n525 & ~n6193 ) | ( n6192 & ~n6193 ) ;
  assign n6195 = x71 & n6104 ;
  assign n6196 = ( x73 & n6105 ) | ( x73 & n6195 ) | ( n6105 & n6195 ) ;
  assign n6197 = n6195 | n6196 ;
  assign n6198 = x72 & ~n6107 ;
  assign n6199 = ( x72 & n6197 ) | ( x72 & ~n6198 ) | ( n6197 & ~n6198 ) ;
  assign n6200 = n370 & ~n6108 ;
  assign n6201 = ( n370 & n6199 ) | ( n370 & ~n6200 ) | ( n6199 & ~n6200 ) ;
  assign n6202 = x75 & n6104 ;
  assign n6203 = ( x77 & n6105 ) | ( x77 & n6202 ) | ( n6105 & n6202 ) ;
  assign n6204 = n6202 | n6203 ;
  assign n6205 = x76 & ~n6107 ;
  assign n6206 = ( x76 & n6204 ) | ( x76 & ~n6205 ) | ( n6204 & ~n6205 ) ;
  assign n6207 = n690 & ~n6108 ;
  assign n6208 = ( n690 & n6206 ) | ( n690 & ~n6207 ) | ( n6206 & ~n6207 ) ;
  assign n6209 = x72 & n6104 ;
  assign n6210 = ( x74 & n6105 ) | ( x74 & n6209 ) | ( n6105 & n6209 ) ;
  assign n6211 = n6209 | n6210 ;
  assign n6212 = x73 & ~n6107 ;
  assign n6213 = ( x73 & n6211 ) | ( x73 & ~n6212 ) | ( n6211 & ~n6212 ) ;
  assign n6214 = n504 & ~n6108 ;
  assign n6215 = ( n504 & n6213 ) | ( n504 & ~n6214 ) | ( n6213 & ~n6214 ) ;
  assign n6216 = n6215 ^ x2 ^ 1'b0 ;
  assign n6217 = x76 & n6104 ;
  assign n6218 = n6201 ^ x2 ^ 1'b0 ;
  assign n6219 = ( n6030 & n6185 ) | ( n6030 & n6218 ) | ( n6185 & n6218 ) ;
  assign n6220 = n6218 ^ n6185 ^ n6030 ;
  assign n6221 = x74 & n6104 ;
  assign n6222 = ( n6041 & n6216 ) | ( n6041 & n6219 ) | ( n6216 & n6219 ) ;
  assign n6223 = n6219 ^ n6216 ^ n6041 ;
  assign n6224 = n664 & ~n6108 ;
  assign n6225 = ( x76 & n6105 ) | ( x76 & n6221 ) | ( n6105 & n6221 ) ;
  assign n6226 = n6221 | n6225 ;
  assign n6227 = x75 & ~n6107 ;
  assign n6228 = ( x75 & n6226 ) | ( x75 & ~n6227 ) | ( n6226 & ~n6227 ) ;
  assign n6229 = ( n664 & ~n6224 ) | ( n664 & n6228 ) | ( ~n6224 & n6228 ) ;
  assign n6230 = n6194 ^ x2 ^ 1'b0 ;
  assign n6231 = ( n6051 & n6222 ) | ( n6051 & n6230 ) | ( n6222 & n6230 ) ;
  assign n6232 = n6229 ^ x2 ^ 1'b0 ;
  assign n6233 = n6208 ^ x2 ^ 1'b0 ;
  assign n6234 = n6230 ^ n6222 ^ n6051 ;
  assign n6235 = x76 & n5979 ;
  assign n6236 = ( x78 & n5969 ) | ( x78 & n6235 ) | ( n5969 & n6235 ) ;
  assign n6237 = ( n6061 & n6231 ) | ( n6061 & n6232 ) | ( n6231 & n6232 ) ;
  assign n6238 = n6237 ^ n6233 ^ n6070 ;
  assign n6239 = ( n6070 & n6233 ) | ( n6070 & n6237 ) | ( n6233 & n6237 ) ;
  assign n6240 = n709 & n5968 ;
  assign n6241 = n6235 | n6236 ;
  assign n6242 = x77 & ~n6107 ;
  assign n6243 = ( x78 & n6105 ) | ( x78 & n6217 ) | ( n6105 & n6217 ) ;
  assign n6244 = n6217 | n6243 ;
  assign n6245 = n709 & ~n6108 ;
  assign n6246 = ( x77 & ~n6242 ) | ( x77 & n6244 ) | ( ~n6242 & n6244 ) ;
  assign n6247 = ( n709 & ~n6245 ) | ( n709 & n6246 ) | ( ~n6245 & n6246 ) ;
  assign n6248 = n6247 ^ x2 ^ 1'b0 ;
  assign n6249 = x77 & ~n5970 ;
  assign n6250 = ( x77 & n6241 ) | ( x77 & ~n6249 ) | ( n6241 & ~n6249 ) ;
  assign n6251 = n6240 | n6250 ;
  assign n6252 = n6248 ^ n6239 ^ n6081 ;
  assign n6253 = ( n6081 & n6239 ) | ( n6081 & n6248 ) | ( n6239 & n6248 ) ;
  assign n6254 = n6232 ^ n6231 ^ n6061 ;
  assign n6255 = n6251 ^ x5 ^ 1'b0 ;
  assign n6256 = ( n5830 & n6100 ) | ( n5830 & n6255 ) | ( n6100 & n6255 ) ;
  assign n6257 = n6255 ^ n6100 ^ n5830 ;
  assign n6258 = x77 & n6104 ;
  assign n6259 = ( x79 & n6105 ) | ( x79 & n6258 ) | ( n6105 & n6258 ) ;
  assign n6260 = n6258 | n6259 ;
  assign n6261 = x78 & ~n6107 ;
  assign n6262 = ( x78 & n6260 ) | ( x78 & ~n6261 ) | ( n6260 & ~n6261 ) ;
  assign n6263 = n1015 & ~n6108 ;
  assign n6264 = ( n1015 & n6262 ) | ( n1015 & ~n6263 ) | ( n6262 & ~n6263 ) ;
  assign n6265 = n6264 ^ x2 ^ 1'b0 ;
  assign n6266 = n6265 ^ n6253 ^ n6091 ;
  assign n6267 = ( n6091 & n6253 ) | ( n6091 & n6265 ) | ( n6253 & n6265 ) ;
  assign n6268 = x77 & n5979 ;
  assign n6269 = ( x79 & n5969 ) | ( x79 & n6268 ) | ( n5969 & n6268 ) ;
  assign n6270 = n6268 | n6269 ;
  assign n6271 = x78 & ~n5970 ;
  assign n6272 = ( x78 & n6270 ) | ( x78 & ~n6271 ) | ( n6270 & ~n6271 ) ;
  assign n6273 = x78 & n6104 ;
  assign n6274 = n1015 & n5968 ;
  assign n6275 = n6272 | n6274 ;
  assign n6276 = n6275 ^ x5 ^ 1'b0 ;
  assign n6277 = ( x80 & n6105 ) | ( x80 & n6273 ) | ( n6105 & n6273 ) ;
  assign n6278 = n6273 | n6277 ;
  assign n6279 = n6276 ^ n6256 ^ n5840 ;
  assign n6280 = ( n5840 & n6256 ) | ( n5840 & n6276 ) | ( n6256 & n6276 ) ;
  assign n6281 = x78 & n5979 ;
  assign n6282 = x79 & ~n6107 ;
  assign n6283 = ( x79 & n6278 ) | ( x79 & ~n6282 ) | ( n6278 & ~n6282 ) ;
  assign n6284 = n1216 & ~n6108 ;
  assign n6285 = ( n1216 & n6283 ) | ( n1216 & ~n6284 ) | ( n6283 & ~n6284 ) ;
  assign n6286 = ( x80 & n5969 ) | ( x80 & n6281 ) | ( n5969 & n6281 ) ;
  assign n6287 = n6281 | n6286 ;
  assign n6288 = n6285 ^ x2 ^ 1'b0 ;
  assign n6289 = ( n6101 & n6267 ) | ( n6101 & n6288 ) | ( n6267 & n6288 ) ;
  assign n6290 = n6288 ^ n6267 ^ n6101 ;
  assign n6291 = x79 & ~n5970 ;
  assign n6292 = ( x79 & n6287 ) | ( x79 & ~n6291 ) | ( n6287 & ~n6291 ) ;
  assign n6293 = n1216 & n5968 ;
  assign n6294 = x80 & n5979 ;
  assign n6295 = x81 & ~n5970 ;
  assign n6296 = n6292 | n6293 ;
  assign n6297 = ( x82 & n5969 ) | ( x82 & n6294 ) | ( n5969 & n6294 ) ;
  assign n6298 = n6294 | n6297 ;
  assign n6299 = ( x81 & ~n6295 ) | ( x81 & n6298 ) | ( ~n6295 & n6298 ) ;
  assign n6300 = n1301 & n5968 ;
  assign n6301 = n6299 | n6300 ;
  assign n6302 = x79 & n5979 ;
  assign n6303 = ( x81 & n5969 ) | ( x81 & n6302 ) | ( n5969 & n6302 ) ;
  assign n6304 = n6302 | n6303 ;
  assign n6305 = n6301 ^ x5 ^ 1'b0 ;
  assign n6306 = x80 & ~n5970 ;
  assign n6307 = ( x80 & n6304 ) | ( x80 & ~n6306 ) | ( n6304 & ~n6306 ) ;
  assign n6308 = n1258 & n5968 ;
  assign n6309 = n6296 ^ x5 ^ 1'b0 ;
  assign n6310 = n6307 | n6308 ;
  assign n6311 = n6309 ^ n6280 ^ n5850 ;
  assign n6312 = ( n5850 & n6280 ) | ( n5850 & n6309 ) | ( n6280 & n6309 ) ;
  assign n6313 = n6310 ^ x5 ^ 1'b0 ;
  assign n6314 = n6313 ^ n6312 ^ n5860 ;
  assign n6315 = ( n5860 & n6312 ) | ( n5860 & n6313 ) | ( n6312 & n6313 ) ;
  assign n6316 = n6315 ^ n6305 ^ n5871 ;
  assign n6317 = ( n5871 & n6305 ) | ( n5871 & n6315 ) | ( n6305 & n6315 ) ;
  assign n6318 = x79 & n6104 ;
  assign n6319 = ( x81 & n6105 ) | ( x81 & n6318 ) | ( n6105 & n6318 ) ;
  assign n6320 = n6318 | n6319 ;
  assign n6321 = n1258 & ~n6108 ;
  assign n6322 = x80 & ~n6107 ;
  assign n6323 = ( x80 & n6320 ) | ( x80 & ~n6322 ) | ( n6320 & ~n6322 ) ;
  assign n6324 = ( n1258 & ~n6321 ) | ( n1258 & n6323 ) | ( ~n6321 & n6323 ) ;
  assign n6325 = n6324 ^ x2 ^ 1'b0 ;
  assign n6326 = n6325 ^ n6289 ^ n6257 ;
  assign n6327 = ( n6257 & n6289 ) | ( n6257 & n6325 ) | ( n6289 & n6325 ) ;
  assign n6328 = x81 & n5979 ;
  assign n6329 = ( x83 & n5969 ) | ( x83 & n6328 ) | ( n5969 & n6328 ) ;
  assign n6330 = n6328 | n6329 ;
  assign n6331 = x82 & ~n5970 ;
  assign n6332 = ( x82 & n6330 ) | ( x82 & ~n6331 ) | ( n6330 & ~n6331 ) ;
  assign n6333 = n1329 & n5968 ;
  assign n6334 = n6332 | n6333 ;
  assign n6335 = n6334 ^ x5 ^ 1'b0 ;
  assign n6336 = n6335 ^ n6317 ^ n5881 ;
  assign n6337 = ( n5881 & n6317 ) | ( n5881 & n6335 ) | ( n6317 & n6335 ) ;
  assign n6338 = x82 & n5979 ;
  assign n6339 = ( x84 & n5969 ) | ( x84 & n6338 ) | ( n5969 & n6338 ) ;
  assign n6340 = n6338 | n6339 ;
  assign n6341 = x83 & ~n5970 ;
  assign n6342 = ( x83 & n6340 ) | ( x83 & ~n6341 ) | ( n6340 & ~n6341 ) ;
  assign n6343 = n1355 & n5968 ;
  assign n6344 = n6342 | n6343 ;
  assign n6345 = n6344 ^ x5 ^ 1'b0 ;
  assign n6346 = n6345 ^ n6337 ^ n5890 ;
  assign n6347 = ( n5890 & n6337 ) | ( n5890 & n6345 ) | ( n6337 & n6345 ) ;
  assign n6348 = x83 & n5979 ;
  assign n6349 = ( x85 & n5969 ) | ( x85 & n6348 ) | ( n5969 & n6348 ) ;
  assign n6350 = n6348 | n6349 ;
  assign n6351 = x84 & ~n5970 ;
  assign n6352 = ( x84 & n6350 ) | ( x84 & ~n6351 ) | ( n6350 & ~n6351 ) ;
  assign n6353 = n1392 & n5968 ;
  assign n6354 = n6352 | n6353 ;
  assign n6355 = n6354 ^ x5 ^ 1'b0 ;
  assign n6356 = n6355 ^ n6347 ^ n5901 ;
  assign n6357 = ( n5901 & n6347 ) | ( n5901 & n6355 ) | ( n6347 & n6355 ) ;
  assign n6358 = x84 & n5979 ;
  assign n6359 = ( x86 & n5969 ) | ( x86 & n6358 ) | ( n5969 & n6358 ) ;
  assign n6360 = n6358 | n6359 ;
  assign n6361 = x85 & ~n5970 ;
  assign n6362 = ( x85 & n6360 ) | ( x85 & ~n6361 ) | ( n6360 & ~n6361 ) ;
  assign n6363 = n1419 & n5968 ;
  assign n6364 = n6362 | n6363 ;
  assign n6365 = n6364 ^ x5 ^ 1'b0 ;
  assign n6366 = n6365 ^ n6357 ^ n5913 ;
  assign n6367 = ( n5913 & n6357 ) | ( n5913 & n6365 ) | ( n6357 & n6365 ) ;
  assign n6368 = x85 & n5979 ;
  assign n6369 = ( x87 & n5969 ) | ( x87 & n6368 ) | ( n5969 & n6368 ) ;
  assign n6370 = n6368 | n6369 ;
  assign n6371 = x86 & ~n5970 ;
  assign n6372 = ( x86 & n6370 ) | ( x86 & ~n6371 ) | ( n6370 & ~n6371 ) ;
  assign n6373 = n1484 & n5968 ;
  assign n6374 = n6372 | n6373 ;
  assign n6375 = n6374 ^ x5 ^ 1'b0 ;
  assign n6376 = ( n5921 & n6367 ) | ( n5921 & n6375 ) | ( n6367 & n6375 ) ;
  assign n6377 = n6375 ^ n6367 ^ n5921 ;
  assign n6378 = x86 & n5979 ;
  assign n6379 = ( x88 & n5969 ) | ( x88 & n6378 ) | ( n5969 & n6378 ) ;
  assign n6380 = n6378 | n6379 ;
  assign n6381 = x87 & ~n5970 ;
  assign n6382 = ( x87 & n6380 ) | ( x87 & ~n6381 ) | ( n6380 & ~n6381 ) ;
  assign n6383 = n1569 & n5968 ;
  assign n6384 = n6382 | n6383 ;
  assign n6385 = n6384 ^ x5 ^ 1'b0 ;
  assign n6386 = n6385 ^ n6376 ^ n5936 ;
  assign n6387 = ( n5936 & n6376 ) | ( n5936 & n6385 ) | ( n6376 & n6385 ) ;
  assign n6388 = x80 & n6104 ;
  assign n6389 = ( x82 & n6105 ) | ( x82 & n6388 ) | ( n6105 & n6388 ) ;
  assign n6390 = n6388 | n6389 ;
  assign n6391 = x81 & ~n6107 ;
  assign n6392 = ( x81 & n6390 ) | ( x81 & ~n6391 ) | ( n6390 & ~n6391 ) ;
  assign n6393 = n1301 & ~n6108 ;
  assign n6394 = ( n1301 & n6392 ) | ( n1301 & ~n6393 ) | ( n6392 & ~n6393 ) ;
  assign n6395 = n6394 ^ x2 ^ 1'b0 ;
  assign n6396 = n1301 & n4608 ;
  assign n6397 = ( n6279 & n6327 ) | ( n6279 & n6395 ) | ( n6327 & n6395 ) ;
  assign n6398 = n6395 ^ n6327 ^ n6279 ;
  assign n6399 = x81 & n6104 ;
  assign n6400 = ( x83 & n6105 ) | ( x83 & n6399 ) | ( n6105 & n6399 ) ;
  assign n6401 = n6399 | n6400 ;
  assign n6402 = x82 & ~n6107 ;
  assign n6403 = ( x82 & n6401 ) | ( x82 & ~n6402 ) | ( n6401 & ~n6402 ) ;
  assign n6404 = n1329 & ~n6108 ;
  assign n6405 = ( n1329 & n6403 ) | ( n1329 & ~n6404 ) | ( n6403 & ~n6404 ) ;
  assign n6406 = n6405 ^ x2 ^ 1'b0 ;
  assign n6407 = n6406 ^ n6397 ^ n6311 ;
  assign n6408 = ( n6311 & n6397 ) | ( n6311 & n6406 ) | ( n6397 & n6406 ) ;
  assign n6409 = x82 & n6104 ;
  assign n6410 = ( x84 & n6105 ) | ( x84 & n6409 ) | ( n6105 & n6409 ) ;
  assign n6411 = n6409 | n6410 ;
  assign n6412 = x83 & ~n6107 ;
  assign n6413 = ( x83 & n6411 ) | ( x83 & ~n6412 ) | ( n6411 & ~n6412 ) ;
  assign n6414 = n1355 & ~n6108 ;
  assign n6415 = ( n1355 & n6413 ) | ( n1355 & ~n6414 ) | ( n6413 & ~n6414 ) ;
  assign n6416 = n6415 ^ x2 ^ 1'b0 ;
  assign n6417 = n6416 ^ n6408 ^ n6314 ;
  assign n6418 = ( n6314 & n6408 ) | ( n6314 & n6416 ) | ( n6408 & n6416 ) ;
  assign n6419 = x83 & n6104 ;
  assign n6420 = ( x85 & n6105 ) | ( x85 & n6419 ) | ( n6105 & n6419 ) ;
  assign n6421 = n6419 | n6420 ;
  assign n6422 = x84 & ~n6107 ;
  assign n6423 = ( x84 & n6421 ) | ( x84 & ~n6422 ) | ( n6421 & ~n6422 ) ;
  assign n6424 = n1392 & ~n6108 ;
  assign n6425 = ( n1392 & n6423 ) | ( n1392 & ~n6424 ) | ( n6423 & ~n6424 ) ;
  assign n6426 = n6425 ^ x2 ^ 1'b0 ;
  assign n6427 = ( n6316 & n6418 ) | ( n6316 & n6426 ) | ( n6418 & n6426 ) ;
  assign n6428 = n6426 ^ n6418 ^ n6316 ;
  assign n6429 = x84 & n6104 ;
  assign n6430 = ( x86 & n6105 ) | ( x86 & n6429 ) | ( n6105 & n6429 ) ;
  assign n6431 = n6429 | n6430 ;
  assign n6432 = x85 & ~n6107 ;
  assign n6433 = ( x85 & n6431 ) | ( x85 & ~n6432 ) | ( n6431 & ~n6432 ) ;
  assign n6434 = n1419 & ~n6108 ;
  assign n6435 = ( n1419 & n6433 ) | ( n1419 & ~n6434 ) | ( n6433 & ~n6434 ) ;
  assign n6436 = n6435 ^ x2 ^ 1'b0 ;
  assign n6437 = n6436 ^ n6427 ^ n6336 ;
  assign n6438 = ( n6336 & n6427 ) | ( n6336 & n6436 ) | ( n6427 & n6436 ) ;
  assign n6439 = x85 & n6104 ;
  assign n6440 = ( x87 & n6105 ) | ( x87 & n6439 ) | ( n6105 & n6439 ) ;
  assign n6441 = n6439 | n6440 ;
  assign n6442 = x86 & ~n6107 ;
  assign n6443 = ( x86 & n6441 ) | ( x86 & ~n6442 ) | ( n6441 & ~n6442 ) ;
  assign n6444 = n1484 & ~n6108 ;
  assign n6445 = ( n1484 & n6443 ) | ( n1484 & ~n6444 ) | ( n6443 & ~n6444 ) ;
  assign n6446 = n6445 ^ x2 ^ 1'b0 ;
  assign n6447 = ( n6346 & n6438 ) | ( n6346 & n6446 ) | ( n6438 & n6446 ) ;
  assign n6448 = n6446 ^ n6438 ^ n6346 ;
  assign n6449 = x86 & n6104 ;
  assign n6450 = ( x88 & n6105 ) | ( x88 & n6449 ) | ( n6105 & n6449 ) ;
  assign n6451 = n6449 | n6450 ;
  assign n6452 = x87 & ~n6107 ;
  assign n6453 = ( x87 & n6451 ) | ( x87 & ~n6452 ) | ( n6451 & ~n6452 ) ;
  assign n6454 = n1569 & ~n6108 ;
  assign n6455 = ( n1569 & n6453 ) | ( n1569 & ~n6454 ) | ( n6453 & ~n6454 ) ;
  assign n6456 = n6455 ^ x2 ^ 1'b0 ;
  assign n6457 = n6456 ^ n6447 ^ n6356 ;
  assign n6458 = ( n6356 & n6447 ) | ( n6356 & n6456 ) | ( n6447 & n6456 ) ;
  assign n6459 = x87 & n6104 ;
  assign n6460 = ( x89 & n6105 ) | ( x89 & n6459 ) | ( n6105 & n6459 ) ;
  assign n6461 = n6459 | n6460 ;
  assign n6462 = x88 & ~n6107 ;
  assign n6463 = ( x88 & n6461 ) | ( x88 & ~n6462 ) | ( n6461 & ~n6462 ) ;
  assign n6464 = n1654 & ~n6108 ;
  assign n6465 = ( n1654 & n6463 ) | ( n1654 & ~n6464 ) | ( n6463 & ~n6464 ) ;
  assign n6466 = n6465 ^ x2 ^ 1'b0 ;
  assign n6467 = ( n6366 & n6458 ) | ( n6366 & n6466 ) | ( n6458 & n6466 ) ;
  assign n6468 = n6466 ^ n6458 ^ n6366 ;
  assign n6469 = x88 & n6104 ;
  assign n6470 = ( x90 & n6105 ) | ( x90 & n6469 ) | ( n6105 & n6469 ) ;
  assign n6471 = n6469 | n6470 ;
  assign n6472 = x89 & ~n6107 ;
  assign n6473 = ( x89 & n6471 ) | ( x89 & ~n6472 ) | ( n6471 & ~n6472 ) ;
  assign n6474 = n1741 & ~n6108 ;
  assign n6475 = ( n1741 & n6473 ) | ( n1741 & ~n6474 ) | ( n6473 & ~n6474 ) ;
  assign n6476 = n6475 ^ x2 ^ 1'b0 ;
  assign n6477 = n6476 ^ n6467 ^ n6377 ;
  assign n6478 = ( n6377 & n6467 ) | ( n6377 & n6476 ) | ( n6467 & n6476 ) ;
  assign n6479 = x89 & n6104 ;
  assign n6480 = ( x91 & n6105 ) | ( x91 & n6479 ) | ( n6105 & n6479 ) ;
  assign n6481 = n6479 | n6480 ;
  assign n6482 = x90 & ~n6107 ;
  assign n6483 = ( x90 & n6481 ) | ( x90 & ~n6482 ) | ( n6481 & ~n6482 ) ;
  assign n6484 = n2114 & ~n6108 ;
  assign n6485 = ( n2114 & n6483 ) | ( n2114 & ~n6484 ) | ( n6483 & ~n6484 ) ;
  assign n6486 = n6485 ^ x2 ^ 1'b0 ;
  assign n6487 = ( n6386 & n6478 ) | ( n6386 & n6486 ) | ( n6478 & n6486 ) ;
  assign n6488 = n6486 ^ n6478 ^ n6386 ;
  assign n6489 = x87 & n5979 ;
  assign n6490 = ( x89 & n5969 ) | ( x89 & n6489 ) | ( n5969 & n6489 ) ;
  assign n6491 = n6489 | n6490 ;
  assign n6492 = x88 & ~n5970 ;
  assign n6493 = ( x88 & n6491 ) | ( x88 & ~n6492 ) | ( n6491 & ~n6492 ) ;
  assign n6494 = n1654 & n5968 ;
  assign n6495 = n6493 | n6494 ;
  assign n6496 = n6495 ^ x5 ^ 1'b0 ;
  assign n6497 = n6496 ^ n6387 ^ n5946 ;
  assign n6498 = ( n5946 & n6387 ) | ( n5946 & n6496 ) | ( n6387 & n6496 ) ;
  assign n6499 = x90 & n6104 ;
  assign n6500 = ( x92 & n6105 ) | ( x92 & n6499 ) | ( n6105 & n6499 ) ;
  assign n6501 = n6499 | n6500 ;
  assign n6502 = x91 & ~n6107 ;
  assign n6503 = ( x91 & n6501 ) | ( x91 & ~n6502 ) | ( n6501 & ~n6502 ) ;
  assign n6504 = n2420 & ~n6108 ;
  assign n6505 = ( n2420 & n6503 ) | ( n2420 & ~n6504 ) | ( n6503 & ~n6504 ) ;
  assign n6506 = n6505 ^ x2 ^ 1'b0 ;
  assign n6507 = n6506 ^ n6497 ^ n6487 ;
  assign n6508 = ( n6487 & n6497 ) | ( n6487 & n6506 ) | ( n6497 & n6506 ) ;
  assign n6509 = x80 & n4616 ;
  assign n6510 = ( x82 & n4606 ) | ( x82 & n6509 ) | ( n4606 & n6509 ) ;
  assign n6511 = n6509 | n6510 ;
  assign n6512 = x81 & ~n4605 ;
  assign n6513 = ( x81 & n6511 ) | ( x81 & ~n6512 ) | ( n6511 & ~n6512 ) ;
  assign n6514 = n6396 | n6513 ;
  assign n6515 = n6514 ^ x23 ^ 1'b0 ;
  assign n6516 = x83 & n5499 ;
  assign n6517 = ( x85 & n5497 ) | ( x85 & n6516 ) | ( n5497 & n6516 ) ;
  assign n6518 = n6516 | n6517 ;
  assign n6519 = ( n3885 & n4778 ) | ( n3885 & n6515 ) | ( n4778 & n6515 ) ;
  assign n6520 = x84 & ~n5502 ;
  assign n6521 = ( x84 & n6518 ) | ( x84 & ~n6520 ) | ( n6518 & ~n6520 ) ;
  assign n6522 = n1355 & n5501 ;
  assign n6523 = n1355 & n4608 ;
  assign n6524 = n6515 ^ n4778 ^ n3885 ;
  assign n6525 = x82 & n5499 ;
  assign n6526 = ( x84 & n5497 ) | ( x84 & n6525 ) | ( n5497 & n6525 ) ;
  assign n6527 = n6525 | n6526 ;
  assign n6528 = x83 & ~n5502 ;
  assign n6529 = ( x83 & n6527 ) | ( x83 & ~n6528 ) | ( n6527 & ~n6528 ) ;
  assign n6530 = x83 & n4790 ;
  assign n6531 = n6522 | n6529 ;
  assign n6532 = n6531 ^ x11 ^ 1'b0 ;
  assign n6533 = n6532 ^ n5703 ^ n5403 ;
  assign n6534 = ( n5403 & n5703 ) | ( n5403 & n6532 ) | ( n5703 & n6532 ) ;
  assign n6535 = ( x85 & n4792 ) | ( x85 & n6530 ) | ( n4792 & n6530 ) ;
  assign n6536 = x84 & ~n4786 ;
  assign n6537 = n6530 | n6535 ;
  assign n6538 = n1392 & n4787 ;
  assign n6539 = ( x84 & ~n6536 ) | ( x84 & n6537 ) | ( ~n6536 & n6537 ) ;
  assign n6540 = n6538 | n6539 ;
  assign n6541 = x83 & n4616 ;
  assign n6542 = ( x85 & n4606 ) | ( x85 & n6541 ) | ( n4606 & n6541 ) ;
  assign n6543 = n6541 | n6542 ;
  assign n6544 = n1392 & n5501 ;
  assign n6545 = n6521 | n6544 ;
  assign n6546 = n1392 & n4608 ;
  assign n6547 = n6545 ^ x11 ^ 1'b0 ;
  assign n6548 = x84 & ~n4605 ;
  assign n6549 = ( x84 & n6543 ) | ( x84 & ~n6548 ) | ( n6543 & ~n6548 ) ;
  assign n6550 = n6546 | n6549 ;
  assign n6551 = x81 & n4616 ;
  assign n6552 = ( x83 & n4606 ) | ( x83 & n6551 ) | ( n4606 & n6551 ) ;
  assign n6553 = n6551 | n6552 ;
  assign n6554 = n6547 ^ n6534 ^ n5412 ;
  assign n6555 = n1329 & n4608 ;
  assign n6556 = ( n5412 & n6534 ) | ( n5412 & n6547 ) | ( n6534 & n6547 ) ;
  assign n6557 = x82 & n4616 ;
  assign n6558 = x82 & ~n4605 ;
  assign n6559 = ( x82 & n6553 ) | ( x82 & ~n6558 ) | ( n6553 & ~n6558 ) ;
  assign n6560 = x83 & ~n4605 ;
  assign n6561 = n6550 ^ x23 ^ 1'b0 ;
  assign n6562 = n6555 | n6559 ;
  assign n6563 = n6540 ^ x20 ^ 1'b0 ;
  assign n6564 = ( x84 & n4606 ) | ( x84 & n6557 ) | ( n4606 & n6557 ) ;
  assign n6565 = n6557 | n6564 ;
  assign n6566 = ( x83 & ~n6560 ) | ( x83 & n6565 ) | ( ~n6560 & n6565 ) ;
  assign n6567 = n6523 | n6566 ;
  assign n6568 = ( n4996 & n6524 ) | ( n4996 & n6563 ) | ( n6524 & n6563 ) ;
  assign n6569 = n6563 ^ n6524 ^ n4996 ;
  assign n6570 = x84 & n4790 ;
  assign n6571 = n6567 ^ x23 ^ 1'b0 ;
  assign n6572 = ( x86 & n4792 ) | ( x86 & n6570 ) | ( n4792 & n6570 ) ;
  assign n6573 = x85 & ~n4786 ;
  assign n6574 = n6562 ^ x23 ^ 1'b0 ;
  assign n6575 = ( n3896 & n6519 ) | ( n3896 & n6574 ) | ( n6519 & n6574 ) ;
  assign n6576 = n6570 | n6572 ;
  assign n6577 = n6575 ^ n6571 ^ n3906 ;
  assign n6578 = ( n3906 & n6571 ) | ( n3906 & n6575 ) | ( n6571 & n6575 ) ;
  assign n6579 = ( n3915 & n6561 ) | ( n3915 & n6578 ) | ( n6561 & n6578 ) ;
  assign n6580 = ( x85 & ~n6573 ) | ( x85 & n6576 ) | ( ~n6573 & n6576 ) ;
  assign n6581 = n1419 & n4787 ;
  assign n6582 = n6580 | n6581 ;
  assign n6583 = n6582 ^ x20 ^ 1'b0 ;
  assign n6584 = n6574 ^ n6519 ^ n3896 ;
  assign n6585 = n6584 ^ n6583 ^ n6568 ;
  assign n6586 = ( n6568 & n6583 ) | ( n6568 & n6584 ) | ( n6583 & n6584 ) ;
  assign n6587 = n6578 ^ n6561 ^ n3915 ;
  assign n6588 = x84 & n4616 ;
  assign n6589 = ( x86 & n4606 ) | ( x86 & n6588 ) | ( n4606 & n6588 ) ;
  assign n6590 = n6588 | n6589 ;
  assign n6591 = x85 & ~n4605 ;
  assign n6592 = ( x85 & n6590 ) | ( x85 & ~n6591 ) | ( n6590 & ~n6591 ) ;
  assign n6593 = n1419 & n4608 ;
  assign n6594 = n6592 | n6593 ;
  assign n6595 = n6594 ^ x23 ^ 1'b0 ;
  assign n6596 = n6595 ^ n6579 ^ n3926 ;
  assign n6597 = ( n3926 & n6579 ) | ( n3926 & n6595 ) | ( n6579 & n6595 ) ;
  assign n6598 = x85 & n4616 ;
  assign n6599 = ( x87 & n4606 ) | ( x87 & n6598 ) | ( n4606 & n6598 ) ;
  assign n6600 = n6598 | n6599 ;
  assign n6601 = x86 & ~n4605 ;
  assign n6602 = ( x86 & n6600 ) | ( x86 & ~n6601 ) | ( n6600 & ~n6601 ) ;
  assign n6603 = n1484 & n4608 ;
  assign n6604 = n6602 | n6603 ;
  assign n6605 = n6604 ^ x23 ^ 1'b0 ;
  assign n6606 = n6605 ^ n6597 ^ n3936 ;
  assign n6607 = ( n3936 & n6597 ) | ( n3936 & n6605 ) | ( n6597 & n6605 ) ;
  assign n6608 = x86 & n5011 ;
  assign n6609 = ( x88 & n5012 ) | ( x88 & n6608 ) | ( n5012 & n6608 ) ;
  assign n6610 = n6608 | n6609 ;
  assign n6611 = x87 & ~n5008 ;
  assign n6612 = ( x87 & n6610 ) | ( x87 & ~n6611 ) | ( n6610 & ~n6611 ) ;
  assign n6613 = n1569 & n5020 ;
  assign n6614 = n6612 | n6613 ;
  assign n6615 = n6614 ^ x17 ^ 1'b0 ;
  assign n6616 = n6615 ^ n6569 ^ n5242 ;
  assign n6617 = ( n5242 & n6569 ) | ( n5242 & n6615 ) | ( n6569 & n6615 ) ;
  assign n6618 = x87 & n5011 ;
  assign n6619 = ( x89 & n5012 ) | ( x89 & n6618 ) | ( n5012 & n6618 ) ;
  assign n6620 = n6618 | n6619 ;
  assign n6621 = x88 & ~n5008 ;
  assign n6622 = ( x88 & n6620 ) | ( x88 & ~n6621 ) | ( n6620 & ~n6621 ) ;
  assign n6623 = n1654 & n5020 ;
  assign n6624 = n6622 | n6623 ;
  assign n6625 = n6624 ^ x17 ^ 1'b0 ;
  assign n6626 = ( n6585 & n6617 ) | ( n6585 & n6625 ) | ( n6617 & n6625 ) ;
  assign n6627 = n6625 ^ n6617 ^ n6585 ;
  assign n6628 = x86 & n4616 ;
  assign n6629 = ( x88 & n4606 ) | ( x88 & n6628 ) | ( n4606 & n6628 ) ;
  assign n6630 = n6628 | n6629 ;
  assign n6631 = x87 & ~n4605 ;
  assign n6632 = ( x87 & n6630 ) | ( x87 & ~n6631 ) | ( n6630 & ~n6631 ) ;
  assign n6633 = n1569 & n4608 ;
  assign n6634 = n6632 | n6633 ;
  assign n6635 = n6634 ^ x23 ^ 1'b0 ;
  assign n6636 = ( n3946 & n6607 ) | ( n3946 & n6635 ) | ( n6607 & n6635 ) ;
  assign n6637 = n6635 ^ n6607 ^ n3946 ;
  assign n6638 = x87 & n4616 ;
  assign n6639 = ( x89 & n4606 ) | ( x89 & n6638 ) | ( n4606 & n6638 ) ;
  assign n6640 = n6638 | n6639 ;
  assign n6641 = x88 & ~n4605 ;
  assign n6642 = ( x88 & n6640 ) | ( x88 & ~n6641 ) | ( n6640 & ~n6641 ) ;
  assign n6643 = n1654 & n4608 ;
  assign n6644 = n6642 | n6643 ;
  assign n6645 = n6644 ^ x23 ^ 1'b0 ;
  assign n6646 = ( n3955 & n6636 ) | ( n3955 & n6645 ) | ( n6636 & n6645 ) ;
  assign n6647 = n6645 ^ n6636 ^ n3955 ;
  assign n6648 = x85 & n4790 ;
  assign n6649 = ( x87 & n4792 ) | ( x87 & n6648 ) | ( n4792 & n6648 ) ;
  assign n6650 = n6648 | n6649 ;
  assign n6651 = x86 & ~n4786 ;
  assign n6652 = ( x86 & n6650 ) | ( x86 & ~n6651 ) | ( n6650 & ~n6651 ) ;
  assign n6653 = n1484 & n4787 ;
  assign n6654 = n6652 | n6653 ;
  assign n6655 = n6654 ^ x20 ^ 1'b0 ;
  assign n6656 = ( n6577 & n6586 ) | ( n6577 & n6655 ) | ( n6586 & n6655 ) ;
  assign n6657 = n6655 ^ n6586 ^ n6577 ;
  assign n6658 = x86 & n4790 ;
  assign n6659 = ( x88 & n4792 ) | ( x88 & n6658 ) | ( n4792 & n6658 ) ;
  assign n6660 = n6658 | n6659 ;
  assign n6661 = x87 & ~n4786 ;
  assign n6662 = ( x87 & n6660 ) | ( x87 & ~n6661 ) | ( n6660 & ~n6661 ) ;
  assign n6663 = n1569 & n4787 ;
  assign n6664 = n6662 | n6663 ;
  assign n6665 = n6664 ^ x20 ^ 1'b0 ;
  assign n6666 = n6665 ^ n6656 ^ n6587 ;
  assign n6667 = ( n6587 & n6656 ) | ( n6587 & n6665 ) | ( n6656 & n6665 ) ;
  assign n6668 = x88 & n5011 ;
  assign n6669 = ( x90 & n5012 ) | ( x90 & n6668 ) | ( n5012 & n6668 ) ;
  assign n6670 = n6668 | n6669 ;
  assign n6671 = x89 & ~n5008 ;
  assign n6672 = ( x89 & n6670 ) | ( x89 & ~n6671 ) | ( n6670 & ~n6671 ) ;
  assign n6673 = n1741 & n5020 ;
  assign n6674 = n6672 | n6673 ;
  assign n6675 = n6674 ^ x17 ^ 1'b0 ;
  assign n6676 = n6675 ^ n6657 ^ n6626 ;
  assign n6677 = ( n6626 & n6657 ) | ( n6626 & n6675 ) | ( n6657 & n6675 ) ;
  assign n6678 = x87 & n4790 ;
  assign n6679 = ( x89 & n4792 ) | ( x89 & n6678 ) | ( n4792 & n6678 ) ;
  assign n6680 = n6678 | n6679 ;
  assign n6681 = x88 & ~n4786 ;
  assign n6682 = ( x88 & n6680 ) | ( x88 & ~n6681 ) | ( n6680 & ~n6681 ) ;
  assign n6683 = n1654 & n4787 ;
  assign n6684 = n6682 | n6683 ;
  assign n6685 = n6684 ^ x20 ^ 1'b0 ;
  assign n6686 = ( n6596 & n6667 ) | ( n6596 & n6685 ) | ( n6667 & n6685 ) ;
  assign n6687 = n6685 ^ n6667 ^ n6596 ;
  assign n6688 = x84 & n5499 ;
  assign n6689 = ( x86 & n5497 ) | ( x86 & n6688 ) | ( n5497 & n6688 ) ;
  assign n6690 = n6688 | n6689 ;
  assign n6691 = x85 & ~n5502 ;
  assign n6692 = ( x85 & n6690 ) | ( x85 & ~n6691 ) | ( n6690 & ~n6691 ) ;
  assign n6693 = n1419 & n5501 ;
  assign n6694 = n6692 | n6693 ;
  assign n6695 = n6694 ^ x11 ^ 1'b0 ;
  assign n6696 = n6695 ^ n6556 ^ n5422 ;
  assign n6697 = ( n5422 & n6556 ) | ( n5422 & n6695 ) | ( n6556 & n6695 ) ;
  assign n6698 = x88 & n4790 ;
  assign n6699 = ( x90 & n4792 ) | ( x90 & n6698 ) | ( n4792 & n6698 ) ;
  assign n6700 = n6698 | n6699 ;
  assign n6701 = x89 & ~n4786 ;
  assign n6702 = ( x89 & n6700 ) | ( x89 & ~n6701 ) | ( n6700 & ~n6701 ) ;
  assign n6703 = n1741 & n4787 ;
  assign n6704 = n6702 | n6703 ;
  assign n6705 = n6704 ^ x20 ^ 1'b0 ;
  assign n6706 = ( n6606 & n6686 ) | ( n6606 & n6705 ) | ( n6686 & n6705 ) ;
  assign n6707 = n6705 ^ n6686 ^ n6606 ;
  assign n6708 = x89 & n5011 ;
  assign n6709 = ( x91 & n5012 ) | ( x91 & n6708 ) | ( n5012 & n6708 ) ;
  assign n6710 = n6708 | n6709 ;
  assign n6711 = x90 & ~n5008 ;
  assign n6712 = ( x90 & n6710 ) | ( x90 & ~n6711 ) | ( n6710 & ~n6711 ) ;
  assign n6713 = n2114 & n5020 ;
  assign n6714 = n6712 | n6713 ;
  assign n6715 = n6714 ^ x17 ^ 1'b0 ;
  assign n6716 = n6715 ^ n6677 ^ n6666 ;
  assign n6717 = ( n6666 & n6677 ) | ( n6666 & n6715 ) | ( n6677 & n6715 ) ;
  assign n6718 = x90 & n5011 ;
  assign n6719 = ( x92 & n5012 ) | ( x92 & n6718 ) | ( n5012 & n6718 ) ;
  assign n6720 = n6718 | n6719 ;
  assign n6721 = x91 & ~n5008 ;
  assign n6722 = ( x91 & n6720 ) | ( x91 & ~n6721 ) | ( n6720 & ~n6721 ) ;
  assign n6723 = n2420 & n5020 ;
  assign n6724 = n6722 | n6723 ;
  assign n6725 = n6724 ^ x17 ^ 1'b0 ;
  assign n6726 = n6725 ^ n6717 ^ n6687 ;
  assign n6727 = ( n6687 & n6717 ) | ( n6687 & n6725 ) | ( n6717 & n6725 ) ;
  assign n6728 = x89 & n4790 ;
  assign n6729 = ( x91 & n4792 ) | ( x91 & n6728 ) | ( n4792 & n6728 ) ;
  assign n6730 = n6728 | n6729 ;
  assign n6731 = x90 & ~n4786 ;
  assign n6732 = ( x90 & n6730 ) | ( x90 & ~n6731 ) | ( n6730 & ~n6731 ) ;
  assign n6733 = n2114 & n4787 ;
  assign n6734 = n6732 | n6733 ;
  assign n6735 = n6734 ^ x20 ^ 1'b0 ;
  assign n6736 = ( n6637 & n6706 ) | ( n6637 & n6735 ) | ( n6706 & n6735 ) ;
  assign n6737 = n6735 ^ n6706 ^ n6637 ;
  assign n6738 = x85 & n5499 ;
  assign n6739 = ( x87 & n5497 ) | ( x87 & n6738 ) | ( n5497 & n6738 ) ;
  assign n6740 = n6738 | n6739 ;
  assign n6741 = x86 & ~n5502 ;
  assign n6742 = ( x86 & n6740 ) | ( x86 & ~n6741 ) | ( n6740 & ~n6741 ) ;
  assign n6743 = n1484 & n5501 ;
  assign n6744 = n6742 | n6743 ;
  assign n6745 = n6744 ^ x11 ^ 1'b0 ;
  assign n6746 = ( n5432 & n6697 ) | ( n5432 & n6745 ) | ( n6697 & n6745 ) ;
  assign n6747 = n6745 ^ n6697 ^ n5432 ;
  assign n6748 = x85 & n5718 ;
  assign n6749 = ( x87 & n5720 ) | ( x87 & n6748 ) | ( n5720 & n6748 ) ;
  assign n6750 = n6748 | n6749 ;
  assign n6751 = x86 & ~n5727 ;
  assign n6752 = ( x86 & n6750 ) | ( x86 & ~n6751 ) | ( n6750 & ~n6751 ) ;
  assign n6753 = n1484 & n5726 ;
  assign n6754 = n6752 | n6753 ;
  assign n6755 = n6754 ^ x8 ^ 1'b0 ;
  assign n6756 = n6755 ^ n6533 ^ n5945 ;
  assign n6757 = ( n5945 & n6533 ) | ( n5945 & n6755 ) | ( n6533 & n6755 ) ;
  assign n6758 = x88 & n4616 ;
  assign n6759 = ( x90 & n4606 ) | ( x90 & n6758 ) | ( n4606 & n6758 ) ;
  assign n6760 = n6758 | n6759 ;
  assign n6761 = x89 & ~n4605 ;
  assign n6762 = ( x89 & n6760 ) | ( x89 & ~n6761 ) | ( n6760 & ~n6761 ) ;
  assign n6763 = n1741 & n4608 ;
  assign n6764 = n6762 | n6763 ;
  assign n6765 = n6764 ^ x23 ^ 1'b0 ;
  assign n6766 = ( n3965 & n6646 ) | ( n3965 & n6765 ) | ( n6646 & n6765 ) ;
  assign n6767 = n6765 ^ n6646 ^ n3965 ;
  assign n6768 = x89 & n4972 ;
  assign n6769 = ( x91 & n4985 ) | ( x91 & n6768 ) | ( n4985 & n6768 ) ;
  assign n6770 = n6768 | n6769 ;
  assign n6771 = x90 & ~n4980 ;
  assign n6772 = ( x90 & n6770 ) | ( x90 & ~n6771 ) | ( n6770 & ~n6771 ) ;
  assign n6773 = n2114 & n4987 ;
  assign n6774 = n6772 | n6773 ;
  assign n6775 = n6774 ^ x14 ^ 1'b0 ;
  assign n6776 = n6775 ^ n6616 ^ n5493 ;
  assign n6777 = ( n5493 & n6616 ) | ( n5493 & n6775 ) | ( n6616 & n6775 ) ;
  assign n6778 = x86 & n5499 ;
  assign n6779 = ( x88 & n5497 ) | ( x88 & n6778 ) | ( n5497 & n6778 ) ;
  assign n6780 = n6778 | n6779 ;
  assign n6781 = x87 & ~n5502 ;
  assign n6782 = ( x87 & n6780 ) | ( x87 & ~n6781 ) | ( n6780 & ~n6781 ) ;
  assign n6783 = n1569 & n5501 ;
  assign n6784 = n6782 | n6783 ;
  assign n6785 = n6784 ^ x11 ^ 1'b0 ;
  assign n6786 = n6785 ^ n6746 ^ n5443 ;
  assign n6787 = ( n5443 & n6746 ) | ( n5443 & n6785 ) | ( n6746 & n6785 ) ;
  assign n6788 = x90 & n4972 ;
  assign n6789 = ( x92 & n4985 ) | ( x92 & n6788 ) | ( n4985 & n6788 ) ;
  assign n6790 = n6788 | n6789 ;
  assign n6791 = x91 & ~n4980 ;
  assign n6792 = ( x91 & n6790 ) | ( x91 & ~n6791 ) | ( n6790 & ~n6791 ) ;
  assign n6793 = n2420 & n4987 ;
  assign n6794 = n6792 | n6793 ;
  assign n6795 = n6794 ^ x14 ^ 1'b0 ;
  assign n6796 = ( n6627 & n6777 ) | ( n6627 & n6795 ) | ( n6777 & n6795 ) ;
  assign n6797 = n6795 ^ n6777 ^ n6627 ;
  assign n6798 = x87 & n5499 ;
  assign n6799 = ( x89 & n5497 ) | ( x89 & n6798 ) | ( n5497 & n6798 ) ;
  assign n6800 = n6798 | n6799 ;
  assign n6801 = x88 & ~n5502 ;
  assign n6802 = ( x88 & n6800 ) | ( x88 & ~n6801 ) | ( n6800 & ~n6801 ) ;
  assign n6803 = n1654 & n5501 ;
  assign n6804 = n6802 | n6803 ;
  assign n6805 = n6804 ^ x11 ^ 1'b0 ;
  assign n6806 = n6805 ^ n6787 ^ n5453 ;
  assign n6807 = ( n5453 & n6787 ) | ( n5453 & n6805 ) | ( n6787 & n6805 ) ;
  assign n6808 = x88 & n5499 ;
  assign n6809 = ( x90 & n5497 ) | ( x90 & n6808 ) | ( n5497 & n6808 ) ;
  assign n6810 = n6808 | n6809 ;
  assign n6811 = x89 & ~n5502 ;
  assign n6812 = ( x89 & n6810 ) | ( x89 & ~n6811 ) | ( n6810 & ~n6811 ) ;
  assign n6813 = n1741 & n5501 ;
  assign n6814 = n6812 | n6813 ;
  assign n6815 = n6814 ^ x11 ^ 1'b0 ;
  assign n6816 = ( n5462 & n6807 ) | ( n5462 & n6815 ) | ( n6807 & n6815 ) ;
  assign n6817 = n6815 ^ n6807 ^ n5462 ;
  assign n6818 = x91 & n4972 ;
  assign n6819 = ( x93 & n4985 ) | ( x93 & n6818 ) | ( n4985 & n6818 ) ;
  assign n6820 = n6818 | n6819 ;
  assign n6821 = x92 & ~n4980 ;
  assign n6822 = ( x92 & n6820 ) | ( x92 & ~n6821 ) | ( n6820 & ~n6821 ) ;
  assign n6823 = n2476 & n4987 ;
  assign n6824 = n6822 | n6823 ;
  assign n6825 = n6824 ^ x14 ^ 1'b0 ;
  assign n6826 = ( n6676 & n6796 ) | ( n6676 & n6825 ) | ( n6796 & n6825 ) ;
  assign n6827 = n6825 ^ n6796 ^ n6676 ;
  assign n6828 = x89 & n5499 ;
  assign n6829 = ( x91 & n5497 ) | ( x91 & n6828 ) | ( n5497 & n6828 ) ;
  assign n6830 = n6828 | n6829 ;
  assign n6831 = x90 & ~n5502 ;
  assign n6832 = ( x90 & n6830 ) | ( x90 & ~n6831 ) | ( n6830 & ~n6831 ) ;
  assign n6833 = n2114 & n5501 ;
  assign n6834 = n6832 | n6833 ;
  assign n6835 = n6834 ^ x11 ^ 1'b0 ;
  assign n6836 = n6835 ^ n6816 ^ n5473 ;
  assign n6837 = ( n5473 & n6816 ) | ( n5473 & n6835 ) | ( n6816 & n6835 ) ;
  assign n6838 = x92 & n4972 ;
  assign n6839 = ( x94 & n4985 ) | ( x94 & n6838 ) | ( n4985 & n6838 ) ;
  assign n6840 = n6838 | n6839 ;
  assign n6841 = x93 & ~n4980 ;
  assign n6842 = ( x93 & n6840 ) | ( x93 & ~n6841 ) | ( n6840 & ~n6841 ) ;
  assign n6843 = n2518 & n4987 ;
  assign n6844 = n6842 | n6843 ;
  assign n6845 = n6844 ^ x14 ^ 1'b0 ;
  assign n6846 = n6845 ^ n6826 ^ n6716 ;
  assign n6847 = ( n6716 & n6826 ) | ( n6716 & n6845 ) | ( n6826 & n6845 ) ;
  assign n6848 = x91 & n5011 ;
  assign n6849 = ( x93 & n5012 ) | ( x93 & n6848 ) | ( n5012 & n6848 ) ;
  assign n6850 = n6848 | n6849 ;
  assign n6851 = x92 & ~n5008 ;
  assign n6852 = ( x92 & n6850 ) | ( x92 & ~n6851 ) | ( n6850 & ~n6851 ) ;
  assign n6853 = n2476 & n5020 ;
  assign n6854 = n6852 | n6853 ;
  assign n6855 = n6854 ^ x17 ^ 1'b0 ;
  assign n6856 = n6855 ^ n6727 ^ n6707 ;
  assign n6857 = ( n6707 & n6727 ) | ( n6707 & n6855 ) | ( n6727 & n6855 ) ;
  assign n6858 = x92 & n5011 ;
  assign n6859 = ( x94 & n5012 ) | ( x94 & n6858 ) | ( n5012 & n6858 ) ;
  assign n6860 = n6858 | n6859 ;
  assign n6861 = x93 & ~n5008 ;
  assign n6862 = ( x93 & n6860 ) | ( x93 & ~n6861 ) | ( n6860 & ~n6861 ) ;
  assign n6863 = n2518 & n5020 ;
  assign n6864 = n6862 | n6863 ;
  assign n6865 = n6864 ^ x17 ^ 1'b0 ;
  assign n6866 = ( n6737 & n6857 ) | ( n6737 & n6865 ) | ( n6857 & n6865 ) ;
  assign n6867 = n6865 ^ n6857 ^ n6737 ;
  assign n6868 = x89 & n4616 ;
  assign n6869 = ( x91 & n4606 ) | ( x91 & n6868 ) | ( n4606 & n6868 ) ;
  assign n6870 = n6868 | n6869 ;
  assign n6871 = x90 & ~n4605 ;
  assign n6872 = ( x90 & n6870 ) | ( x90 & ~n6871 ) | ( n6870 & ~n6871 ) ;
  assign n6873 = n2114 & n4608 ;
  assign n6874 = n6872 | n6873 ;
  assign n6875 = n6874 ^ x23 ^ 1'b0 ;
  assign n6876 = ( n3975 & n6766 ) | ( n3975 & n6875 ) | ( n6766 & n6875 ) ;
  assign n6877 = n6875 ^ n6766 ^ n3975 ;
  assign n6878 = x90 & n4616 ;
  assign n6879 = ( x92 & n4606 ) | ( x92 & n6878 ) | ( n4606 & n6878 ) ;
  assign n6880 = n6878 | n6879 ;
  assign n6881 = x91 & ~n4605 ;
  assign n6882 = ( x91 & n6880 ) | ( x91 & ~n6881 ) | ( n6880 & ~n6881 ) ;
  assign n6883 = n2420 & n4608 ;
  assign n6884 = n6882 | n6883 ;
  assign n6885 = n6884 ^ x23 ^ 1'b0 ;
  assign n6886 = n6885 ^ n6876 ^ n3986 ;
  assign n6887 = ( n3986 & n6876 ) | ( n3986 & n6885 ) | ( n6876 & n6885 ) ;
  assign n6888 = x90 & n4790 ;
  assign n6889 = ( x92 & n4792 ) | ( x92 & n6888 ) | ( n4792 & n6888 ) ;
  assign n6890 = n6888 | n6889 ;
  assign n6891 = x91 & ~n4786 ;
  assign n6892 = ( x91 & n6890 ) | ( x91 & ~n6891 ) | ( n6890 & ~n6891 ) ;
  assign n6893 = n2420 & n4787 ;
  assign n6894 = n6892 | n6893 ;
  assign n6895 = n6894 ^ x20 ^ 1'b0 ;
  assign n6896 = ( n6647 & n6736 ) | ( n6647 & n6895 ) | ( n6736 & n6895 ) ;
  assign n6897 = n6895 ^ n6736 ^ n6647 ;
  assign n6898 = x93 & n5011 ;
  assign n6899 = ( x95 & n5012 ) | ( x95 & n6898 ) | ( n5012 & n6898 ) ;
  assign n6900 = n6898 | n6899 ;
  assign n6901 = x94 & ~n5008 ;
  assign n6902 = ( x94 & n6900 ) | ( x94 & ~n6901 ) | ( n6900 & ~n6901 ) ;
  assign n6903 = n2854 & n5020 ;
  assign n6904 = n6902 | n6903 ;
  assign n6905 = n6904 ^ x17 ^ 1'b0 ;
  assign n6906 = ( n6866 & n6897 ) | ( n6866 & n6905 ) | ( n6897 & n6905 ) ;
  assign n6907 = n6905 ^ n6897 ^ n6866 ;
  assign n6908 = x91 & n4790 ;
  assign n6909 = ( x93 & n4792 ) | ( x93 & n6908 ) | ( n4792 & n6908 ) ;
  assign n6910 = n6908 | n6909 ;
  assign n6911 = x92 & ~n4786 ;
  assign n6912 = ( x92 & n6910 ) | ( x92 & ~n6911 ) | ( n6910 & ~n6911 ) ;
  assign n6913 = n2476 & n4787 ;
  assign n6914 = n6912 | n6913 ;
  assign n6915 = n6914 ^ x20 ^ 1'b0 ;
  assign n6916 = ( n6767 & n6896 ) | ( n6767 & n6915 ) | ( n6896 & n6915 ) ;
  assign n6917 = n6915 ^ n6896 ^ n6767 ;
  assign n6918 = x92 & n4790 ;
  assign n6919 = ( x94 & n4792 ) | ( x94 & n6918 ) | ( n4792 & n6918 ) ;
  assign n6920 = n6918 | n6919 ;
  assign n6921 = x93 & ~n4786 ;
  assign n6922 = ( x93 & n6920 ) | ( x93 & ~n6921 ) | ( n6920 & ~n6921 ) ;
  assign n6923 = n2518 & n4787 ;
  assign n6924 = n6922 | n6923 ;
  assign n6925 = n6924 ^ x20 ^ 1'b0 ;
  assign n6926 = ( n6877 & n6916 ) | ( n6877 & n6925 ) | ( n6916 & n6925 ) ;
  assign n6927 = n6925 ^ n6916 ^ n6877 ;
  assign n6928 = x93 & n4790 ;
  assign n6929 = ( x95 & n4792 ) | ( x95 & n6928 ) | ( n4792 & n6928 ) ;
  assign n6930 = n6928 | n6929 ;
  assign n6931 = x94 & ~n4786 ;
  assign n6932 = ( x94 & n6930 ) | ( x94 & ~n6931 ) | ( n6930 & ~n6931 ) ;
  assign n6933 = n2854 & n4787 ;
  assign n6934 = n6932 | n6933 ;
  assign n6935 = n6934 ^ x20 ^ 1'b0 ;
  assign n6936 = n6935 ^ n6926 ^ n6886 ;
  assign n6937 = ( n6886 & n6926 ) | ( n6886 & n6935 ) | ( n6926 & n6935 ) ;
  assign n6938 = x94 & n5011 ;
  assign n6939 = ( x96 & n5012 ) | ( x96 & n6938 ) | ( n5012 & n6938 ) ;
  assign n6940 = n6938 | n6939 ;
  assign n6941 = x95 & ~n5008 ;
  assign n6942 = ( x95 & n6940 ) | ( x95 & ~n6941 ) | ( n6940 & ~n6941 ) ;
  assign n6943 = n2907 & n5020 ;
  assign n6944 = n6942 | n6943 ;
  assign n6945 = n6944 ^ x17 ^ 1'b0 ;
  assign n6946 = n6945 ^ n6917 ^ n6906 ;
  assign n6947 = ( n6906 & n6917 ) | ( n6906 & n6945 ) | ( n6917 & n6945 ) ;
  assign n6948 = x86 & n5718 ;
  assign n6949 = ( x88 & n5720 ) | ( x88 & n6948 ) | ( n5720 & n6948 ) ;
  assign n6950 = n6948 | n6949 ;
  assign n6951 = x87 & ~n5727 ;
  assign n6952 = ( x87 & n6950 ) | ( x87 & ~n6951 ) | ( n6950 & ~n6951 ) ;
  assign n6953 = n1569 & n5726 ;
  assign n6954 = n6952 | n6953 ;
  assign n6955 = n6954 ^ x8 ^ 1'b0 ;
  assign n6956 = n6955 ^ n6757 ^ n6554 ;
  assign n6957 = ( n6554 & n6757 ) | ( n6554 & n6955 ) | ( n6757 & n6955 ) ;
  assign n6958 = x87 & n5718 ;
  assign n6959 = ( x89 & n5720 ) | ( x89 & n6958 ) | ( n5720 & n6958 ) ;
  assign n6960 = n6958 | n6959 ;
  assign n6961 = x88 & ~n5727 ;
  assign n6962 = ( x88 & n6960 ) | ( x88 & ~n6961 ) | ( n6960 & ~n6961 ) ;
  assign n6963 = n1654 & n5726 ;
  assign n6964 = n6962 | n6963 ;
  assign n6965 = n6964 ^ x8 ^ 1'b0 ;
  assign n6966 = n6965 ^ n6957 ^ n6696 ;
  assign n6967 = ( n6696 & n6957 ) | ( n6696 & n6965 ) | ( n6957 & n6965 ) ;
  assign n6968 = x95 & n5011 ;
  assign n6969 = ( x97 & n5012 ) | ( x97 & n6968 ) | ( n5012 & n6968 ) ;
  assign n6970 = n6968 | n6969 ;
  assign n6971 = x96 & ~n5008 ;
  assign n6972 = ( x96 & n6970 ) | ( x96 & ~n6971 ) | ( n6970 & ~n6971 ) ;
  assign n6973 = n3668 & n5020 ;
  assign n6974 = n6972 | n6973 ;
  assign n6975 = n6974 ^ x17 ^ 1'b0 ;
  assign n6976 = n6975 ^ n6947 ^ n6927 ;
  assign n6977 = ( n6927 & n6947 ) | ( n6927 & n6975 ) | ( n6947 & n6975 ) ;
  assign n6978 = x93 & n4972 ;
  assign n6979 = ( x95 & n4985 ) | ( x95 & n6978 ) | ( n4985 & n6978 ) ;
  assign n6980 = n6978 | n6979 ;
  assign n6981 = x94 & ~n4980 ;
  assign n6982 = ( x94 & n6980 ) | ( x94 & ~n6981 ) | ( n6980 & ~n6981 ) ;
  assign n6983 = n2854 & n4987 ;
  assign n6984 = n6982 | n6983 ;
  assign n6985 = n6984 ^ x14 ^ 1'b0 ;
  assign n6986 = ( n6726 & n6847 ) | ( n6726 & n6985 ) | ( n6847 & n6985 ) ;
  assign n6987 = n6985 ^ n6847 ^ n6726 ;
  assign n6988 = x90 & n5499 ;
  assign n6989 = ( x92 & n5497 ) | ( x92 & n6988 ) | ( n5497 & n6988 ) ;
  assign n6990 = n6988 | n6989 ;
  assign n6991 = x91 & ~n5502 ;
  assign n6992 = ( x91 & n6990 ) | ( x91 & ~n6991 ) | ( n6990 & ~n6991 ) ;
  assign n6993 = n2420 & n5501 ;
  assign n6994 = n6992 | n6993 ;
  assign n6995 = n6994 ^ x11 ^ 1'b0 ;
  assign n6996 = ( n5482 & n6837 ) | ( n5482 & n6995 ) | ( n6837 & n6995 ) ;
  assign n6997 = n6995 ^ n6837 ^ n5482 ;
  assign n6998 = x88 & n5718 ;
  assign n6999 = ( x90 & n5720 ) | ( x90 & n6998 ) | ( n5720 & n6998 ) ;
  assign n7000 = n6998 | n6999 ;
  assign n7001 = x89 & ~n5727 ;
  assign n7002 = ( x89 & n7000 ) | ( x89 & ~n7001 ) | ( n7000 & ~n7001 ) ;
  assign n7003 = n1741 & n5726 ;
  assign n7004 = n7002 | n7003 ;
  assign n7005 = n7004 ^ x8 ^ 1'b0 ;
  assign n7006 = ( n6747 & n6967 ) | ( n6747 & n7005 ) | ( n6967 & n7005 ) ;
  assign n7007 = n7005 ^ n6967 ^ n6747 ;
  assign n7008 = x91 & n5499 ;
  assign n7009 = ( x93 & n5497 ) | ( x93 & n7008 ) | ( n5497 & n7008 ) ;
  assign n7010 = n7008 | n7009 ;
  assign n7011 = x92 & ~n5502 ;
  assign n7012 = ( x92 & n7010 ) | ( x92 & ~n7011 ) | ( n7010 & ~n7011 ) ;
  assign n7013 = n2476 & n5501 ;
  assign n7014 = n7012 | n7013 ;
  assign n7015 = n7014 ^ x11 ^ 1'b0 ;
  assign n7016 = n7015 ^ n6996 ^ n5492 ;
  assign n7017 = ( n5492 & n6996 ) | ( n5492 & n7015 ) | ( n6996 & n7015 ) ;
  assign n7018 = x92 & n5499 ;
  assign n7019 = ( x94 & n5497 ) | ( x94 & n7018 ) | ( n5497 & n7018 ) ;
  assign n7020 = n7018 | n7019 ;
  assign n7021 = x93 & ~n5502 ;
  assign n7022 = ( x93 & n7020 ) | ( x93 & ~n7021 ) | ( n7020 & ~n7021 ) ;
  assign n7023 = n2518 & n5501 ;
  assign n7024 = n7022 | n7023 ;
  assign n7025 = n7024 ^ x11 ^ 1'b0 ;
  assign n7026 = n7025 ^ n7017 ^ n6776 ;
  assign n7027 = ( n6776 & n7017 ) | ( n6776 & n7025 ) | ( n7017 & n7025 ) ;
  assign n7028 = x93 & n5499 ;
  assign n7029 = ( x95 & n5497 ) | ( x95 & n7028 ) | ( n5497 & n7028 ) ;
  assign n7030 = n7028 | n7029 ;
  assign n7031 = x94 & ~n5502 ;
  assign n7032 = ( x94 & n7030 ) | ( x94 & ~n7031 ) | ( n7030 & ~n7031 ) ;
  assign n7033 = n2854 & n5501 ;
  assign n7034 = n7032 | n7033 ;
  assign n7035 = n7034 ^ x11 ^ 1'b0 ;
  assign n7036 = n7035 ^ n7027 ^ n6797 ;
  assign n7037 = ( n6797 & n7027 ) | ( n6797 & n7035 ) | ( n7027 & n7035 ) ;
  assign n7038 = x94 & n5499 ;
  assign n7039 = ( x96 & n5497 ) | ( x96 & n7038 ) | ( n5497 & n7038 ) ;
  assign n7040 = n7038 | n7039 ;
  assign n7041 = x95 & ~n5502 ;
  assign n7042 = ( x95 & n7040 ) | ( x95 & ~n7041 ) | ( n7040 & ~n7041 ) ;
  assign n7043 = n2907 & n5501 ;
  assign n7044 = n7042 | n7043 ;
  assign n7045 = n7044 ^ x11 ^ 1'b0 ;
  assign n7046 = ( n6827 & n7037 ) | ( n6827 & n7045 ) | ( n7037 & n7045 ) ;
  assign n7047 = n7045 ^ n7037 ^ n6827 ;
  assign n7048 = x89 & n5718 ;
  assign n7049 = ( x91 & n5720 ) | ( x91 & n7048 ) | ( n5720 & n7048 ) ;
  assign n7050 = n7048 | n7049 ;
  assign n7051 = x90 & ~n5727 ;
  assign n7052 = ( x90 & n7050 ) | ( x90 & ~n7051 ) | ( n7050 & ~n7051 ) ;
  assign n7053 = n2114 & n5726 ;
  assign n7054 = n7052 | n7053 ;
  assign n7055 = n7054 ^ x8 ^ 1'b0 ;
  assign n7056 = ( n6786 & n7006 ) | ( n6786 & n7055 ) | ( n7006 & n7055 ) ;
  assign n7057 = n7055 ^ n7006 ^ n6786 ;
  assign n7058 = x90 & n5718 ;
  assign n7059 = ( x92 & n5720 ) | ( x92 & n7058 ) | ( n5720 & n7058 ) ;
  assign n7060 = n7058 | n7059 ;
  assign n7061 = x91 & ~n5727 ;
  assign n7062 = ( x91 & n7060 ) | ( x91 & ~n7061 ) | ( n7060 & ~n7061 ) ;
  assign n7063 = n2420 & n5726 ;
  assign n7064 = n7062 | n7063 ;
  assign n7065 = n7064 ^ x8 ^ 1'b0 ;
  assign n7066 = ( n6806 & n7056 ) | ( n6806 & n7065 ) | ( n7056 & n7065 ) ;
  assign n7067 = n7065 ^ n7056 ^ n6806 ;
  assign n7068 = x91 & n6104 ;
  assign n7069 = ( x93 & n6105 ) | ( x93 & n7068 ) | ( n6105 & n7068 ) ;
  assign n7070 = x88 & n5979 ;
  assign n7071 = x89 & ~n5970 ;
  assign n7072 = n7068 | n7069 ;
  assign n7073 = x92 & ~n5727 ;
  assign n7074 = ( x90 & n5969 ) | ( x90 & n7070 ) | ( n5969 & n7070 ) ;
  assign n7075 = n7070 | n7074 ;
  assign n7076 = x91 & n5718 ;
  assign n7077 = ( x93 & n5720 ) | ( x93 & n7076 ) | ( n5720 & n7076 ) ;
  assign n7078 = n7076 | n7077 ;
  assign n7079 = ( x92 & ~n7073 ) | ( x92 & n7078 ) | ( ~n7073 & n7078 ) ;
  assign n7080 = x92 & ~n6107 ;
  assign n7081 = ( x92 & n7072 ) | ( x92 & ~n7080 ) | ( n7072 & ~n7080 ) ;
  assign n7082 = ( x89 & ~n7071 ) | ( x89 & n7075 ) | ( ~n7071 & n7075 ) ;
  assign n7083 = n1741 & n5968 ;
  assign n7084 = n2476 & n5726 ;
  assign n7085 = n7082 | n7083 ;
  assign n7086 = n7085 ^ x5 ^ 1'b0 ;
  assign n7087 = n2476 & ~n6108 ;
  assign n7088 = n7079 | n7084 ;
  assign n7089 = n7088 ^ x8 ^ 1'b0 ;
  assign n7090 = n7089 ^ n7066 ^ n6817 ;
  assign n7091 = ( n6817 & n7066 ) | ( n6817 & n7089 ) | ( n7066 & n7089 ) ;
  assign n7092 = x89 & n5979 ;
  assign n7093 = ( x91 & n5969 ) | ( x91 & n7092 ) | ( n5969 & n7092 ) ;
  assign n7094 = ( n2476 & n7081 ) | ( n2476 & ~n7087 ) | ( n7081 & ~n7087 ) ;
  assign n7095 = n7094 ^ x2 ^ 1'b0 ;
  assign n7096 = n7086 ^ n6756 ^ n6498 ;
  assign n7097 = ( n6508 & n7095 ) | ( n6508 & n7096 ) | ( n7095 & n7096 ) ;
  assign n7098 = n7092 | n7093 ;
  assign n7099 = x90 & ~n5970 ;
  assign n7100 = ( x90 & n7098 ) | ( x90 & ~n7099 ) | ( n7098 & ~n7099 ) ;
  assign n7101 = n2114 & n5968 ;
  assign n7102 = n7100 | n7101 ;
  assign n7103 = ( n6498 & n6756 ) | ( n6498 & n7086 ) | ( n6756 & n7086 ) ;
  assign n7104 = n7102 ^ x5 ^ 1'b0 ;
  assign n7105 = n7104 ^ n7103 ^ n6956 ;
  assign n7106 = x90 & n5979 ;
  assign n7107 = ( x92 & n5969 ) | ( x92 & n7106 ) | ( n5969 & n7106 ) ;
  assign n7108 = n7106 | n7107 ;
  assign n7109 = n7096 ^ n7095 ^ n6508 ;
  assign n7110 = x93 & n5718 ;
  assign n7111 = ( x95 & n5720 ) | ( x95 & n7110 ) | ( n5720 & n7110 ) ;
  assign n7112 = n7110 | n7111 ;
  assign n7113 = x91 & ~n5970 ;
  assign n7114 = x93 & ~n5727 ;
  assign n7115 = ( x91 & n7108 ) | ( x91 & ~n7113 ) | ( n7108 & ~n7113 ) ;
  assign n7116 = n2420 & n5968 ;
  assign n7117 = n7115 | n7116 ;
  assign n7118 = x94 & ~n5727 ;
  assign n7119 = ( n6956 & n7103 ) | ( n6956 & n7104 ) | ( n7103 & n7104 ) ;
  assign n7120 = ( x94 & n7112 ) | ( x94 & ~n7118 ) | ( n7112 & ~n7118 ) ;
  assign n7121 = n2854 & n5726 ;
  assign n7122 = n3668 & n5501 ;
  assign n7123 = n7120 | n7121 ;
  assign n7124 = n7117 ^ x5 ^ 1'b0 ;
  assign n7125 = n7124 ^ n7119 ^ n6966 ;
  assign n7126 = ( n6966 & n7119 ) | ( n6966 & n7124 ) | ( n7119 & n7124 ) ;
  assign n7127 = x92 & n5718 ;
  assign n7128 = x96 & ~n5502 ;
  assign n7129 = ( x94 & n5720 ) | ( x94 & n7127 ) | ( n5720 & n7127 ) ;
  assign n7130 = n7127 | n7129 ;
  assign n7131 = n2518 & n5726 ;
  assign n7132 = n7123 ^ x8 ^ 1'b0 ;
  assign n7133 = ( x93 & ~n7114 ) | ( x93 & n7130 ) | ( ~n7114 & n7130 ) ;
  assign n7134 = x95 & n5499 ;
  assign n7135 = n7131 | n7133 ;
  assign n7136 = ( x97 & n5497 ) | ( x97 & n7134 ) | ( n5497 & n7134 ) ;
  assign n7137 = n7134 | n7136 ;
  assign n7138 = ( x96 & ~n7128 ) | ( x96 & n7137 ) | ( ~n7128 & n7137 ) ;
  assign n7139 = n7122 | n7138 ;
  assign n7140 = n7135 ^ x8 ^ 1'b0 ;
  assign n7141 = ( n6836 & n7091 ) | ( n6836 & n7140 ) | ( n7091 & n7140 ) ;
  assign n7142 = n7141 ^ n7132 ^ n6997 ;
  assign n7143 = n7140 ^ n7091 ^ n6836 ;
  assign n7144 = n7139 ^ x11 ^ 1'b0 ;
  assign n7145 = n7144 ^ n7046 ^ n6846 ;
  assign n7146 = ( n6846 & n7046 ) | ( n6846 & n7144 ) | ( n7046 & n7144 ) ;
  assign n7147 = ( n6997 & n7132 ) | ( n6997 & n7141 ) | ( n7132 & n7141 ) ;
  assign n7148 = x94 & n4972 ;
  assign n7149 = ( x96 & n4985 ) | ( x96 & n7148 ) | ( n4985 & n7148 ) ;
  assign n7150 = n7148 | n7149 ;
  assign n7151 = x95 & ~n4980 ;
  assign n7152 = ( x95 & n7150 ) | ( x95 & ~n7151 ) | ( n7150 & ~n7151 ) ;
  assign n7153 = n2907 & n4987 ;
  assign n7154 = n7152 | n7153 ;
  assign n7155 = n7154 ^ x14 ^ 1'b0 ;
  assign n7156 = ( n6856 & n6986 ) | ( n6856 & n7155 ) | ( n6986 & n7155 ) ;
  assign n7157 = n7155 ^ n6986 ^ n6856 ;
  assign n7158 = x91 & n5979 ;
  assign n7159 = ( x93 & n5969 ) | ( x93 & n7158 ) | ( n5969 & n7158 ) ;
  assign n7160 = n7158 | n7159 ;
  assign n7161 = x92 & ~n5970 ;
  assign n7162 = ( x92 & n7160 ) | ( x92 & ~n7161 ) | ( n7160 & ~n7161 ) ;
  assign n7163 = n2476 & n5968 ;
  assign n7164 = n7162 | n7163 ;
  assign n7165 = n7164 ^ x5 ^ 1'b0 ;
  assign n7166 = ( n7007 & n7126 ) | ( n7007 & n7165 ) | ( n7126 & n7165 ) ;
  assign n7167 = n7165 ^ n7126 ^ n7007 ;
  assign n7168 = x95 & n4972 ;
  assign n7169 = ( x97 & n4985 ) | ( x97 & n7168 ) | ( n4985 & n7168 ) ;
  assign n7170 = n7168 | n7169 ;
  assign n7171 = x96 & ~n4980 ;
  assign n7172 = ( x96 & n7170 ) | ( x96 & ~n7171 ) | ( n7170 & ~n7171 ) ;
  assign n7173 = n3668 & n4987 ;
  assign n7174 = n7172 | n7173 ;
  assign n7175 = n7174 ^ x14 ^ 1'b0 ;
  assign n7176 = n7175 ^ n7156 ^ n6867 ;
  assign n7177 = ( n6867 & n7156 ) | ( n6867 & n7175 ) | ( n7156 & n7175 ) ;
  assign n7178 = x92 & n5979 ;
  assign n7179 = ( x94 & n5969 ) | ( x94 & n7178 ) | ( n5969 & n7178 ) ;
  assign n7180 = n7178 | n7179 ;
  assign n7181 = x93 & ~n5970 ;
  assign n7182 = ( x93 & n7180 ) | ( x93 & ~n7181 ) | ( n7180 & ~n7181 ) ;
  assign n7183 = n2518 & n5968 ;
  assign n7184 = n7182 | n7183 ;
  assign n7185 = n7184 ^ x5 ^ 1'b0 ;
  assign n7186 = n7185 ^ n7166 ^ n7057 ;
  assign n7187 = ( n7057 & n7166 ) | ( n7057 & n7185 ) | ( n7166 & n7185 ) ;
  assign n7188 = x93 & n5979 ;
  assign n7189 = ( x95 & n5969 ) | ( x95 & n7188 ) | ( n5969 & n7188 ) ;
  assign n7190 = n7188 | n7189 ;
  assign n7191 = x94 & ~n5970 ;
  assign n7192 = ( x94 & n7190 ) | ( x94 & ~n7191 ) | ( n7190 & ~n7191 ) ;
  assign n7193 = n2854 & n5968 ;
  assign n7194 = n7192 | n7193 ;
  assign n7195 = n7194 ^ x5 ^ 1'b0 ;
  assign n7196 = n7195 ^ n7187 ^ n7067 ;
  assign n7197 = ( n7067 & n7187 ) | ( n7067 & n7195 ) | ( n7187 & n7195 ) ;
  assign n7198 = x94 & n5979 ;
  assign n7199 = ( x96 & n5969 ) | ( x96 & n7198 ) | ( n5969 & n7198 ) ;
  assign n7200 = n7198 | n7199 ;
  assign n7201 = x95 & ~n5970 ;
  assign n7202 = ( x95 & n7200 ) | ( x95 & ~n7201 ) | ( n7200 & ~n7201 ) ;
  assign n7203 = n2907 & n5968 ;
  assign n7204 = n7202 | n7203 ;
  assign n7205 = n7204 ^ x5 ^ 1'b0 ;
  assign n7206 = ( n7090 & n7197 ) | ( n7090 & n7205 ) | ( n7197 & n7205 ) ;
  assign n7207 = n7205 ^ n7197 ^ n7090 ;
  assign n7208 = x95 & n5979 ;
  assign n7209 = ( x97 & n5969 ) | ( x97 & n7208 ) | ( n5969 & n7208 ) ;
  assign n7210 = n7208 | n7209 ;
  assign n7211 = x96 & ~n5970 ;
  assign n7212 = ( x96 & n7210 ) | ( x96 & ~n7211 ) | ( n7210 & ~n7211 ) ;
  assign n7213 = n3668 & n5968 ;
  assign n7214 = n7212 | n7213 ;
  assign n7215 = n7214 ^ x5 ^ 1'b0 ;
  assign n7216 = ( n7143 & n7206 ) | ( n7143 & n7215 ) | ( n7206 & n7215 ) ;
  assign n7217 = n7215 ^ n7206 ^ n7143 ;
  assign n7218 = x96 & n5979 ;
  assign n7219 = ( x98 & n5969 ) | ( x98 & n7218 ) | ( n5969 & n7218 ) ;
  assign n7220 = n7218 | n7219 ;
  assign n7221 = x97 & ~n5970 ;
  assign n7222 = ( x97 & n7220 ) | ( x97 & ~n7221 ) | ( n7220 & ~n7221 ) ;
  assign n7223 = n4052 & n5968 ;
  assign n7224 = n7222 | n7223 ;
  assign n7225 = n7224 ^ x5 ^ 1'b0 ;
  assign n7226 = n7225 ^ n7216 ^ n7142 ;
  assign n7227 = ( n7142 & n7216 ) | ( n7142 & n7225 ) | ( n7216 & n7225 ) ;
  assign n7228 = x94 & n5718 ;
  assign n7229 = ( x96 & n5720 ) | ( x96 & n7228 ) | ( n5720 & n7228 ) ;
  assign n7230 = n7228 | n7229 ;
  assign n7231 = x95 & ~n5727 ;
  assign n7232 = ( x95 & n7230 ) | ( x95 & ~n7231 ) | ( n7230 & ~n7231 ) ;
  assign n7233 = n2907 & n5726 ;
  assign n7234 = n7232 | n7233 ;
  assign n7235 = n7234 ^ x8 ^ 1'b0 ;
  assign n7236 = n7235 ^ n7147 ^ n7016 ;
  assign n7237 = ( n7016 & n7147 ) | ( n7016 & n7235 ) | ( n7147 & n7235 ) ;
  assign n7238 = x96 & n4972 ;
  assign n7239 = ( x98 & n4985 ) | ( x98 & n7238 ) | ( n4985 & n7238 ) ;
  assign n7240 = n7238 | n7239 ;
  assign n7241 = x97 & ~n4980 ;
  assign n7242 = ( x97 & n7240 ) | ( x97 & ~n7241 ) | ( n7240 & ~n7241 ) ;
  assign n7243 = n4052 & n4987 ;
  assign n7244 = n7242 | n7243 ;
  assign n7245 = n7244 ^ x14 ^ 1'b0 ;
  assign n7246 = n7245 ^ n7177 ^ n6907 ;
  assign n7247 = ( n6907 & n7177 ) | ( n6907 & n7245 ) | ( n7177 & n7245 ) ;
  assign n7248 = x97 & n4972 ;
  assign n7249 = ( x99 & n4985 ) | ( x99 & n7248 ) | ( n4985 & n7248 ) ;
  assign n7250 = n7248 | n7249 ;
  assign n7251 = x98 & ~n4980 ;
  assign n7252 = ( x98 & n7250 ) | ( x98 & ~n7251 ) | ( n7250 & ~n7251 ) ;
  assign n7253 = n4270 & n4987 ;
  assign n7254 = n7252 | n7253 ;
  assign n7255 = n7254 ^ x14 ^ 1'b0 ;
  assign n7256 = n7255 ^ n7247 ^ n6946 ;
  assign n7257 = ( n6946 & n7247 ) | ( n6946 & n7255 ) | ( n7247 & n7255 ) ;
  assign n7258 = x97 & n5979 ;
  assign n7259 = ( x99 & n5969 ) | ( x99 & n7258 ) | ( n5969 & n7258 ) ;
  assign n7260 = n7258 | n7259 ;
  assign n7261 = x98 & ~n5970 ;
  assign n7262 = ( x98 & n7260 ) | ( x98 & ~n7261 ) | ( n7260 & ~n7261 ) ;
  assign n7263 = n4270 & n5968 ;
  assign n7264 = n7262 | n7263 ;
  assign n7265 = n7264 ^ x5 ^ 1'b0 ;
  assign n7266 = n7265 ^ n7236 ^ n7227 ;
  assign n7267 = ( n7227 & n7236 ) | ( n7227 & n7265 ) | ( n7236 & n7265 ) ;
  assign n7268 = x95 & n5718 ;
  assign n7269 = ( x97 & n5720 ) | ( x97 & n7268 ) | ( n5720 & n7268 ) ;
  assign n7270 = n7268 | n7269 ;
  assign n7271 = x96 & ~n5727 ;
  assign n7272 = ( x96 & n7270 ) | ( x96 & ~n7271 ) | ( n7270 & ~n7271 ) ;
  assign n7273 = n3668 & n5726 ;
  assign n7274 = n7272 | n7273 ;
  assign n7275 = n7274 ^ x8 ^ 1'b0 ;
  assign n7276 = n7275 ^ n7237 ^ n7026 ;
  assign n7277 = ( n7026 & n7237 ) | ( n7026 & n7275 ) | ( n7237 & n7275 ) ;
  assign n7278 = x96 & n5718 ;
  assign n7279 = ( x98 & n5720 ) | ( x98 & n7278 ) | ( n5720 & n7278 ) ;
  assign n7280 = n7278 | n7279 ;
  assign n7281 = x97 & ~n5727 ;
  assign n7282 = ( x97 & n7280 ) | ( x97 & ~n7281 ) | ( n7280 & ~n7281 ) ;
  assign n7283 = n4052 & n5726 ;
  assign n7284 = n7282 | n7283 ;
  assign n7285 = n7284 ^ x8 ^ 1'b0 ;
  assign n7286 = ( n7036 & n7277 ) | ( n7036 & n7285 ) | ( n7277 & n7285 ) ;
  assign n7287 = n7285 ^ n7277 ^ n7036 ;
  assign n7288 = x96 & n5499 ;
  assign n7289 = ( x98 & n5497 ) | ( x98 & n7288 ) | ( n5497 & n7288 ) ;
  assign n7290 = n7288 | n7289 ;
  assign n7291 = x97 & ~n5502 ;
  assign n7292 = ( x97 & n7290 ) | ( x97 & ~n7291 ) | ( n7290 & ~n7291 ) ;
  assign n7293 = n4052 & n5501 ;
  assign n7294 = n7292 | n7293 ;
  assign n7295 = n7294 ^ x11 ^ 1'b0 ;
  assign n7296 = ( n6987 & n7146 ) | ( n6987 & n7295 ) | ( n7146 & n7295 ) ;
  assign n7297 = n7295 ^ n7146 ^ n6987 ;
  assign n7298 = x92 & n6104 ;
  assign n7299 = ( x94 & n6105 ) | ( x94 & n7298 ) | ( n6105 & n7298 ) ;
  assign n7300 = n7298 | n7299 ;
  assign n7301 = x93 & ~n6107 ;
  assign n7302 = ( x93 & n7300 ) | ( x93 & ~n7301 ) | ( n7300 & ~n7301 ) ;
  assign n7303 = n2518 & ~n6108 ;
  assign n7304 = ( n2518 & n7302 ) | ( n2518 & ~n7303 ) | ( n7302 & ~n7303 ) ;
  assign n7305 = n7304 ^ x2 ^ 1'b0 ;
  assign n7306 = ( n7097 & n7105 ) | ( n7097 & n7305 ) | ( n7105 & n7305 ) ;
  assign n7307 = n7305 ^ n7105 ^ n7097 ;
  assign n7308 = x97 & n5718 ;
  assign n7309 = ( x99 & n5720 ) | ( x99 & n7308 ) | ( n5720 & n7308 ) ;
  assign n7310 = n7308 | n7309 ;
  assign n7311 = x98 & ~n5727 ;
  assign n7312 = ( x98 & n7310 ) | ( x98 & ~n7311 ) | ( n7310 & ~n7311 ) ;
  assign n7313 = n4270 & n5726 ;
  assign n7314 = n7312 | n7313 ;
  assign n7315 = n7314 ^ x8 ^ 1'b0 ;
  assign n7316 = ( n7047 & n7286 ) | ( n7047 & n7315 ) | ( n7286 & n7315 ) ;
  assign n7317 = n7315 ^ n7286 ^ n7047 ;
  assign n7318 = x93 & n6104 ;
  assign n7319 = ( x95 & n6105 ) | ( x95 & n7318 ) | ( n6105 & n7318 ) ;
  assign n7320 = n7318 | n7319 ;
  assign n7321 = x94 & ~n6107 ;
  assign n7322 = ( x94 & n7320 ) | ( x94 & ~n7321 ) | ( n7320 & ~n7321 ) ;
  assign n7323 = n2854 & ~n6108 ;
  assign n7324 = ( n2854 & n7322 ) | ( n2854 & ~n7323 ) | ( n7322 & ~n7323 ) ;
  assign n7325 = n7324 ^ x2 ^ 1'b0 ;
  assign n7326 = n7325 ^ n7306 ^ n7125 ;
  assign n7327 = ( n7125 & n7306 ) | ( n7125 & n7325 ) | ( n7306 & n7325 ) ;
  assign n7328 = x94 & n6104 ;
  assign n7329 = ( x96 & n6105 ) | ( x96 & n7328 ) | ( n6105 & n7328 ) ;
  assign n7330 = n7328 | n7329 ;
  assign n7331 = x95 & ~n6107 ;
  assign n7332 = ( x95 & n7330 ) | ( x95 & ~n7331 ) | ( n7330 & ~n7331 ) ;
  assign n7333 = n2907 & ~n6108 ;
  assign n7334 = ( n2907 & n7332 ) | ( n2907 & ~n7333 ) | ( n7332 & ~n7333 ) ;
  assign n7335 = n7334 ^ x2 ^ 1'b0 ;
  assign n7336 = ( n7167 & n7327 ) | ( n7167 & n7335 ) | ( n7327 & n7335 ) ;
  assign n7337 = n7335 ^ n7327 ^ n7167 ;
  assign n7338 = x95 & n6104 ;
  assign n7339 = ( x97 & n6105 ) | ( x97 & n7338 ) | ( n6105 & n7338 ) ;
  assign n7340 = n7338 | n7339 ;
  assign n7341 = x96 & ~n6107 ;
  assign n7342 = ( x96 & n7340 ) | ( x96 & ~n7341 ) | ( n7340 & ~n7341 ) ;
  assign n7343 = n3668 & ~n6108 ;
  assign n7344 = ( n3668 & n7342 ) | ( n3668 & ~n7343 ) | ( n7342 & ~n7343 ) ;
  assign n7345 = n7344 ^ x2 ^ 1'b0 ;
  assign n7346 = n7345 ^ n7336 ^ n7186 ;
  assign n7347 = ( n7186 & n7336 ) | ( n7186 & n7345 ) | ( n7336 & n7345 ) ;
  assign n7348 = x96 & n6104 ;
  assign n7349 = ( x98 & n6105 ) | ( x98 & n7348 ) | ( n6105 & n7348 ) ;
  assign n7350 = n7348 | n7349 ;
  assign n7351 = x97 & ~n6107 ;
  assign n7352 = ( x97 & n7350 ) | ( x97 & ~n7351 ) | ( n7350 & ~n7351 ) ;
  assign n7353 = n4052 & ~n6108 ;
  assign n7354 = ( n4052 & n7352 ) | ( n4052 & ~n7353 ) | ( n7352 & ~n7353 ) ;
  assign n7355 = n7354 ^ x2 ^ 1'b0 ;
  assign n7356 = ( n7196 & n7347 ) | ( n7196 & n7355 ) | ( n7347 & n7355 ) ;
  assign n7357 = n7355 ^ n7347 ^ n7196 ;
  assign n7358 = x97 & n6104 ;
  assign n7359 = ( x99 & n6105 ) | ( x99 & n7358 ) | ( n6105 & n7358 ) ;
  assign n7360 = n7358 | n7359 ;
  assign n7361 = x98 & ~n6107 ;
  assign n7362 = ( x98 & n7360 ) | ( x98 & ~n7361 ) | ( n7360 & ~n7361 ) ;
  assign n7363 = n4270 & ~n6108 ;
  assign n7364 = ( n4270 & n7362 ) | ( n4270 & ~n7363 ) | ( n7362 & ~n7363 ) ;
  assign n7365 = n7364 ^ x2 ^ 1'b0 ;
  assign n7366 = ( n7207 & n7356 ) | ( n7207 & n7365 ) | ( n7356 & n7365 ) ;
  assign n7367 = n7365 ^ n7356 ^ n7207 ;
  assign n7368 = x98 & n5979 ;
  assign n7369 = ( x100 & n5969 ) | ( x100 & n7368 ) | ( n5969 & n7368 ) ;
  assign n7370 = n7368 | n7369 ;
  assign n7371 = x99 & ~n5970 ;
  assign n7372 = ( x99 & n7370 ) | ( x99 & ~n7371 ) | ( n7370 & ~n7371 ) ;
  assign n7373 = n4334 & n5968 ;
  assign n7374 = n7372 | n7373 ;
  assign n7375 = n7374 ^ x5 ^ 1'b0 ;
  assign n7376 = ( n7267 & n7276 ) | ( n7267 & n7375 ) | ( n7276 & n7375 ) ;
  assign n7377 = n7375 ^ n7276 ^ n7267 ;
  assign n7378 = x99 & n5979 ;
  assign n7379 = ( x101 & n5969 ) | ( x101 & n7378 ) | ( n5969 & n7378 ) ;
  assign n7380 = n7378 | n7379 ;
  assign n7381 = x100 & ~n5970 ;
  assign n7382 = ( x100 & n7380 ) | ( x100 & ~n7381 ) | ( n7380 & ~n7381 ) ;
  assign n7383 = n5687 & n5968 ;
  assign n7384 = n7382 | n7383 ;
  assign n7385 = n7384 ^ x5 ^ 1'b0 ;
  assign n7386 = n7385 ^ n7376 ^ n7287 ;
  assign n7387 = ( n7287 & n7376 ) | ( n7287 & n7385 ) | ( n7376 & n7385 ) ;
  assign n7388 = x100 & n5979 ;
  assign n7389 = ( x102 & n5969 ) | ( x102 & n7388 ) | ( n5969 & n7388 ) ;
  assign n7390 = n7388 | n7389 ;
  assign n7391 = x101 & ~n5970 ;
  assign n7392 = ( x101 & n7390 ) | ( x101 & ~n7391 ) | ( n7390 & ~n7391 ) ;
  assign n7393 = n5947 & n5968 ;
  assign n7394 = n7392 | n7393 ;
  assign n7395 = n7394 ^ x5 ^ 1'b0 ;
  assign n7396 = n7395 ^ n7387 ^ n7317 ;
  assign n7397 = ( n7317 & n7387 ) | ( n7317 & n7395 ) | ( n7387 & n7395 ) ;
  assign n7398 = x98 & n5718 ;
  assign n7399 = ( x100 & n5720 ) | ( x100 & n7398 ) | ( n5720 & n7398 ) ;
  assign n7400 = n7398 | n7399 ;
  assign n7401 = x99 & ~n5727 ;
  assign n7402 = ( x99 & n7400 ) | ( x99 & ~n7401 ) | ( n7400 & ~n7401 ) ;
  assign n7403 = n4334 & n5726 ;
  assign n7404 = n7402 | n7403 ;
  assign n7405 = n7404 ^ x8 ^ 1'b0 ;
  assign n7406 = n7405 ^ n7316 ^ n7145 ;
  assign n7407 = ( n7145 & n7316 ) | ( n7145 & n7405 ) | ( n7316 & n7405 ) ;
  assign n7408 = x98 & n6104 ;
  assign n7409 = ( x100 & n6105 ) | ( x100 & n7408 ) | ( n6105 & n7408 ) ;
  assign n7410 = n7408 | n7409 ;
  assign n7411 = x99 & ~n6107 ;
  assign n7412 = ( x99 & n7410 ) | ( x99 & ~n7411 ) | ( n7410 & ~n7411 ) ;
  assign n7413 = n4334 & ~n6108 ;
  assign n7414 = ( n4334 & n7412 ) | ( n4334 & ~n7413 ) | ( n7412 & ~n7413 ) ;
  assign n7415 = n7414 ^ x2 ^ 1'b0 ;
  assign n7416 = n7415 ^ n7366 ^ n7217 ;
  assign n7417 = ( n7217 & n7366 ) | ( n7217 & n7415 ) | ( n7366 & n7415 ) ;
  assign n7418 = x99 & n6104 ;
  assign n7419 = ( x101 & n6105 ) | ( x101 & n7418 ) | ( n6105 & n7418 ) ;
  assign n7420 = n7418 | n7419 ;
  assign n7421 = x100 & ~n6107 ;
  assign n7422 = ( x100 & n7420 ) | ( x100 & ~n7421 ) | ( n7420 & ~n7421 ) ;
  assign n7423 = n5687 & ~n6108 ;
  assign n7424 = ( n5687 & n7422 ) | ( n5687 & ~n7423 ) | ( n7422 & ~n7423 ) ;
  assign n7425 = n7424 ^ x2 ^ 1'b0 ;
  assign n7426 = n7425 ^ n7417 ^ n7226 ;
  assign n7427 = ( n7226 & n7417 ) | ( n7226 & n7425 ) | ( n7417 & n7425 ) ;
  assign n7428 = x96 & n5011 ;
  assign n7429 = ( x98 & n5012 ) | ( x98 & n7428 ) | ( n5012 & n7428 ) ;
  assign n7430 = n7428 | n7429 ;
  assign n7431 = x97 & ~n5008 ;
  assign n7432 = ( x97 & n7430 ) | ( x97 & ~n7431 ) | ( n7430 & ~n7431 ) ;
  assign n7433 = n4052 & n5020 ;
  assign n7434 = n7432 | n7433 ;
  assign n7435 = n7434 ^ x17 ^ 1'b0 ;
  assign n7436 = ( n6936 & n6977 ) | ( n6936 & n7435 ) | ( n6977 & n7435 ) ;
  assign n7437 = n7435 ^ n6977 ^ n6936 ;
  assign n7438 = x91 & n4616 ;
  assign n7439 = ( x93 & n4606 ) | ( x93 & n7438 ) | ( n4606 & n7438 ) ;
  assign n7440 = n7438 | n7439 ;
  assign n7441 = x92 & ~n4605 ;
  assign n7442 = ( x92 & n7440 ) | ( x92 & ~n7441 ) | ( n7440 & ~n7441 ) ;
  assign n7443 = n2476 & n4608 ;
  assign n7444 = n7442 | n7443 ;
  assign n7445 = n7444 ^ x23 ^ 1'b0 ;
  assign n7446 = n7445 ^ n6887 ^ n3995 ;
  assign n7447 = ( n3995 & n6887 ) | ( n3995 & n7445 ) | ( n6887 & n7445 ) ;
  assign n7448 = x94 & n4790 ;
  assign n7449 = ( x96 & n4792 ) | ( x96 & n7448 ) | ( n4792 & n7448 ) ;
  assign n7450 = n7448 | n7449 ;
  assign n7451 = x95 & ~n4786 ;
  assign n7452 = ( x95 & n7450 ) | ( x95 & ~n7451 ) | ( n7450 & ~n7451 ) ;
  assign n7453 = n2907 & n4787 ;
  assign n7454 = n7452 | n7453 ;
  assign n7455 = n7454 ^ x20 ^ 1'b0 ;
  assign n7456 = ( n6937 & n7446 ) | ( n6937 & n7455 ) | ( n7446 & n7455 ) ;
  assign n7457 = n197 & n1419 ;
  assign n7458 = n7455 ^ n7446 ^ n6937 ;
  assign n7459 = x97 & n5011 ;
  assign n7460 = ( x99 & n5012 ) | ( x99 & n7459 ) | ( n5012 & n7459 ) ;
  assign n7461 = n7459 | n7460 ;
  assign n7462 = x98 & ~n5008 ;
  assign n7463 = ( x98 & n7461 ) | ( x98 & ~n7462 ) | ( n7461 & ~n7462 ) ;
  assign n7464 = n4270 & n5020 ;
  assign n7465 = n7463 | n7464 ;
  assign n7466 = n7465 ^ x17 ^ 1'b0 ;
  assign n7467 = ( n7436 & n7458 ) | ( n7436 & n7466 ) | ( n7458 & n7466 ) ;
  assign n7468 = n7466 ^ n7458 ^ n7436 ;
  assign n7469 = x100 & n6104 ;
  assign n7470 = ( x102 & n6105 ) | ( x102 & n7469 ) | ( n6105 & n7469 ) ;
  assign n7471 = n7469 | n7470 ;
  assign n7472 = x101 & ~n6107 ;
  assign n7473 = ( x101 & n7471 ) | ( x101 & ~n7472 ) | ( n7471 & ~n7472 ) ;
  assign n7474 = n5947 & ~n6108 ;
  assign n7475 = ( n5947 & n7473 ) | ( n5947 & ~n7474 ) | ( n7473 & ~n7474 ) ;
  assign n7476 = n7475 ^ x2 ^ 1'b0 ;
  assign n7477 = n7476 ^ n7427 ^ n7266 ;
  assign n7478 = ( n7266 & n7427 ) | ( n7266 & n7476 ) | ( n7427 & n7476 ) ;
  assign n7479 = x97 & n5499 ;
  assign n7480 = ( x99 & n5497 ) | ( x99 & n7479 ) | ( n5497 & n7479 ) ;
  assign n7481 = n7479 | n7480 ;
  assign n7482 = x98 & ~n5502 ;
  assign n7483 = ( x98 & n7481 ) | ( x98 & ~n7482 ) | ( n7481 & ~n7482 ) ;
  assign n7484 = n4270 & n5501 ;
  assign n7485 = n7483 | n7484 ;
  assign n7486 = n7485 ^ x11 ^ 1'b0 ;
  assign n7487 = n7486 ^ n7296 ^ n7157 ;
  assign n7488 = ( n7157 & n7296 ) | ( n7157 & n7486 ) | ( n7296 & n7486 ) ;
  assign n7489 = x98 & n4972 ;
  assign n7490 = ( x100 & n4985 ) | ( x100 & n7489 ) | ( n4985 & n7489 ) ;
  assign n7491 = n7489 | n7490 ;
  assign n7492 = x99 & ~n4980 ;
  assign n7493 = ( x99 & n7491 ) | ( x99 & ~n7492 ) | ( n7491 & ~n7492 ) ;
  assign n7494 = n4334 & n4987 ;
  assign n7495 = n7493 | n7494 ;
  assign n7496 = n7495 ^ x14 ^ 1'b0 ;
  assign n7497 = n7496 ^ n7257 ^ n6976 ;
  assign n7498 = ( n6976 & n7257 ) | ( n6976 & n7496 ) | ( n7257 & n7496 ) ;
  assign n7499 = x98 & n5499 ;
  assign n7500 = ( x100 & n5497 ) | ( x100 & n7499 ) | ( n5497 & n7499 ) ;
  assign n7501 = n7499 | n7500 ;
  assign n7502 = x99 & ~n5502 ;
  assign n7503 = ( x99 & n7501 ) | ( x99 & ~n7502 ) | ( n7501 & ~n7502 ) ;
  assign n7504 = n4334 & n5501 ;
  assign n7505 = n7503 | n7504 ;
  assign n7506 = n7505 ^ x11 ^ 1'b0 ;
  assign n7507 = ( n7176 & n7488 ) | ( n7176 & n7506 ) | ( n7488 & n7506 ) ;
  assign n7508 = n7506 ^ n7488 ^ n7176 ;
  assign n7509 = x99 & n4972 ;
  assign n7510 = ( x101 & n4985 ) | ( x101 & n7509 ) | ( n4985 & n7509 ) ;
  assign n7511 = n7509 | n7510 ;
  assign n7512 = x100 & ~n4980 ;
  assign n7513 = ( x100 & n7511 ) | ( x100 & ~n7512 ) | ( n7511 & ~n7512 ) ;
  assign n7514 = n4987 & n5687 ;
  assign n7515 = n7513 | n7514 ;
  assign n7516 = n7515 ^ x14 ^ 1'b0 ;
  assign n7517 = ( n7437 & n7498 ) | ( n7437 & n7516 ) | ( n7498 & n7516 ) ;
  assign n7518 = n7516 ^ n7498 ^ n7437 ;
  assign n7519 = x99 & n5499 ;
  assign n7520 = ( x101 & n5497 ) | ( x101 & n7519 ) | ( n5497 & n7519 ) ;
  assign n7521 = n7519 | n7520 ;
  assign n7522 = x100 & ~n5502 ;
  assign n7523 = ( x100 & n7521 ) | ( x100 & ~n7522 ) | ( n7521 & ~n7522 ) ;
  assign n7524 = n5501 & n5687 ;
  assign n7525 = n7523 | n7524 ;
  assign n7526 = n7525 ^ x11 ^ 1'b0 ;
  assign n7527 = ( n7246 & n7507 ) | ( n7246 & n7526 ) | ( n7507 & n7526 ) ;
  assign n7528 = n7526 ^ n7507 ^ n7246 ;
  assign n7529 = x100 & n5499 ;
  assign n7530 = ( x102 & n5497 ) | ( x102 & n7529 ) | ( n5497 & n7529 ) ;
  assign n7531 = n7529 | n7530 ;
  assign n7532 = x101 & ~n5502 ;
  assign n7533 = ( x101 & n7531 ) | ( x101 & ~n7532 ) | ( n7531 & ~n7532 ) ;
  assign n7534 = n5501 & n5947 ;
  assign n7535 = n7533 | n7534 ;
  assign n7536 = n7535 ^ x11 ^ 1'b0 ;
  assign n7537 = n7536 ^ n7527 ^ n7256 ;
  assign n7538 = ( n7256 & n7527 ) | ( n7256 & n7536 ) | ( n7527 & n7536 ) ;
  assign n7539 = x99 & n5718 ;
  assign n7540 = ( x101 & n5720 ) | ( x101 & n7539 ) | ( n5720 & n7539 ) ;
  assign n7541 = n7539 | n7540 ;
  assign n7542 = x100 & ~n5727 ;
  assign n7543 = ( x100 & n7541 ) | ( x100 & ~n7542 ) | ( n7541 & ~n7542 ) ;
  assign n7544 = n5687 & n5726 ;
  assign n7545 = n7543 | n7544 ;
  assign n7546 = n7545 ^ x8 ^ 1'b0 ;
  assign n7547 = ( n7297 & n7407 ) | ( n7297 & n7546 ) | ( n7407 & n7546 ) ;
  assign n7548 = n7546 ^ n7407 ^ n7297 ;
  assign n7549 = x100 & n5718 ;
  assign n7550 = ( x102 & n5720 ) | ( x102 & n7549 ) | ( n5720 & n7549 ) ;
  assign n7551 = n7549 | n7550 ;
  assign n7552 = x101 & ~n5727 ;
  assign n7553 = ( x101 & n7551 ) | ( x101 & ~n7552 ) | ( n7551 & ~n7552 ) ;
  assign n7554 = n5726 & n5947 ;
  assign n7555 = n7553 | n7554 ;
  assign n7556 = n7555 ^ x8 ^ 1'b0 ;
  assign n7557 = ( n7487 & n7547 ) | ( n7487 & n7556 ) | ( n7547 & n7556 ) ;
  assign n7558 = n7556 ^ n7547 ^ n7487 ;
  assign n7559 = x92 & n4616 ;
  assign n7560 = ( x94 & n4606 ) | ( x94 & n7559 ) | ( n4606 & n7559 ) ;
  assign n7561 = n7559 | n7560 ;
  assign n7562 = x93 & ~n4605 ;
  assign n7563 = ( x93 & n7561 ) | ( x93 & ~n7562 ) | ( n7561 & ~n7562 ) ;
  assign n7564 = n2518 & n4608 ;
  assign n7565 = n7563 | n7564 ;
  assign n7566 = n7565 ^ x23 ^ 1'b0 ;
  assign n7567 = ( n4005 & n7447 ) | ( n4005 & n7566 ) | ( n7447 & n7566 ) ;
  assign n7568 = n7566 ^ n7447 ^ n4005 ;
  assign n7569 = x93 & n4616 ;
  assign n7570 = ( x95 & n4606 ) | ( x95 & n7569 ) | ( n4606 & n7569 ) ;
  assign n7571 = n7569 | n7570 ;
  assign n7572 = x94 & ~n4605 ;
  assign n7573 = ( x94 & n7571 ) | ( x94 & ~n7572 ) | ( n7571 & ~n7572 ) ;
  assign n7574 = n2854 & n4608 ;
  assign n7575 = n7573 | n7574 ;
  assign n7576 = n7575 ^ x23 ^ 1'b0 ;
  assign n7577 = n7576 ^ n7567 ^ n4016 ;
  assign n7578 = ( n4016 & n7567 ) | ( n4016 & n7576 ) | ( n7567 & n7576 ) ;
  assign n7579 = x94 & n4616 ;
  assign n7580 = ( x96 & n4606 ) | ( x96 & n7579 ) | ( n4606 & n7579 ) ;
  assign n7581 = n7579 | n7580 ;
  assign n7582 = x95 & ~n4605 ;
  assign n7583 = ( x95 & n7581 ) | ( x95 & ~n7582 ) | ( n7581 & ~n7582 ) ;
  assign n7584 = n2907 & n4608 ;
  assign n7585 = n7583 | n7584 ;
  assign n7586 = n7585 ^ x23 ^ 1'b0 ;
  assign n7587 = n7586 ^ n7578 ^ n4025 ;
  assign n7588 = ( n4025 & n7578 ) | ( n4025 & n7586 ) | ( n7578 & n7586 ) ;
  assign n7589 = x95 & n4616 ;
  assign n7590 = ( x97 & n4606 ) | ( x97 & n7589 ) | ( n4606 & n7589 ) ;
  assign n7591 = n7589 | n7590 ;
  assign n7592 = x96 & ~n4605 ;
  assign n7593 = ( x96 & n7591 ) | ( x96 & ~n7592 ) | ( n7591 & ~n7592 ) ;
  assign n7594 = n3668 & n4608 ;
  assign n7595 = n7593 | n7594 ;
  assign n7596 = n7595 ^ x23 ^ 1'b0 ;
  assign n7597 = n7596 ^ n7588 ^ n4036 ;
  assign n7598 = ( n4036 & n7588 ) | ( n4036 & n7596 ) | ( n7588 & n7596 ) ;
  assign n7599 = x96 & n4616 ;
  assign n7600 = ( x98 & n4606 ) | ( x98 & n7599 ) | ( n4606 & n7599 ) ;
  assign n7601 = n7599 | n7600 ;
  assign n7602 = x97 & ~n4605 ;
  assign n7603 = ( x97 & n7601 ) | ( x97 & ~n7602 ) | ( n7601 & ~n7602 ) ;
  assign n7604 = n4052 & n4608 ;
  assign n7605 = n7603 | n7604 ;
  assign n7606 = n7605 ^ x23 ^ 1'b0 ;
  assign n7607 = n7606 ^ n7598 ^ n4051 ;
  assign n7608 = ( n4051 & n7598 ) | ( n4051 & n7606 ) | ( n7598 & n7606 ) ;
  assign n7609 = x97 & n4616 ;
  assign n7610 = ( x99 & n4606 ) | ( x99 & n7609 ) | ( n4606 & n7609 ) ;
  assign n7611 = n7609 | n7610 ;
  assign n7612 = x98 & ~n4605 ;
  assign n7613 = ( x98 & n7611 ) | ( x98 & ~n7612 ) | ( n7611 & ~n7612 ) ;
  assign n7614 = n4270 & n4608 ;
  assign n7615 = n7613 | n7614 ;
  assign n7616 = n7615 ^ x23 ^ 1'b0 ;
  assign n7617 = n7616 ^ n7608 ^ n4066 ;
  assign n7618 = ( n4066 & n7608 ) | ( n4066 & n7616 ) | ( n7608 & n7616 ) ;
  assign n7619 = x95 & n4790 ;
  assign n7620 = ( x97 & n4792 ) | ( x97 & n7619 ) | ( n4792 & n7619 ) ;
  assign n7621 = n7619 | n7620 ;
  assign n7622 = x96 & ~n4786 ;
  assign n7623 = ( x96 & n7621 ) | ( x96 & ~n7622 ) | ( n7621 & ~n7622 ) ;
  assign n7624 = n3668 & n4787 ;
  assign n7625 = n7623 | n7624 ;
  assign n7626 = n7625 ^ x20 ^ 1'b0 ;
  assign n7627 = n7626 ^ n7568 ^ n7456 ;
  assign n7628 = ( n7456 & n7568 ) | ( n7456 & n7626 ) | ( n7568 & n7626 ) ;
  assign n7629 = x96 & n4790 ;
  assign n7630 = ( x98 & n4792 ) | ( x98 & n7629 ) | ( n4792 & n7629 ) ;
  assign n7631 = n7629 | n7630 ;
  assign n7632 = x97 & ~n4786 ;
  assign n7633 = ( x97 & n7631 ) | ( x97 & ~n7632 ) | ( n7631 & ~n7632 ) ;
  assign n7634 = n4052 & n4787 ;
  assign n7635 = n7633 | n7634 ;
  assign n7636 = n7635 ^ x20 ^ 1'b0 ;
  assign n7637 = ( n7577 & n7628 ) | ( n7577 & n7636 ) | ( n7628 & n7636 ) ;
  assign n7638 = n7636 ^ n7628 ^ n7577 ;
  assign n7639 = x97 & n4790 ;
  assign n7640 = ( x99 & n4792 ) | ( x99 & n7639 ) | ( n4792 & n7639 ) ;
  assign n7641 = n7639 | n7640 ;
  assign n7642 = x98 & ~n4786 ;
  assign n7643 = ( x98 & n7641 ) | ( x98 & ~n7642 ) | ( n7641 & ~n7642 ) ;
  assign n7644 = n4270 & n4787 ;
  assign n7645 = n7643 | n7644 ;
  assign n7646 = n7645 ^ x20 ^ 1'b0 ;
  assign n7647 = ( n7587 & n7637 ) | ( n7587 & n7646 ) | ( n7637 & n7646 ) ;
  assign n7648 = n7646 ^ n7637 ^ n7587 ;
  assign n7649 = x98 & n4790 ;
  assign n7650 = ( x100 & n4792 ) | ( x100 & n7649 ) | ( n4792 & n7649 ) ;
  assign n7651 = n7649 | n7650 ;
  assign n7652 = x99 & ~n4786 ;
  assign n7653 = ( x99 & n7651 ) | ( x99 & ~n7652 ) | ( n7651 & ~n7652 ) ;
  assign n7654 = n4334 & n4787 ;
  assign n7655 = n7653 | n7654 ;
  assign n7656 = n7655 ^ x20 ^ 1'b0 ;
  assign n7657 = ( n7597 & n7647 ) | ( n7597 & n7656 ) | ( n7647 & n7656 ) ;
  assign n7658 = n7656 ^ n7647 ^ n7597 ;
  assign n7659 = x99 & n4790 ;
  assign n7660 = ( x101 & n4792 ) | ( x101 & n7659 ) | ( n4792 & n7659 ) ;
  assign n7661 = n7659 | n7660 ;
  assign n7662 = x100 & ~n4786 ;
  assign n7663 = ( x100 & n7661 ) | ( x100 & ~n7662 ) | ( n7661 & ~n7662 ) ;
  assign n7664 = n4787 & n5687 ;
  assign n7665 = n7663 | n7664 ;
  assign n7666 = n7665 ^ x20 ^ 1'b0 ;
  assign n7667 = ( n7607 & n7657 ) | ( n7607 & n7666 ) | ( n7657 & n7666 ) ;
  assign n7668 = n7666 ^ n7657 ^ n7607 ;
  assign n7669 = x100 & n4790 ;
  assign n7670 = ( x102 & n4792 ) | ( x102 & n7669 ) | ( n4792 & n7669 ) ;
  assign n7671 = n7669 | n7670 ;
  assign n7672 = x101 & ~n4786 ;
  assign n7673 = ( x101 & n7671 ) | ( x101 & ~n7672 ) | ( n7671 & ~n7672 ) ;
  assign n7674 = n4787 & n5947 ;
  assign n7675 = n7673 | n7674 ;
  assign n7676 = n7675 ^ x20 ^ 1'b0 ;
  assign n7677 = ( n7617 & n7667 ) | ( n7617 & n7676 ) | ( n7667 & n7676 ) ;
  assign n7678 = n7676 ^ n7667 ^ n7617 ;
  assign n7679 = x84 & n208 ;
  assign n7680 = ( x86 & n194 ) | ( x86 & n7679 ) | ( n194 & n7679 ) ;
  assign n7681 = n7679 | n7680 ;
  assign n7682 = x85 & ~n192 ;
  assign n7683 = ( x85 & n7681 ) | ( x85 & ~n7682 ) | ( n7681 & ~n7682 ) ;
  assign n7684 = n7457 | n7683 ;
  assign n7685 = x99 & n3734 ;
  assign n7686 = ( x101 & n3732 ) | ( x101 & n7685 ) | ( n3732 & n7685 ) ;
  assign n7687 = n7685 | n7686 ;
  assign n7688 = x100 & ~n3737 ;
  assign n7689 = ( x100 & n7687 ) | ( x100 & ~n7688 ) | ( n7687 & ~n7688 ) ;
  assign n7690 = n3736 & n5687 ;
  assign n7691 = n7689 | n7690 ;
  assign n7692 = n7691 ^ x26 ^ 1'b0 ;
  assign n7693 = ( n4127 & n4349 ) | ( n4127 & n7692 ) | ( n4349 & n7692 ) ;
  assign n7694 = n7692 ^ n4349 ^ n4127 ;
  assign n7695 = x100 & n3734 ;
  assign n7696 = ( x102 & n3732 ) | ( x102 & n7695 ) | ( n3732 & n7695 ) ;
  assign n7697 = n7695 | n7696 ;
  assign n7698 = x101 & ~n3737 ;
  assign n7699 = ( x101 & n7697 ) | ( x101 & ~n7698 ) | ( n7697 & ~n7698 ) ;
  assign n7700 = n3736 & n5947 ;
  assign n7701 = n7699 | n7700 ;
  assign n7702 = n7701 ^ x26 ^ 1'b0 ;
  assign n7703 = n7702 ^ n7693 ^ n4308 ;
  assign n7704 = ( n4308 & n7693 ) | ( n4308 & n7702 ) | ( n7693 & n7702 ) ;
  assign n7705 = x98 & n5011 ;
  assign n7706 = ( x100 & n5012 ) | ( x100 & n7705 ) | ( n5012 & n7705 ) ;
  assign n7707 = n7705 | n7706 ;
  assign n7708 = x99 & ~n5008 ;
  assign n7709 = ( x99 & n7707 ) | ( x99 & ~n7708 ) | ( n7707 & ~n7708 ) ;
  assign n7710 = n4334 & n5020 ;
  assign n7711 = n7709 | n7710 ;
  assign n7712 = n7711 ^ x17 ^ 1'b0 ;
  assign n7713 = n7712 ^ n7627 ^ n7467 ;
  assign n7714 = ( n7467 & n7627 ) | ( n7467 & n7712 ) | ( n7627 & n7712 ) ;
  assign n7715 = x98 & n4616 ;
  assign n7716 = ( x100 & n4606 ) | ( x100 & n7715 ) | ( n4606 & n7715 ) ;
  assign n7717 = n7715 | n7716 ;
  assign n7718 = x99 & ~n4605 ;
  assign n7719 = ( x99 & n7717 ) | ( x99 & ~n7718 ) | ( n7717 & ~n7718 ) ;
  assign n7720 = n4334 & n4608 ;
  assign n7721 = n7719 | n7720 ;
  assign n7722 = n7721 ^ x23 ^ 1'b0 ;
  assign n7723 = ( n4076 & n7618 ) | ( n4076 & n7722 ) | ( n7618 & n7722 ) ;
  assign n7724 = n7722 ^ n7618 ^ n4076 ;
  assign n7725 = x99 & n5011 ;
  assign n7726 = ( x101 & n5012 ) | ( x101 & n7725 ) | ( n5012 & n7725 ) ;
  assign n7727 = n7725 | n7726 ;
  assign n7728 = x100 & ~n5008 ;
  assign n7729 = ( x100 & n7727 ) | ( x100 & ~n7728 ) | ( n7727 & ~n7728 ) ;
  assign n7730 = n5020 & n5687 ;
  assign n7731 = n7729 | n7730 ;
  assign n7732 = n7731 ^ x17 ^ 1'b0 ;
  assign n7733 = n7732 ^ n7714 ^ n7638 ;
  assign n7734 = ( n7638 & n7714 ) | ( n7638 & n7732 ) | ( n7714 & n7732 ) ;
  assign n7735 = x99 & n4616 ;
  assign n7736 = ( x101 & n4606 ) | ( x101 & n7735 ) | ( n4606 & n7735 ) ;
  assign n7737 = n7735 | n7736 ;
  assign n7738 = x100 & ~n4605 ;
  assign n7739 = ( x100 & n7737 ) | ( x100 & ~n7738 ) | ( n7737 & ~n7738 ) ;
  assign n7740 = n4608 & n5687 ;
  assign n7741 = n7739 | n7740 ;
  assign n7742 = n7741 ^ x23 ^ 1'b0 ;
  assign n7743 = ( n4087 & n7723 ) | ( n4087 & n7742 ) | ( n7723 & n7742 ) ;
  assign n7744 = n7742 ^ n7723 ^ n4087 ;
  assign n7745 = x100 & n4616 ;
  assign n7746 = ( x102 & n4606 ) | ( x102 & n7745 ) | ( n4606 & n7745 ) ;
  assign n7747 = n7745 | n7746 ;
  assign n7748 = x101 & ~n4605 ;
  assign n7749 = ( x101 & n7747 ) | ( x101 & ~n7748 ) | ( n7747 & ~n7748 ) ;
  assign n7750 = n4608 & n5947 ;
  assign n7751 = n7749 | n7750 ;
  assign n7752 = n7751 ^ x23 ^ 1'b0 ;
  assign n7753 = n7752 ^ n7743 ^ n4297 ;
  assign n7754 = ( n4297 & n7743 ) | ( n4297 & n7752 ) | ( n7743 & n7752 ) ;
  assign n7755 = x99 & n3344 ;
  assign n7756 = ( x101 & n3342 ) | ( x101 & n7755 ) | ( n3342 & n7755 ) ;
  assign n7757 = n7755 | n7756 ;
  assign n7758 = x100 & ~n3347 ;
  assign n7759 = ( x100 & n7757 ) | ( x100 & ~n7758 ) | ( n7757 & ~n7758 ) ;
  assign n7760 = n3346 & n5687 ;
  assign n7761 = n7759 | n7760 ;
  assign n7762 = n7761 ^ x29 ^ 1'b0 ;
  assign n7763 = ( n4108 & n4359 ) | ( n4108 & n7762 ) | ( n4359 & n7762 ) ;
  assign n7764 = n7762 ^ n4359 ^ n4108 ;
  assign n7765 = x100 & n2156 ;
  assign n7766 = ( x102 & n2163 ) | ( x102 & n7765 ) | ( n2163 & n7765 ) ;
  assign n7767 = n7765 | n7766 ;
  assign n7768 = x101 & ~n2158 ;
  assign n7769 = ( x101 & n7767 ) | ( x101 & ~n7768 ) | ( n7767 & ~n7768 ) ;
  assign n7770 = n2161 & n5947 ;
  assign n7771 = n7769 | n7770 ;
  assign n7772 = n7771 ^ x38 ^ 1'b0 ;
  assign n7773 = n7772 ^ n4471 ^ n4097 ;
  assign n7774 = ( n4097 & n4471 ) | ( n4097 & n7772 ) | ( n4471 & n7772 ) ;
  assign n7775 = x100 & n2560 ;
  assign n7776 = ( x102 & n2567 ) | ( x102 & n7775 ) | ( n2567 & n7775 ) ;
  assign n7777 = n7775 | n7776 ;
  assign n7778 = x101 & ~n2562 ;
  assign n7779 = ( x101 & n7777 ) | ( x101 & ~n7778 ) | ( n7777 & ~n7778 ) ;
  assign n7780 = n2565 & n5947 ;
  assign n7781 = n7779 | n7780 ;
  assign n7782 = n7781 ^ x35 ^ 1'b0 ;
  assign n7783 = n7782 ^ n4318 ^ n4118 ;
  assign n7784 = ( n4118 & n4318 ) | ( n4118 & n7782 ) | ( n4318 & n7782 ) ;
  assign n7785 = x100 & n5011 ;
  assign n7786 = ( x102 & n5012 ) | ( x102 & n7785 ) | ( n5012 & n7785 ) ;
  assign n7787 = n7785 | n7786 ;
  assign n7788 = x101 & ~n5008 ;
  assign n7789 = ( x101 & n7787 ) | ( x101 & ~n7788 ) | ( n7787 & ~n7788 ) ;
  assign n7790 = n5020 & n5947 ;
  assign n7791 = n7789 | n7790 ;
  assign n7792 = n7791 ^ x17 ^ 1'b0 ;
  assign n7793 = n7792 ^ n7734 ^ n7648 ;
  assign n7794 = ( n7648 & n7734 ) | ( n7648 & n7792 ) | ( n7734 & n7792 ) ;
  assign n7795 = x100 & n3344 ;
  assign n7796 = ( x102 & n3342 ) | ( x102 & n7795 ) | ( n3342 & n7795 ) ;
  assign n7797 = n7795 | n7796 ;
  assign n7798 = x101 & ~n3347 ;
  assign n7799 = ( x101 & n7797 ) | ( x101 & ~n7798 ) | ( n7797 & ~n7798 ) ;
  assign n7800 = n3346 & n5947 ;
  assign n7801 = n7799 | n7800 ;
  assign n7802 = n7801 ^ x29 ^ 1'b0 ;
  assign n7803 = ( n4276 & n7763 ) | ( n4276 & n7802 ) | ( n7763 & n7802 ) ;
  assign n7804 = n7802 ^ n7763 ^ n4276 ;
  assign n7805 = x99 & n2156 ;
  assign n7806 = ( x101 & n2163 ) | ( x101 & n7805 ) | ( n2163 & n7805 ) ;
  assign n7807 = n7805 | n7806 ;
  assign n7808 = x100 & ~n2158 ;
  assign n7809 = ( x100 & n7807 ) | ( x100 & ~n7808 ) | ( n7807 & ~n7808 ) ;
  assign n7810 = n2161 & n5687 ;
  assign n7811 = n7809 | n7810 ;
  assign n7812 = n7811 ^ x38 ^ 1'b0 ;
  assign n7813 = ( n3708 & n4098 ) | ( n3708 & n7812 ) | ( n4098 & n7812 ) ;
  assign n7814 = n7812 ^ n4098 ^ n3708 ;
  assign n7815 = x100 & n3025 ;
  assign n7816 = ( x102 & n3015 ) | ( x102 & n7815 ) | ( n3015 & n7815 ) ;
  assign n7817 = n7815 | n7816 ;
  assign n7818 = x101 & ~n3014 ;
  assign n7819 = ( x101 & n7817 ) | ( x101 & ~n7818 ) | ( n7817 & ~n7818 ) ;
  assign n7820 = ( n3017 & n5947 ) | ( n3017 & n7819 ) | ( n5947 & n7819 ) ;
  assign n7821 = n7819 | n7820 ;
  assign n7822 = n7821 ^ x32 ^ 1'b0 ;
  assign n7823 = n7822 ^ n4288 ^ n4138 ;
  assign n7824 = ( n4138 & n4288 ) | ( n4138 & n7822 ) | ( n4288 & n7822 ) ;
  assign n7825 = x100 & n4972 ;
  assign n7826 = ( x102 & n4985 ) | ( x102 & n7825 ) | ( n4985 & n7825 ) ;
  assign n7827 = n7825 | n7826 ;
  assign n7828 = x101 & ~n4980 ;
  assign n7829 = ( x101 & n7827 ) | ( x101 & ~n7828 ) | ( n7827 & ~n7828 ) ;
  assign n7830 = n4987 & n5947 ;
  assign n7831 = n7829 | n7830 ;
  assign n7832 = n7831 ^ x14 ^ 1'b0 ;
  assign n7833 = n7832 ^ n7517 ^ n7468 ;
  assign n7834 = ( n7468 & n7517 ) | ( n7468 & n7832 ) | ( n7517 & n7832 ) ;
  assign n7835 = x99 & n3025 ;
  assign n7836 = ( x101 & n3015 ) | ( x101 & n7835 ) | ( n3015 & n7835 ) ;
  assign n7837 = n7835 | n7836 ;
  assign n7838 = x100 & ~n3014 ;
  assign n7839 = ( x100 & n7837 ) | ( x100 & ~n7838 ) | ( n7837 & ~n7838 ) ;
  assign n7840 = ( n3017 & n5687 ) | ( n3017 & n7839 ) | ( n5687 & n7839 ) ;
  assign n7841 = n7839 | n7840 ;
  assign n7842 = n7841 ^ x32 ^ 1'b0 ;
  assign n7843 = ( n3697 & n4137 ) | ( n3697 & n7842 ) | ( n4137 & n7842 ) ;
  assign n7844 = n7842 ^ n4137 ^ n3697 ;
  assign n7845 = x99 & n2560 ;
  assign n7846 = ( x101 & n2567 ) | ( x101 & n7845 ) | ( n2567 & n7845 ) ;
  assign n7847 = n7845 | n7846 ;
  assign n7848 = x100 & ~n2562 ;
  assign n7849 = ( x100 & n7847 ) | ( x100 & ~n7848 ) | ( n7847 & ~n7848 ) ;
  assign n7850 = n2565 & n5687 ;
  assign n7851 = n7849 | n7850 ;
  assign n7852 = n7851 ^ x35 ^ 1'b0 ;
  assign n7853 = ( n3728 & n4117 ) | ( n3728 & n7852 ) | ( n4117 & n7852 ) ;
  assign n7854 = n7852 ^ n4117 ^ n3728 ;
  assign n7855 = x101 & n2560 ;
  assign n7856 = ( x103 & n2567 ) | ( x103 & n7855 ) | ( n2567 & n7855 ) ;
  assign n7857 = n7855 | n7856 ;
  assign n7858 = x102 & ~n2562 ;
  assign n7859 = ( x102 & n7857 ) | ( x102 & ~n7858 ) | ( n7857 & ~n7858 ) ;
  assign n7860 = n5952 ^ x103 ^ x102 ;
  assign n7861 = n2565 & n7860 ;
  assign n7862 = n7859 | n7861 ;
  assign n7863 = n7862 ^ x35 ^ 1'b0 ;
  assign n7864 = n7863 ^ n7784 ^ n4338 ;
  assign n7865 = ( n4338 & n7784 ) | ( n4338 & n7863 ) | ( n7784 & n7863 ) ;
  assign n7866 = x101 & n888 ;
  assign n7867 = ( x103 & n878 ) | ( x103 & n7866 ) | ( n878 & n7866 ) ;
  assign n7868 = n7866 | n7867 ;
  assign n7869 = x102 & ~n877 ;
  assign n7870 = ( x102 & n7868 ) | ( x102 & ~n7869 ) | ( n7868 & ~n7869 ) ;
  assign n7871 = n880 & n7860 ;
  assign n7872 = n7870 | n7871 ;
  assign n7873 = n7872 ^ x44 ^ 1'b0 ;
  assign n7874 = n7684 ^ x62 ^ 1'b0 ;
  assign n7875 = ( n4600 & n5962 ) | ( n4600 & ~n7873 ) | ( n5962 & ~n7873 ) ;
  assign n7876 = n7873 ^ n5962 ^ n4600 ;
  assign n7877 = x101 & n1058 ;
  assign n7878 = ( x103 & n1065 ) | ( x103 & n7877 ) | ( n1065 & n7877 ) ;
  assign n7879 = n7877 | n7878 ;
  assign n7880 = x102 & ~n1060 ;
  assign n7881 = ( x102 & n7879 ) | ( x102 & ~n7880 ) | ( n7879 & ~n7880 ) ;
  assign n7882 = n1063 & n7860 ;
  assign n7883 = n7881 | n7882 ;
  assign n7884 = n7883 ^ x41 ^ 1'b0 ;
  assign n7885 = n7884 ^ n5951 ^ n4368 ;
  assign n7886 = ( n4368 & n5951 ) | ( n4368 & n7884 ) | ( n5951 & n7884 ) ;
  assign n7887 = x101 & n2156 ;
  assign n7888 = ( x103 & n2163 ) | ( x103 & n7887 ) | ( n2163 & n7887 ) ;
  assign n7889 = n7887 | n7888 ;
  assign n7890 = x102 & ~n2158 ;
  assign n7891 = ( x102 & n7889 ) | ( x102 & ~n7890 ) | ( n7889 & ~n7890 ) ;
  assign n7892 = n2161 & n7860 ;
  assign n7893 = n7891 | n7892 ;
  assign n7894 = n7893 ^ x38 ^ 1'b0 ;
  assign n7895 = ( n4480 & n7774 ) | ( n4480 & n7894 ) | ( n7774 & n7894 ) ;
  assign n7896 = n7894 ^ n7774 ^ n4480 ;
  assign n7897 = x101 & n5979 ;
  assign n7898 = ( x103 & n5969 ) | ( x103 & n7897 ) | ( n5969 & n7897 ) ;
  assign n7899 = n7897 | n7898 ;
  assign n7900 = x102 & ~n5970 ;
  assign n7901 = ( x102 & n7899 ) | ( x102 & ~n7900 ) | ( n7899 & ~n7900 ) ;
  assign n7902 = n5968 & n7860 ;
  assign n7903 = n7901 | n7902 ;
  assign n7904 = n7903 ^ x5 ^ 1'b0 ;
  assign n7905 = n7904 ^ n7406 ^ n7397 ;
  assign n7906 = ( n7397 & n7406 ) | ( n7397 & n7904 ) | ( n7406 & n7904 ) ;
  assign n7907 = x101 & n5011 ;
  assign n7908 = ( x103 & n5012 ) | ( x103 & n7907 ) | ( n5012 & n7907 ) ;
  assign n7909 = n7907 | n7908 ;
  assign n7910 = x102 & ~n5008 ;
  assign n7911 = ( x102 & n7909 ) | ( x102 & ~n7910 ) | ( n7909 & ~n7910 ) ;
  assign n7912 = n5020 & n7860 ;
  assign n7913 = n7911 | n7912 ;
  assign n7914 = n7913 ^ x17 ^ 1'b0 ;
  assign n7915 = ( n7658 & n7794 ) | ( n7658 & n7914 ) | ( n7794 & n7914 ) ;
  assign n7916 = n7914 ^ n7794 ^ n7658 ;
  assign n7917 = x101 & n3344 ;
  assign n7918 = ( x103 & n3342 ) | ( x103 & n7917 ) | ( n3342 & n7917 ) ;
  assign n7919 = n7917 | n7918 ;
  assign n7920 = x102 & ~n3347 ;
  assign n7921 = ( x102 & n7919 ) | ( x102 & ~n7920 ) | ( n7919 & ~n7920 ) ;
  assign n7922 = ( n3346 & n7860 ) | ( n3346 & n7921 ) | ( n7860 & n7921 ) ;
  assign n7923 = n7921 | n7922 ;
  assign n7924 = n7923 ^ x29 ^ 1'b0 ;
  assign n7925 = ( n4277 & n4389 ) | ( n4277 & n7924 ) | ( n4389 & n7924 ) ;
  assign n7926 = n7924 ^ n4389 ^ n4277 ;
  assign n7927 = x101 & n5718 ;
  assign n7928 = ( x103 & n5720 ) | ( x103 & n7927 ) | ( n5720 & n7927 ) ;
  assign n7929 = n7927 | n7928 ;
  assign n7930 = x102 & ~n5727 ;
  assign n7931 = ( x102 & n7929 ) | ( x102 & ~n7930 ) | ( n7929 & ~n7930 ) ;
  assign n7932 = n5726 & n7860 ;
  assign n7933 = n7931 | n7932 ;
  assign n7934 = n7933 ^ x8 ^ 1'b0 ;
  assign n7935 = ( n7508 & n7557 ) | ( n7508 & n7934 ) | ( n7557 & n7934 ) ;
  assign n7936 = n7934 ^ n7557 ^ n7508 ;
  assign n7937 = x101 & n3025 ;
  assign n7938 = ( x103 & n3015 ) | ( x103 & n7937 ) | ( n3015 & n7937 ) ;
  assign n7939 = n7937 | n7938 ;
  assign n7940 = x102 & ~n3014 ;
  assign n7941 = ( x102 & n7939 ) | ( x102 & ~n7940 ) | ( n7939 & ~n7940 ) ;
  assign n7942 = n3017 & n7860 ;
  assign n7943 = n7941 | n7942 ;
  assign n7944 = n7943 ^ x32 ^ 1'b0 ;
  assign n7945 = ( n4378 & n7824 ) | ( n4378 & n7944 ) | ( n7824 & n7944 ) ;
  assign n7946 = n7944 ^ n7824 ^ n4378 ;
  assign n7947 = x101 & n3734 ;
  assign n7948 = ( x103 & n3732 ) | ( x103 & n7947 ) | ( n3732 & n7947 ) ;
  assign n7949 = n7947 | n7948 ;
  assign n7950 = x102 & ~n3737 ;
  assign n7951 = ( x102 & n7949 ) | ( x102 & ~n7950 ) | ( n7949 & ~n7950 ) ;
  assign n7952 = n3736 & n7860 ;
  assign n7953 = n7951 | n7952 ;
  assign n7954 = n7953 ^ x26 ^ 1'b0 ;
  assign n7955 = n7954 ^ n7704 ^ n4358 ;
  assign n7956 = ( n4358 & n7704 ) | ( n4358 & n7954 ) | ( n7704 & n7954 ) ;
  assign n7957 = x101 & n5499 ;
  assign n7958 = ( x103 & n5497 ) | ( x103 & n7957 ) | ( n5497 & n7957 ) ;
  assign n7959 = n7957 | n7958 ;
  assign n7960 = x102 & ~n5502 ;
  assign n7961 = ( x102 & n7959 ) | ( x102 & ~n7960 ) | ( n7959 & ~n7960 ) ;
  assign n7962 = n5501 & n7860 ;
  assign n7963 = n7961 | n7962 ;
  assign n7964 = n7963 ^ x11 ^ 1'b0 ;
  assign n7965 = n7964 ^ n7538 ^ n7497 ;
  assign n7966 = ( n7497 & n7538 ) | ( n7497 & n7964 ) | ( n7538 & n7964 ) ;
  assign n7967 = x101 & n4616 ;
  assign n7968 = ( x103 & n4606 ) | ( x103 & n7967 ) | ( n4606 & n7967 ) ;
  assign n7969 = n7967 | n7968 ;
  assign n7970 = x102 & ~n4605 ;
  assign n7971 = ( x102 & n7969 ) | ( x102 & ~n7970 ) | ( n7969 & ~n7970 ) ;
  assign n7972 = n4608 & n7860 ;
  assign n7973 = n7971 | n7972 ;
  assign n7974 = n7973 ^ x23 ^ 1'b0 ;
  assign n7975 = n7974 ^ n7754 ^ n4348 ;
  assign n7976 = ( n4348 & n7754 ) | ( n4348 & n7974 ) | ( n7754 & n7974 ) ;
  assign n7977 = x101 & n4972 ;
  assign n7978 = ( x102 & x103 ) | ( x102 & n5952 ) | ( x103 & n5952 ) ;
  assign n7979 = ( x103 & n4985 ) | ( x103 & n7977 ) | ( n4985 & n7977 ) ;
  assign n7980 = n7977 | n7979 ;
  assign n7981 = x102 & ~n4980 ;
  assign n7982 = ( x102 & n7980 ) | ( x102 & ~n7981 ) | ( n7980 & ~n7981 ) ;
  assign n7983 = n4987 & n7860 ;
  assign n7984 = n7982 | n7983 ;
  assign n7985 = n7984 ^ x14 ^ 1'b0 ;
  assign n7986 = ( n7713 & n7834 ) | ( n7713 & n7985 ) | ( n7834 & n7985 ) ;
  assign n7987 = n7985 ^ n7834 ^ n7713 ;
  assign n7988 = x101 & n4790 ;
  assign n7989 = ( x103 & n4792 ) | ( x103 & n7988 ) | ( n4792 & n7988 ) ;
  assign n7990 = n7988 | n7989 ;
  assign n7991 = x102 & ~n4786 ;
  assign n7992 = ( x102 & n7990 ) | ( x102 & ~n7991 ) | ( n7990 & ~n7991 ) ;
  assign n7993 = n4787 & n7860 ;
  assign n7994 = n7992 | n7993 ;
  assign n7995 = n7994 ^ x20 ^ 1'b0 ;
  assign n7996 = ( n7677 & n7724 ) | ( n7677 & n7995 ) | ( n7724 & n7995 ) ;
  assign n7997 = n7995 ^ n7724 ^ n7677 ;
  assign n7998 = x101 & n6104 ;
  assign n7999 = ( x103 & n6105 ) | ( x103 & n7998 ) | ( n6105 & n7998 ) ;
  assign n8000 = n7998 | n7999 ;
  assign n8001 = x102 & ~n6107 ;
  assign n8002 = ( x102 & n8000 ) | ( x102 & ~n8001 ) | ( n8000 & ~n8001 ) ;
  assign n8003 = ~n6108 & n7860 ;
  assign n8004 = ( n7860 & n8002 ) | ( n7860 & ~n8003 ) | ( n8002 & ~n8003 ) ;
  assign n8005 = n8004 ^ x2 ^ 1'b0 ;
  assign n8006 = n8005 ^ n7478 ^ n7377 ;
  assign n8007 = ( n7377 & n7478 ) | ( n7377 & n8005 ) | ( n7478 & n8005 ) ;
  assign n8008 = x103 & ~n5008 ;
  assign n8009 = x102 & n5011 ;
  assign n8010 = ( x104 & n5012 ) | ( x104 & n8009 ) | ( n5012 & n8009 ) ;
  assign n8011 = n8009 | n8010 ;
  assign n8012 = n7978 ^ x104 ^ x103 ;
  assign n8013 = ( x103 & ~n8008 ) | ( x103 & n8011 ) | ( ~n8008 & n8011 ) ;
  assign n8014 = n5020 & n8012 ;
  assign n8015 = n8013 | n8014 ;
  assign n8016 = n8015 ^ x17 ^ 1'b0 ;
  assign n8017 = n8016 ^ n7915 ^ n7668 ;
  assign n8018 = ( n7668 & n7915 ) | ( n7668 & n8016 ) | ( n7915 & n8016 ) ;
  assign n8019 = x102 & n4616 ;
  assign n8020 = ( x104 & n4606 ) | ( x104 & n8019 ) | ( n4606 & n8019 ) ;
  assign n8021 = n8019 | n8020 ;
  assign n8022 = x103 & ~n4605 ;
  assign n8023 = ( x103 & n8021 ) | ( x103 & ~n8022 ) | ( n8021 & ~n8022 ) ;
  assign n8024 = n4608 & n8012 ;
  assign n8025 = n8023 | n8024 ;
  assign n8026 = n8025 ^ x23 ^ 1'b0 ;
  assign n8027 = n8026 ^ n7976 ^ n7694 ;
  assign n8028 = ( n7694 & n7976 ) | ( n7694 & n8026 ) | ( n7976 & n8026 ) ;
  assign n8029 = x102 & n3344 ;
  assign n8030 = ( x104 & n3342 ) | ( x104 & n8029 ) | ( n3342 & n8029 ) ;
  assign n8031 = n8029 | n8030 ;
  assign n8032 = x103 & ~n3347 ;
  assign n8033 = ( x103 & n8031 ) | ( x103 & ~n8032 ) | ( n8031 & ~n8032 ) ;
  assign n8034 = ( n3346 & n8012 ) | ( n3346 & n8033 ) | ( n8012 & n8033 ) ;
  assign n8035 = n8033 | n8034 ;
  assign n8036 = n8035 ^ x29 ^ 1'b0 ;
  assign n8037 = ( n4388 & n7844 ) | ( n4388 & n8036 ) | ( n7844 & n8036 ) ;
  assign n8038 = n8036 ^ n7844 ^ n4388 ;
  assign n8039 = x102 & n6104 ;
  assign n8040 = ( x104 & n6105 ) | ( x104 & n8039 ) | ( n6105 & n8039 ) ;
  assign n8041 = ( x103 & x104 ) | ( x103 & n7978 ) | ( x104 & n7978 ) ;
  assign n8042 = n8039 | n8040 ;
  assign n8043 = x103 & ~n6107 ;
  assign n8044 = ( x103 & n8042 ) | ( x103 & ~n8043 ) | ( n8042 & ~n8043 ) ;
  assign n8045 = ~n6108 & n8012 ;
  assign n8046 = ( n8012 & n8044 ) | ( n8012 & ~n8045 ) | ( n8044 & ~n8045 ) ;
  assign n8047 = n8046 ^ x2 ^ 1'b0 ;
  assign n8048 = ( n7386 & n8007 ) | ( n7386 & n8047 ) | ( n8007 & n8047 ) ;
  assign n8049 = n8047 ^ n8007 ^ n7386 ;
  assign n8050 = x102 & n2156 ;
  assign n8051 = ( x104 & n2163 ) | ( x104 & n8050 ) | ( n2163 & n8050 ) ;
  assign n8052 = n8050 | n8051 ;
  assign n8053 = x103 & ~n2158 ;
  assign n8054 = ( x103 & n8052 ) | ( x103 & ~n8053 ) | ( n8052 & ~n8053 ) ;
  assign n8055 = n2161 & n8012 ;
  assign n8056 = n8054 | n8055 ;
  assign n8057 = n8056 ^ x38 ^ 1'b0 ;
  assign n8058 = ( n4481 & n5691 ) | ( n4481 & n8057 ) | ( n5691 & n8057 ) ;
  assign n8059 = n8057 ^ n5691 ^ n4481 ;
  assign n8060 = x102 & n5718 ;
  assign n8061 = ( x104 & n5720 ) | ( x104 & n8060 ) | ( n5720 & n8060 ) ;
  assign n8062 = n8060 | n8061 ;
  assign n8063 = x103 & ~n5727 ;
  assign n8064 = ( x103 & n8062 ) | ( x103 & ~n8063 ) | ( n8062 & ~n8063 ) ;
  assign n8065 = n5726 & n8012 ;
  assign n8066 = n8064 | n8065 ;
  assign n8067 = n8066 ^ x8 ^ 1'b0 ;
  assign n8068 = ( n7528 & n7935 ) | ( n7528 & n8067 ) | ( n7935 & n8067 ) ;
  assign n8069 = n8067 ^ n7935 ^ n7528 ;
  assign n8070 = x102 & n3734 ;
  assign n8071 = ( x104 & n3732 ) | ( x104 & n8070 ) | ( n3732 & n8070 ) ;
  assign n8072 = n8070 | n8071 ;
  assign n8073 = x103 & ~n3737 ;
  assign n8074 = ( x103 & n8072 ) | ( x103 & ~n8073 ) | ( n8072 & ~n8073 ) ;
  assign n8075 = n3736 & n8012 ;
  assign n8076 = n8074 | n8075 ;
  assign n8077 = n8076 ^ x26 ^ 1'b0 ;
  assign n8078 = n8077 ^ n7956 ^ n7764 ;
  assign n8079 = ( n7764 & n7956 ) | ( n7764 & n8077 ) | ( n7956 & n8077 ) ;
  assign n8080 = x102 & n5979 ;
  assign n8081 = ( x104 & n5969 ) | ( x104 & n8080 ) | ( n5969 & n8080 ) ;
  assign n8082 = n8080 | n8081 ;
  assign n8083 = x103 & ~n5970 ;
  assign n8084 = ( x103 & n8082 ) | ( x103 & ~n8083 ) | ( n8082 & ~n8083 ) ;
  assign n8085 = n5968 & n8012 ;
  assign n8086 = n8084 | n8085 ;
  assign n8087 = n8086 ^ x5 ^ 1'b0 ;
  assign n8088 = n8087 ^ n7906 ^ n7548 ;
  assign n8089 = ( n7548 & n7906 ) | ( n7548 & n8087 ) | ( n7906 & n8087 ) ;
  assign n8090 = x102 & n4972 ;
  assign n8091 = ( x104 & n4985 ) | ( x104 & n8090 ) | ( n4985 & n8090 ) ;
  assign n8092 = n8090 | n8091 ;
  assign n8093 = x103 & ~n4980 ;
  assign n8094 = ( x103 & n8092 ) | ( x103 & ~n8093 ) | ( n8092 & ~n8093 ) ;
  assign n8095 = n4987 & n8012 ;
  assign n8096 = n8094 | n8095 ;
  assign n8097 = n8096 ^ x14 ^ 1'b0 ;
  assign n8098 = n8097 ^ n7986 ^ n7733 ;
  assign n8099 = ( n7733 & n7986 ) | ( n7733 & n8097 ) | ( n7986 & n8097 ) ;
  assign n8100 = x103 & n1058 ;
  assign n8101 = ( x105 & n1065 ) | ( x105 & n8100 ) | ( n1065 & n8100 ) ;
  assign n8102 = n8100 | n8101 ;
  assign n8103 = x104 & ~n1060 ;
  assign n8104 = ( x104 & n8102 ) | ( x104 & ~n8103 ) | ( n8102 & ~n8103 ) ;
  assign n8105 = n8041 ^ x105 ^ x104 ;
  assign n8106 = n1063 & n8105 ;
  assign n8107 = n8104 | n8106 ;
  assign n8108 = n8107 ^ x41 ^ 1'b0 ;
  assign n8109 = ( n5712 & n5963 ) | ( n5712 & n8108 ) | ( n5963 & n8108 ) ;
  assign n8110 = n8108 ^ n5963 ^ n5712 ;
  assign n8111 = x103 & n6104 ;
  assign n8112 = ( x105 & n6105 ) | ( x105 & n8111 ) | ( n6105 & n8111 ) ;
  assign n8113 = n8111 | n8112 ;
  assign n8114 = x104 & ~n6107 ;
  assign n8115 = ( x104 & n8113 ) | ( x104 & ~n8114 ) | ( n8113 & ~n8114 ) ;
  assign n8116 = ~n6108 & n8105 ;
  assign n8117 = ( n8105 & n8115 ) | ( n8105 & ~n8116 ) | ( n8115 & ~n8116 ) ;
  assign n8118 = n8117 ^ x2 ^ 1'b0 ;
  assign n8119 = ( n7396 & n8048 ) | ( n7396 & n8118 ) | ( n8048 & n8118 ) ;
  assign n8120 = n8118 ^ n8048 ^ n7396 ;
  assign n8121 = x103 & n4616 ;
  assign n8122 = ( x105 & n4606 ) | ( x105 & n8121 ) | ( n4606 & n8121 ) ;
  assign n8123 = n8121 | n8122 ;
  assign n8124 = x104 & ~n4605 ;
  assign n8125 = ( x104 & n8123 ) | ( x104 & ~n8124 ) | ( n8123 & ~n8124 ) ;
  assign n8126 = n4608 & n8105 ;
  assign n8127 = n8125 | n8126 ;
  assign n8128 = n8127 ^ x23 ^ 1'b0 ;
  assign n8129 = ( n7703 & n8028 ) | ( n7703 & n8128 ) | ( n8028 & n8128 ) ;
  assign n8130 = n8128 ^ n8028 ^ n7703 ;
  assign n8131 = x103 & n5979 ;
  assign n8132 = ( x105 & n5969 ) | ( x105 & n8131 ) | ( n5969 & n8131 ) ;
  assign n8133 = n8131 | n8132 ;
  assign n8134 = x104 & ~n5970 ;
  assign n8135 = ( x104 & n8133 ) | ( x104 & ~n8134 ) | ( n8133 & ~n8134 ) ;
  assign n8136 = n5968 & n8105 ;
  assign n8137 = n8135 | n8136 ;
  assign n8138 = n8137 ^ x5 ^ 1'b0 ;
  assign n8139 = n8138 ^ n8089 ^ n7558 ;
  assign n8140 = ( n7558 & n8089 ) | ( n7558 & n8138 ) | ( n8089 & n8138 ) ;
  assign n8141 = x103 & n3025 ;
  assign n8142 = ( x105 & n3015 ) | ( x105 & n8141 ) | ( n3015 & n8141 ) ;
  assign n8143 = ( x104 & x105 ) | ( x104 & n8041 ) | ( x105 & n8041 ) ;
  assign n8144 = n8141 | n8142 ;
  assign n8145 = x104 & ~n3014 ;
  assign n8146 = ( x104 & n8144 ) | ( x104 & ~n8145 ) | ( n8144 & ~n8145 ) ;
  assign n8147 = n3017 & n8105 ;
  assign n8148 = n8146 | n8147 ;
  assign n8149 = n8148 ^ x32 ^ 1'b0 ;
  assign n8150 = n8149 ^ n7853 ^ n7783 ;
  assign n8151 = ( n7783 & n7853 ) | ( n7783 & n8149 ) | ( n7853 & n8149 ) ;
  assign n8152 = x103 & n2560 ;
  assign n8153 = ( x105 & n2567 ) | ( x105 & n8152 ) | ( n2567 & n8152 ) ;
  assign n8154 = n8152 | n8153 ;
  assign n8155 = x104 & ~n2562 ;
  assign n8156 = ( x104 & n8154 ) | ( x104 & ~n8155 ) | ( n8154 & ~n8155 ) ;
  assign n8157 = n2565 & n8105 ;
  assign n8158 = n8156 | n8157 ;
  assign n8159 = n8158 ^ x35 ^ 1'b0 ;
  assign n8160 = ( n7773 & n7813 ) | ( n7773 & n8159 ) | ( n7813 & n8159 ) ;
  assign n8161 = n8159 ^ n7813 ^ n7773 ;
  assign n8162 = x103 & n5011 ;
  assign n8163 = ( x105 & n5012 ) | ( x105 & n8162 ) | ( n5012 & n8162 ) ;
  assign n8164 = n8162 | n8163 ;
  assign n8165 = x104 & ~n5008 ;
  assign n8166 = ( x104 & n8164 ) | ( x104 & ~n8165 ) | ( n8164 & ~n8165 ) ;
  assign n8167 = n5020 & n8105 ;
  assign n8168 = n8166 | n8167 ;
  assign n8169 = n8168 ^ x17 ^ 1'b0 ;
  assign n8170 = ( n7678 & n8018 ) | ( n7678 & n8169 ) | ( n8018 & n8169 ) ;
  assign n8171 = n8169 ^ n8018 ^ n7678 ;
  assign n8172 = x103 & n3344 ;
  assign n8173 = ( x105 & n3342 ) | ( x105 & n8172 ) | ( n3342 & n8172 ) ;
  assign n8174 = n8172 | n8173 ;
  assign n8175 = x104 & ~n3347 ;
  assign n8176 = ( x104 & n8174 ) | ( x104 & ~n8175 ) | ( n8174 & ~n8175 ) ;
  assign n8177 = n3346 & n8105 ;
  assign n8178 = n8176 | n8177 ;
  assign n8179 = n8178 ^ x29 ^ 1'b0 ;
  assign n8180 = n8179 ^ n7843 ^ n7823 ;
  assign n8181 = ( n7823 & n7843 ) | ( n7823 & n8179 ) | ( n7843 & n8179 ) ;
  assign n8182 = x103 & n5718 ;
  assign n8183 = ( x105 & n5720 ) | ( x105 & n8182 ) | ( n5720 & n8182 ) ;
  assign n8184 = n8182 | n8183 ;
  assign n8185 = x104 & ~n5727 ;
  assign n8186 = ( x104 & n8184 ) | ( x104 & ~n8185 ) | ( n8184 & ~n8185 ) ;
  assign n8187 = n5726 & n8105 ;
  assign n8188 = n8186 | n8187 ;
  assign n8189 = n8188 ^ x8 ^ 1'b0 ;
  assign n8190 = n8189 ^ n8068 ^ n7537 ;
  assign n8191 = ( n7537 & n8068 ) | ( n7537 & n8189 ) | ( n8068 & n8189 ) ;
  assign n8192 = x103 & n3734 ;
  assign n8193 = ( x105 & n3732 ) | ( x105 & n8192 ) | ( n3732 & n8192 ) ;
  assign n8194 = n8192 | n8193 ;
  assign n8195 = x104 & ~n3737 ;
  assign n8196 = ( x104 & n8194 ) | ( x104 & ~n8195 ) | ( n8194 & ~n8195 ) ;
  assign n8197 = n3736 & n8105 ;
  assign n8198 = n8196 | n8197 ;
  assign n8199 = n8198 ^ x26 ^ 1'b0 ;
  assign n8200 = n8199 ^ n8079 ^ n7804 ;
  assign n8201 = ( n7804 & n8079 ) | ( n7804 & n8199 ) | ( n8079 & n8199 ) ;
  assign n8202 = x102 & n5499 ;
  assign n8203 = ( x104 & n5497 ) | ( x104 & n8202 ) | ( n5497 & n8202 ) ;
  assign n8204 = n8202 | n8203 ;
  assign n8205 = x103 & ~n5502 ;
  assign n8206 = ( x103 & n8204 ) | ( x103 & ~n8205 ) | ( n8204 & ~n8205 ) ;
  assign n8207 = n5501 & n8012 ;
  assign n8208 = n8206 | n8207 ;
  assign n8209 = n8208 ^ x11 ^ 1'b0 ;
  assign n8210 = ( n7518 & n7966 ) | ( n7518 & n8209 ) | ( n7966 & n8209 ) ;
  assign n8211 = n8209 ^ n7966 ^ n7518 ;
  assign n8212 = x103 & n5499 ;
  assign n8213 = ( x105 & n5497 ) | ( x105 & n8212 ) | ( n5497 & n8212 ) ;
  assign n8214 = n8212 | n8213 ;
  assign n8215 = x104 & ~n5502 ;
  assign n8216 = ( x104 & n8214 ) | ( x104 & ~n8215 ) | ( n8214 & ~n8215 ) ;
  assign n8217 = n5501 & n8105 ;
  assign n8218 = n8216 | n8217 ;
  assign n8219 = n8218 ^ x11 ^ 1'b0 ;
  assign n8220 = ( n7833 & n8210 ) | ( n7833 & n8219 ) | ( n8210 & n8219 ) ;
  assign n8221 = n8219 ^ n8210 ^ n7833 ;
  assign n8222 = x102 & n4790 ;
  assign n8223 = ( x104 & n4792 ) | ( x104 & n8222 ) | ( n4792 & n8222 ) ;
  assign n8224 = n8222 | n8223 ;
  assign n8225 = x103 & ~n4786 ;
  assign n8226 = ( x103 & n8224 ) | ( x103 & ~n8225 ) | ( n8224 & ~n8225 ) ;
  assign n8227 = n4787 & n8012 ;
  assign n8228 = n8226 | n8227 ;
  assign n8229 = n8228 ^ x20 ^ 1'b0 ;
  assign n8230 = ( n7744 & n7996 ) | ( n7744 & n8229 ) | ( n7996 & n8229 ) ;
  assign n8231 = n8229 ^ n7996 ^ n7744 ;
  assign n8232 = x102 & n2560 ;
  assign n8233 = ( x104 & n2567 ) | ( x104 & n8232 ) | ( n2567 & n8232 ) ;
  assign n8234 = n8232 | n8233 ;
  assign n8235 = x103 & ~n2562 ;
  assign n8236 = ( x103 & n8234 ) | ( x103 & ~n8235 ) | ( n8234 & ~n8235 ) ;
  assign n8237 = n2565 & n8012 ;
  assign n8238 = n8236 | n8237 ;
  assign n8239 = n8238 ^ x35 ^ 1'b0 ;
  assign n8240 = ( n4339 & n7814 ) | ( n4339 & n8239 ) | ( n7814 & n8239 ) ;
  assign n8241 = n8239 ^ n7814 ^ n4339 ;
  assign n8242 = x103 & n4790 ;
  assign n8243 = ( x105 & n4792 ) | ( x105 & n8242 ) | ( n4792 & n8242 ) ;
  assign n8244 = n8242 | n8243 ;
  assign n8245 = x104 & ~n4786 ;
  assign n8246 = ( x104 & n8244 ) | ( x104 & ~n8245 ) | ( n8244 & ~n8245 ) ;
  assign n8247 = n4787 & n8105 ;
  assign n8248 = n8246 | n8247 ;
  assign n8249 = n8248 ^ x20 ^ 1'b0 ;
  assign n8250 = ( n7753 & n8230 ) | ( n7753 & n8249 ) | ( n8230 & n8249 ) ;
  assign n8251 = n8249 ^ n8230 ^ n7753 ;
  assign n8252 = x102 & n3025 ;
  assign n8253 = ( x104 & n3015 ) | ( x104 & n8252 ) | ( n3015 & n8252 ) ;
  assign n8254 = n8252 | n8253 ;
  assign n8255 = x103 & ~n3014 ;
  assign n8256 = ( x103 & n8254 ) | ( x103 & ~n8255 ) | ( n8254 & ~n8255 ) ;
  assign n8257 = n3017 & n8012 ;
  assign n8258 = n8256 | n8257 ;
  assign n8259 = n8258 ^ x32 ^ 1'b0 ;
  assign n8260 = ( n4379 & n7854 ) | ( n4379 & n8259 ) | ( n7854 & n8259 ) ;
  assign n8261 = n8259 ^ n7854 ^ n4379 ;
  assign n8262 = x103 & n4972 ;
  assign n8263 = ( x105 & n4985 ) | ( x105 & n8262 ) | ( n4985 & n8262 ) ;
  assign n8264 = n8262 | n8263 ;
  assign n8265 = x104 & ~n4980 ;
  assign n8266 = n4987 & n8105 ;
  assign n8267 = ( x104 & n8264 ) | ( x104 & ~n8265 ) | ( n8264 & ~n8265 ) ;
  assign n8268 = x102 & n1058 ;
  assign n8269 = n8266 | n8267 ;
  assign n8270 = ( x104 & n1065 ) | ( x104 & n8268 ) | ( n1065 & n8268 ) ;
  assign n8271 = n8268 | n8270 ;
  assign n8272 = x103 & ~n1060 ;
  assign n8273 = ( x103 & n8271 ) | ( x103 & ~n8272 ) | ( n8271 & ~n8272 ) ;
  assign n8274 = n1063 & n8012 ;
  assign n8275 = n8273 | n8274 ;
  assign n8276 = n8275 ^ x41 ^ 1'b0 ;
  assign n8277 = n8269 ^ x14 ^ 1'b0 ;
  assign n8278 = n8277 ^ n8099 ^ n7793 ;
  assign n8279 = ( n7793 & n8099 ) | ( n7793 & n8277 ) | ( n8099 & n8277 ) ;
  assign n8280 = x104 & n1058 ;
  assign n8281 = ( x106 & n1065 ) | ( x106 & n8280 ) | ( n1065 & n8280 ) ;
  assign n8282 = n8280 | n8281 ;
  assign n8283 = x105 & ~n1060 ;
  assign n8284 = ( x105 & n8282 ) | ( x105 & ~n8283 ) | ( n8282 & ~n8283 ) ;
  assign n8285 = ( n4369 & n5713 ) | ( n4369 & n8276 ) | ( n5713 & n8276 ) ;
  assign n8286 = n8276 ^ n5713 ^ n4369 ;
  assign n8287 = n8143 ^ x106 ^ x105 ;
  assign n8288 = n1063 & n8287 ;
  assign n8289 = n8284 | n8288 ;
  assign n8290 = n8289 ^ x41 ^ 1'b0 ;
  assign n8291 = n8290 ^ n8109 ^ n7876 ;
  assign n8292 = ( n7876 & n8109 ) | ( n7876 & n8290 ) | ( n8109 & n8290 ) ;
  assign n8293 = x103 & n2156 ;
  assign n8294 = ( x105 & n2163 ) | ( x105 & n8293 ) | ( n2163 & n8293 ) ;
  assign n8295 = n8293 | n8294 ;
  assign n8296 = x104 & ~n2158 ;
  assign n8297 = ( x104 & n8295 ) | ( x104 & ~n8296 ) | ( n8295 & ~n8296 ) ;
  assign n8298 = n2161 & n8105 ;
  assign n8299 = n8297 | n8298 ;
  assign n8300 = n8299 ^ x38 ^ 1'b0 ;
  assign n8301 = n8300 ^ n5953 ^ n5692 ;
  assign n8302 = ( n5692 & n5953 ) | ( n5692 & n8300 ) | ( n5953 & n8300 ) ;
  assign n8303 = x104 & n3025 ;
  assign n8304 = ( x106 & n3015 ) | ( x106 & n8303 ) | ( n3015 & n8303 ) ;
  assign n8305 = n8303 | n8304 ;
  assign n8306 = x105 & ~n3014 ;
  assign n8307 = ( x105 & n8305 ) | ( x105 & ~n8306 ) | ( n8305 & ~n8306 ) ;
  assign n8308 = n3017 & n8287 ;
  assign n8309 = n8307 | n8308 ;
  assign n8310 = n8309 ^ x32 ^ 1'b0 ;
  assign n8311 = n8310 ^ n8151 ^ n7864 ;
  assign n8312 = ( n7864 & n8151 ) | ( n7864 & n8310 ) | ( n8151 & n8310 ) ;
  assign n8313 = x104 & n2560 ;
  assign n8314 = ( x106 & n2567 ) | ( x106 & n8313 ) | ( n2567 & n8313 ) ;
  assign n8315 = n8313 | n8314 ;
  assign n8316 = x105 & ~n2562 ;
  assign n8317 = ( x105 & n8315 ) | ( x105 & ~n8316 ) | ( n8315 & ~n8316 ) ;
  assign n8318 = n2565 & n8287 ;
  assign n8319 = n8317 | n8318 ;
  assign n8320 = n8319 ^ x35 ^ 1'b0 ;
  assign n8321 = ( n7896 & n8160 ) | ( n7896 & n8320 ) | ( n8160 & n8320 ) ;
  assign n8322 = n8320 ^ n8160 ^ n7896 ;
  assign n8323 = x104 & n5499 ;
  assign n8324 = ( x106 & n5497 ) | ( x106 & n8323 ) | ( n5497 & n8323 ) ;
  assign n8325 = n8323 | n8324 ;
  assign n8326 = x105 & ~n5502 ;
  assign n8327 = ( x105 & n8325 ) | ( x105 & ~n8326 ) | ( n8325 & ~n8326 ) ;
  assign n8328 = n5501 & n8287 ;
  assign n8329 = n8327 | n8328 ;
  assign n8330 = n8329 ^ x11 ^ 1'b0 ;
  assign n8331 = ( n7987 & n8220 ) | ( n7987 & n8330 ) | ( n8220 & n8330 ) ;
  assign n8332 = n8330 ^ n8220 ^ n7987 ;
  assign n8333 = x104 & n5979 ;
  assign n8334 = ( x106 & n5969 ) | ( x106 & n8333 ) | ( n5969 & n8333 ) ;
  assign n8335 = n8333 | n8334 ;
  assign n8336 = x105 & ~n5970 ;
  assign n8337 = ( x105 & n8335 ) | ( x105 & ~n8336 ) | ( n8335 & ~n8336 ) ;
  assign n8338 = n5968 & n8287 ;
  assign n8339 = n8337 | n8338 ;
  assign n8340 = n8339 ^ x5 ^ 1'b0 ;
  assign n8341 = n8340 ^ n8140 ^ n7936 ;
  assign n8342 = ( n7936 & n8140 ) | ( n7936 & n8340 ) | ( n8140 & n8340 ) ;
  assign n8343 = x104 & n4790 ;
  assign n8344 = ( x106 & n4792 ) | ( x106 & n8343 ) | ( n4792 & n8343 ) ;
  assign n8345 = n8343 | n8344 ;
  assign n8346 = x105 & ~n4786 ;
  assign n8347 = ( x105 & n8345 ) | ( x105 & ~n8346 ) | ( n8345 & ~n8346 ) ;
  assign n8348 = n4787 & n8287 ;
  assign n8349 = n8347 | n8348 ;
  assign n8350 = ( x105 & x106 ) | ( x105 & n8143 ) | ( x106 & n8143 ) ;
  assign n8351 = n8349 ^ x20 ^ 1'b0 ;
  assign n8352 = ( n7975 & n8250 ) | ( n7975 & n8351 ) | ( n8250 & n8351 ) ;
  assign n8353 = n8351 ^ n8250 ^ n7975 ;
  assign n8354 = x104 & n5011 ;
  assign n8355 = ( x106 & n5012 ) | ( x106 & n8354 ) | ( n5012 & n8354 ) ;
  assign n8356 = n8354 | n8355 ;
  assign n8357 = x105 & ~n5008 ;
  assign n8358 = ( x105 & n8356 ) | ( x105 & ~n8357 ) | ( n8356 & ~n8357 ) ;
  assign n8359 = n5020 & n8287 ;
  assign n8360 = n8358 | n8359 ;
  assign n8361 = n8360 ^ x17 ^ 1'b0 ;
  assign n8362 = n8361 ^ n8170 ^ n7997 ;
  assign n8363 = ( n7997 & n8170 ) | ( n7997 & n8361 ) | ( n8170 & n8361 ) ;
  assign n8364 = x104 & n3344 ;
  assign n8365 = ( x106 & n3342 ) | ( x106 & n8364 ) | ( n3342 & n8364 ) ;
  assign n8366 = n8364 | n8365 ;
  assign n8367 = x105 & ~n3347 ;
  assign n8368 = ( x105 & n8366 ) | ( x105 & ~n8367 ) | ( n8366 & ~n8367 ) ;
  assign n8369 = n3346 & n8287 ;
  assign n8370 = n8368 | n8369 ;
  assign n8371 = n8370 ^ x29 ^ 1'b0 ;
  assign n8372 = ( n7946 & n8181 ) | ( n7946 & n8371 ) | ( n8181 & n8371 ) ;
  assign n8373 = n8371 ^ n8181 ^ n7946 ;
  assign n8374 = x104 & n3734 ;
  assign n8375 = ( x106 & n3732 ) | ( x106 & n8374 ) | ( n3732 & n8374 ) ;
  assign n8376 = n8374 | n8375 ;
  assign n8377 = x105 & ~n3737 ;
  assign n8378 = ( x105 & n8376 ) | ( x105 & ~n8377 ) | ( n8376 & ~n8377 ) ;
  assign n8379 = n3736 & n8287 ;
  assign n8380 = n8378 | n8379 ;
  assign n8381 = n8380 ^ x26 ^ 1'b0 ;
  assign n8382 = ( n7803 & n7926 ) | ( n7803 & n8381 ) | ( n7926 & n8381 ) ;
  assign n8383 = n8381 ^ n7926 ^ n7803 ;
  assign n8384 = x104 & n4972 ;
  assign n8385 = ( x106 & n4985 ) | ( x106 & n8384 ) | ( n4985 & n8384 ) ;
  assign n8386 = n8384 | n8385 ;
  assign n8387 = x105 & ~n4980 ;
  assign n8388 = ( x105 & n8386 ) | ( x105 & ~n8387 ) | ( n8386 & ~n8387 ) ;
  assign n8389 = n4987 & n8287 ;
  assign n8390 = n8388 | n8389 ;
  assign n8391 = n8390 ^ x14 ^ 1'b0 ;
  assign n8392 = ( n7916 & n8279 ) | ( n7916 & n8391 ) | ( n8279 & n8391 ) ;
  assign n8393 = n8391 ^ n8279 ^ n7916 ;
  assign n8394 = x104 & n6104 ;
  assign n8395 = ( x106 & n6105 ) | ( x106 & n8394 ) | ( n6105 & n8394 ) ;
  assign n8396 = n8394 | n8395 ;
  assign n8397 = x105 & ~n6107 ;
  assign n8398 = ( x105 & n8396 ) | ( x105 & ~n8397 ) | ( n8396 & ~n8397 ) ;
  assign n8399 = ~n6108 & n8287 ;
  assign n8400 = ( n8287 & n8398 ) | ( n8287 & ~n8399 ) | ( n8398 & ~n8399 ) ;
  assign n8401 = n8400 ^ x2 ^ 1'b0 ;
  assign n8402 = ( n7905 & n8119 ) | ( n7905 & n8401 ) | ( n8119 & n8401 ) ;
  assign n8403 = n8401 ^ n8119 ^ n7905 ;
  assign n8404 = x104 & n2156 ;
  assign n8405 = ( x106 & n2163 ) | ( x106 & n8404 ) | ( n2163 & n8404 ) ;
  assign n8406 = n8404 | n8405 ;
  assign n8407 = x105 & ~n2158 ;
  assign n8408 = ( x105 & n8406 ) | ( x105 & ~n8407 ) | ( n8406 & ~n8407 ) ;
  assign n8409 = n2161 & n8287 ;
  assign n8410 = n8408 | n8409 ;
  assign n8411 = n8410 ^ x38 ^ 1'b0 ;
  assign n8412 = ( n7885 & n8302 ) | ( n7885 & n8411 ) | ( n8302 & n8411 ) ;
  assign n8413 = n8411 ^ n8302 ^ n7885 ;
  assign n8414 = x104 & n4616 ;
  assign n8415 = ( x106 & n4606 ) | ( x106 & n8414 ) | ( n4606 & n8414 ) ;
  assign n8416 = n8414 | n8415 ;
  assign n8417 = x105 & ~n4605 ;
  assign n8418 = ( x105 & n8416 ) | ( x105 & ~n8417 ) | ( n8416 & ~n8417 ) ;
  assign n8419 = n4608 & n8287 ;
  assign n8420 = n8418 | n8419 ;
  assign n8421 = n8420 ^ x23 ^ 1'b0 ;
  assign n8422 = ( n7955 & n8129 ) | ( n7955 & n8421 ) | ( n8129 & n8421 ) ;
  assign n8423 = n8421 ^ n8129 ^ n7955 ;
  assign n8424 = x104 & n5718 ;
  assign n8425 = ( x106 & n5720 ) | ( x106 & n8424 ) | ( n5720 & n8424 ) ;
  assign n8426 = n8424 | n8425 ;
  assign n8427 = x105 & ~n5727 ;
  assign n8428 = ( x105 & n8426 ) | ( x105 & ~n8427 ) | ( n8426 & ~n8427 ) ;
  assign n8429 = n5726 & n8287 ;
  assign n8430 = n8428 | n8429 ;
  assign n8431 = n8430 ^ x8 ^ 1'b0 ;
  assign n8432 = n8431 ^ n8191 ^ n7965 ;
  assign n8433 = ( n7965 & n8191 ) | ( n7965 & n8431 ) | ( n8191 & n8431 ) ;
  assign n8434 = x105 & n2156 ;
  assign n8435 = ( x107 & n2163 ) | ( x107 & n8434 ) | ( n2163 & n8434 ) ;
  assign n8436 = x105 & n3344 ;
  assign n8437 = ( x107 & n3342 ) | ( x107 & n8436 ) | ( n3342 & n8436 ) ;
  assign n8438 = n8434 | n8435 ;
  assign n8439 = n8436 | n8437 ;
  assign n8440 = n8350 ^ x107 ^ x106 ;
  assign n8441 = x106 & ~n2158 ;
  assign n8442 = ( x106 & n8438 ) | ( x106 & ~n8441 ) | ( n8438 & ~n8441 ) ;
  assign n8443 = x106 & ~n3347 ;
  assign n8444 = ( x106 & n8439 ) | ( x106 & ~n8443 ) | ( n8439 & ~n8443 ) ;
  assign n8445 = n2161 & n8440 ;
  assign n8446 = n8442 | n8445 ;
  assign n8447 = n3346 & n8440 ;
  assign n8448 = n8444 | n8447 ;
  assign n8449 = n8448 ^ x29 ^ 1'b0 ;
  assign n8450 = ( n7945 & n8261 ) | ( n7945 & n8449 ) | ( n8261 & n8449 ) ;
  assign n8451 = n8449 ^ n8261 ^ n7945 ;
  assign n8452 = x105 & n5011 ;
  assign n8453 = ( x107 & n5012 ) | ( x107 & n8452 ) | ( n5012 & n8452 ) ;
  assign n8454 = n8452 | n8453 ;
  assign n8455 = x106 & ~n5008 ;
  assign n8456 = ( x106 & n8454 ) | ( x106 & ~n8455 ) | ( n8454 & ~n8455 ) ;
  assign n8457 = n5020 & n8440 ;
  assign n8458 = n8456 | n8457 ;
  assign n8459 = n8458 ^ x17 ^ 1'b0 ;
  assign n8460 = n8446 ^ x38 ^ 1'b0 ;
  assign n8461 = n8459 ^ n8363 ^ n8231 ;
  assign n8462 = ( n8231 & n8363 ) | ( n8231 & n8459 ) | ( n8363 & n8459 ) ;
  assign n8463 = n8460 ^ n8286 ^ n7886 ;
  assign n8464 = x105 & n6104 ;
  assign n8465 = ( n7886 & n8286 ) | ( n7886 & n8460 ) | ( n8286 & n8460 ) ;
  assign n8466 = ( x107 & n6105 ) | ( x107 & n8464 ) | ( n6105 & n8464 ) ;
  assign n8467 = n8464 | n8466 ;
  assign n8468 = ( x106 & x107 ) | ( x106 & n8350 ) | ( x107 & n8350 ) ;
  assign n8469 = x106 & ~n6107 ;
  assign n8470 = ( x106 & n8467 ) | ( x106 & ~n8469 ) | ( n8467 & ~n8469 ) ;
  assign n8471 = ~n6108 & n8440 ;
  assign n8472 = ( n8440 & n8470 ) | ( n8440 & ~n8471 ) | ( n8470 & ~n8471 ) ;
  assign n8473 = n8472 ^ x2 ^ 1'b0 ;
  assign n8474 = ( n8088 & n8402 ) | ( n8088 & n8473 ) | ( n8402 & n8473 ) ;
  assign n8475 = n8473 ^ n8402 ^ n8088 ;
  assign n8476 = x105 & n5718 ;
  assign n8477 = ( x107 & n5720 ) | ( x107 & n8476 ) | ( n5720 & n8476 ) ;
  assign n8478 = x106 & ~n5727 ;
  assign n8479 = n8476 | n8477 ;
  assign n8480 = x105 & n3025 ;
  assign n8481 = ( x106 & ~n8478 ) | ( x106 & n8479 ) | ( ~n8478 & n8479 ) ;
  assign n8482 = n5726 & n8440 ;
  assign n8483 = n8481 | n8482 ;
  assign n8484 = ( x107 & n3015 ) | ( x107 & n8480 ) | ( n3015 & n8480 ) ;
  assign n8485 = n8480 | n8484 ;
  assign n8486 = x106 & ~n3014 ;
  assign n8487 = ( x106 & n8485 ) | ( x106 & ~n8486 ) | ( n8485 & ~n8486 ) ;
  assign n8488 = n8483 ^ x8 ^ 1'b0 ;
  assign n8489 = n3017 & n8440 ;
  assign n8490 = n8487 | n8489 ;
  assign n8491 = n8490 ^ x32 ^ 1'b0 ;
  assign n8492 = n8488 ^ n8433 ^ n8211 ;
  assign n8493 = ( n8211 & n8433 ) | ( n8211 & n8488 ) | ( n8433 & n8488 ) ;
  assign n8494 = n8491 ^ n8241 ^ n7865 ;
  assign n8495 = ( n7865 & n8241 ) | ( n7865 & n8491 ) | ( n8241 & n8491 ) ;
  assign n8496 = x105 & n4616 ;
  assign n8497 = ( x107 & n4606 ) | ( x107 & n8496 ) | ( n4606 & n8496 ) ;
  assign n8498 = n8496 | n8497 ;
  assign n8499 = x106 & ~n4605 ;
  assign n8500 = ( x106 & n8498 ) | ( x106 & ~n8499 ) | ( n8498 & ~n8499 ) ;
  assign n8501 = n4608 & n8440 ;
  assign n8502 = n8500 | n8501 ;
  assign n8503 = n8502 ^ x23 ^ 1'b0 ;
  assign n8504 = ( n8078 & n8422 ) | ( n8078 & n8503 ) | ( n8422 & n8503 ) ;
  assign n8505 = n8503 ^ n8422 ^ n8078 ;
  assign n8506 = x105 & n4972 ;
  assign n8507 = ( x107 & n4985 ) | ( x107 & n8506 ) | ( n4985 & n8506 ) ;
  assign n8508 = n8506 | n8507 ;
  assign n8509 = x106 & ~n4980 ;
  assign n8510 = ( x106 & n8508 ) | ( x106 & ~n8509 ) | ( n8508 & ~n8509 ) ;
  assign n8511 = n4987 & n8440 ;
  assign n8512 = n8510 | n8511 ;
  assign n8513 = n8512 ^ x14 ^ 1'b0 ;
  assign n8514 = ( n8017 & n8392 ) | ( n8017 & n8513 ) | ( n8392 & n8513 ) ;
  assign n8515 = n8513 ^ n8392 ^ n8017 ;
  assign n8516 = x105 & n5979 ;
  assign n8517 = ( x107 & n5969 ) | ( x107 & n8516 ) | ( n5969 & n8516 ) ;
  assign n8518 = n8516 | n8517 ;
  assign n8519 = x106 & ~n5970 ;
  assign n8520 = ( x106 & n8518 ) | ( x106 & ~n8519 ) | ( n8518 & ~n8519 ) ;
  assign n8521 = n5968 & n8440 ;
  assign n8522 = n8520 | n8521 ;
  assign n8523 = n8522 ^ x5 ^ 1'b0 ;
  assign n8524 = ( n8069 & n8342 ) | ( n8069 & n8523 ) | ( n8342 & n8523 ) ;
  assign n8525 = n8523 ^ n8342 ^ n8069 ;
  assign n8526 = x105 & n3734 ;
  assign n8527 = ( x107 & n3732 ) | ( x107 & n8526 ) | ( n3732 & n8526 ) ;
  assign n8528 = n8526 | n8527 ;
  assign n8529 = x106 & ~n3737 ;
  assign n8530 = ( x106 & n8528 ) | ( x106 & ~n8529 ) | ( n8528 & ~n8529 ) ;
  assign n8531 = n3736 & n8440 ;
  assign n8532 = n8530 | n8531 ;
  assign n8533 = n8532 ^ x26 ^ 1'b0 ;
  assign n8534 = ( n7925 & n8038 ) | ( n7925 & n8533 ) | ( n8038 & n8533 ) ;
  assign n8535 = n8533 ^ n8038 ^ n7925 ;
  assign n8536 = x105 & n4790 ;
  assign n8537 = ( x107 & n4792 ) | ( x107 & n8536 ) | ( n4792 & n8536 ) ;
  assign n8538 = n8536 | n8537 ;
  assign n8539 = x106 & ~n4786 ;
  assign n8540 = ( x106 & n8538 ) | ( x106 & ~n8539 ) | ( n8538 & ~n8539 ) ;
  assign n8541 = n4787 & n8440 ;
  assign n8542 = n8540 | n8541 ;
  assign n8543 = n8542 ^ x20 ^ 1'b0 ;
  assign n8544 = ( n8027 & n8352 ) | ( n8027 & n8543 ) | ( n8352 & n8543 ) ;
  assign n8545 = n8543 ^ n8352 ^ n8027 ;
  assign n8546 = x105 & n5499 ;
  assign n8547 = ( x107 & n5497 ) | ( x107 & n8546 ) | ( n5497 & n8546 ) ;
  assign n8548 = n8546 | n8547 ;
  assign n8549 = x106 & ~n5502 ;
  assign n8550 = ( x106 & n8548 ) | ( x106 & ~n8549 ) | ( n8548 & ~n8549 ) ;
  assign n8551 = n5501 & n8440 ;
  assign n8552 = n8550 | n8551 ;
  assign n8553 = n8552 ^ x11 ^ 1'b0 ;
  assign n8554 = n8553 ^ n8331 ^ n8098 ;
  assign n8555 = ( n8098 & n8331 ) | ( n8098 & n8553 ) | ( n8331 & n8553 ) ;
  assign n8556 = x106 & n4616 ;
  assign n8557 = n8468 ^ x108 ^ x107 ;
  assign n8558 = ( x108 & n4606 ) | ( x108 & n8556 ) | ( n4606 & n8556 ) ;
  assign n8559 = n8556 | n8558 ;
  assign n8560 = x107 & ~n4605 ;
  assign n8561 = ( x107 & n8559 ) | ( x107 & ~n8560 ) | ( n8559 & ~n8560 ) ;
  assign n8562 = n4608 & n8557 ;
  assign n8563 = n8561 | n8562 ;
  assign n8564 = n8563 ^ x23 ^ 1'b0 ;
  assign n8565 = n8564 ^ n8504 ^ n8200 ;
  assign n8566 = ( n8200 & n8504 ) | ( n8200 & n8564 ) | ( n8504 & n8564 ) ;
  assign n8567 = x106 & n6104 ;
  assign n8568 = ( x108 & n6105 ) | ( x108 & n8567 ) | ( n6105 & n8567 ) ;
  assign n8569 = n8567 | n8568 ;
  assign n8570 = x107 & ~n6107 ;
  assign n8571 = ( x107 & n8569 ) | ( x107 & ~n8570 ) | ( n8569 & ~n8570 ) ;
  assign n8572 = ~n6108 & n8557 ;
  assign n8573 = ( n8557 & n8571 ) | ( n8557 & ~n8572 ) | ( n8571 & ~n8572 ) ;
  assign n8574 = n8573 ^ x2 ^ 1'b0 ;
  assign n8575 = n8574 ^ n8474 ^ n8139 ;
  assign n8576 = ( n8139 & n8474 ) | ( n8139 & n8574 ) | ( n8474 & n8574 ) ;
  assign n8577 = x106 & n2560 ;
  assign n8578 = ( x108 & n2567 ) | ( x108 & n8577 ) | ( n2567 & n8577 ) ;
  assign n8579 = n8577 | n8578 ;
  assign n8580 = x107 & ~n2562 ;
  assign n8581 = ( x107 & n8579 ) | ( x107 & ~n8580 ) | ( n8579 & ~n8580 ) ;
  assign n8582 = n2565 & n8557 ;
  assign n8583 = n8581 | n8582 ;
  assign n8584 = n8583 ^ x35 ^ 1'b0 ;
  assign n8585 = ( x107 & x108 ) | ( x107 & n8468 ) | ( x108 & n8468 ) ;
  assign n8586 = ( n8058 & n8301 ) | ( n8058 & n8584 ) | ( n8301 & n8584 ) ;
  assign n8587 = n8584 ^ n8301 ^ n8058 ;
  assign n8588 = x106 & n3025 ;
  assign n8589 = ( x108 & n3015 ) | ( x108 & n8588 ) | ( n3015 & n8588 ) ;
  assign n8590 = n8588 | n8589 ;
  assign n8591 = x107 & ~n3014 ;
  assign n8592 = ( x107 & n8590 ) | ( x107 & ~n8591 ) | ( n8590 & ~n8591 ) ;
  assign n8593 = ( n3017 & n8557 ) | ( n3017 & n8592 ) | ( n8557 & n8592 ) ;
  assign n8594 = n8592 | n8593 ;
  assign n8595 = n8594 ^ x32 ^ 1'b0 ;
  assign n8596 = n8595 ^ n8240 ^ n8161 ;
  assign n8597 = ( n8161 & n8240 ) | ( n8161 & n8595 ) | ( n8240 & n8595 ) ;
  assign n8598 = x105 & n2560 ;
  assign n8599 = ( x107 & n2567 ) | ( x107 & n8598 ) | ( n2567 & n8598 ) ;
  assign n8600 = n8598 | n8599 ;
  assign n8601 = x106 & ~n2562 ;
  assign n8602 = ( x106 & n8600 ) | ( x106 & ~n8601 ) | ( n8600 & ~n8601 ) ;
  assign n8603 = n2565 & n8440 ;
  assign n8604 = n8602 | n8603 ;
  assign n8605 = n8604 ^ x35 ^ 1'b0 ;
  assign n8606 = n8605 ^ n8059 ^ n7895 ;
  assign n8607 = ( n7895 & n8059 ) | ( n7895 & n8605 ) | ( n8059 & n8605 ) ;
  assign n8608 = x106 & n5011 ;
  assign n8609 = ( x108 & n5012 ) | ( x108 & n8608 ) | ( n5012 & n8608 ) ;
  assign n8610 = n8608 | n8609 ;
  assign n8611 = x107 & ~n5008 ;
  assign n8612 = ( x107 & n8610 ) | ( x107 & ~n8611 ) | ( n8610 & ~n8611 ) ;
  assign n8613 = n5020 & n8557 ;
  assign n8614 = n8612 | n8613 ;
  assign n8615 = n8614 ^ x17 ^ 1'b0 ;
  assign n8616 = ( n8251 & n8462 ) | ( n8251 & n8615 ) | ( n8462 & n8615 ) ;
  assign n8617 = n8615 ^ n8462 ^ n8251 ;
  assign n8618 = x106 & n5499 ;
  assign n8619 = ( x108 & n5497 ) | ( x108 & n8618 ) | ( n5497 & n8618 ) ;
  assign n8620 = n8618 | n8619 ;
  assign n8621 = x107 & ~n5502 ;
  assign n8622 = ( x107 & n8620 ) | ( x107 & ~n8621 ) | ( n8620 & ~n8621 ) ;
  assign n8623 = n5501 & n8557 ;
  assign n8624 = n8622 | n8623 ;
  assign n8625 = n8624 ^ x11 ^ 1'b0 ;
  assign n8626 = ( n8278 & n8555 ) | ( n8278 & n8625 ) | ( n8555 & n8625 ) ;
  assign n8627 = n8625 ^ n8555 ^ n8278 ;
  assign n8628 = x106 & n5979 ;
  assign n8629 = ( x108 & n5969 ) | ( x108 & n8628 ) | ( n5969 & n8628 ) ;
  assign n8630 = n8628 | n8629 ;
  assign n8631 = x107 & ~n5970 ;
  assign n8632 = ( x107 & n8630 ) | ( x107 & ~n8631 ) | ( n8630 & ~n8631 ) ;
  assign n8633 = n5968 & n8557 ;
  assign n8634 = n8632 | n8633 ;
  assign n8635 = n8634 ^ x5 ^ 1'b0 ;
  assign n8636 = ( n8190 & n8524 ) | ( n8190 & n8635 ) | ( n8524 & n8635 ) ;
  assign n8637 = n8635 ^ n8524 ^ n8190 ;
  assign n8638 = x106 & n4790 ;
  assign n8639 = ( x108 & n4792 ) | ( x108 & n8638 ) | ( n4792 & n8638 ) ;
  assign n8640 = n8638 | n8639 ;
  assign n8641 = x107 & ~n4786 ;
  assign n8642 = ( x107 & n8640 ) | ( x107 & ~n8641 ) | ( n8640 & ~n8641 ) ;
  assign n8643 = n4787 & n8557 ;
  assign n8644 = n8642 | n8643 ;
  assign n8645 = n8644 ^ x20 ^ 1'b0 ;
  assign n8646 = ( n8130 & n8544 ) | ( n8130 & n8645 ) | ( n8544 & n8645 ) ;
  assign n8647 = n8645 ^ n8544 ^ n8130 ;
  assign n8648 = x106 & n4972 ;
  assign n8649 = ( x108 & n4985 ) | ( x108 & n8648 ) | ( n4985 & n8648 ) ;
  assign n8650 = n8648 | n8649 ;
  assign n8651 = x107 & ~n4980 ;
  assign n8652 = ( x107 & n8650 ) | ( x107 & ~n8651 ) | ( n8650 & ~n8651 ) ;
  assign n8653 = n4987 & n8557 ;
  assign n8654 = n8652 | n8653 ;
  assign n8655 = n8654 ^ x14 ^ 1'b0 ;
  assign n8656 = ( n8171 & n8514 ) | ( n8171 & n8655 ) | ( n8514 & n8655 ) ;
  assign n8657 = n8655 ^ n8514 ^ n8171 ;
  assign n8658 = x106 & n5718 ;
  assign n8659 = ( x108 & n5720 ) | ( x108 & n8658 ) | ( n5720 & n8658 ) ;
  assign n8660 = n8658 | n8659 ;
  assign n8661 = x107 & ~n5727 ;
  assign n8662 = ( x107 & n8660 ) | ( x107 & ~n8661 ) | ( n8660 & ~n8661 ) ;
  assign n8663 = n5726 & n8557 ;
  assign n8664 = n8662 | n8663 ;
  assign n8665 = n8664 ^ x8 ^ 1'b0 ;
  assign n8666 = n8665 ^ n8493 ^ n8221 ;
  assign n8667 = ( n8221 & n8493 ) | ( n8221 & n8665 ) | ( n8493 & n8665 ) ;
  assign n8668 = x106 & n3734 ;
  assign n8669 = ( x108 & n3732 ) | ( x108 & n8668 ) | ( n3732 & n8668 ) ;
  assign n8670 = n8668 | n8669 ;
  assign n8671 = x107 & ~n3737 ;
  assign n8672 = ( x107 & n8670 ) | ( x107 & ~n8671 ) | ( n8670 & ~n8671 ) ;
  assign n8673 = ( n3736 & n8557 ) | ( n3736 & n8672 ) | ( n8557 & n8672 ) ;
  assign n8674 = n8672 | n8673 ;
  assign n8675 = n8674 ^ x26 ^ 1'b0 ;
  assign n8676 = x107 & n6104 ;
  assign n8677 = ( n8037 & n8180 ) | ( n8037 & n8675 ) | ( n8180 & n8675 ) ;
  assign n8678 = ( x109 & n6105 ) | ( x109 & n8676 ) | ( n6105 & n8676 ) ;
  assign n8679 = n8675 ^ n8180 ^ n8037 ;
  assign n8680 = n8585 ^ x109 ^ x108 ;
  assign n8681 = ~n6108 & n8680 ;
  assign n8682 = n8676 | n8678 ;
  assign n8683 = x108 & ~n6107 ;
  assign n8684 = ( x108 & n8682 ) | ( x108 & ~n8683 ) | ( n8682 & ~n8683 ) ;
  assign n8685 = ( n8680 & ~n8681 ) | ( n8680 & n8684 ) | ( ~n8681 & n8684 ) ;
  assign n8686 = n8685 ^ x2 ^ 1'b0 ;
  assign n8687 = x107 & n2560 ;
  assign n8688 = ( x109 & n2567 ) | ( x109 & n8687 ) | ( n2567 & n8687 ) ;
  assign n8689 = n8687 | n8688 ;
  assign n8690 = x108 & ~n2562 ;
  assign n8691 = ( x108 & n8689 ) | ( x108 & ~n8690 ) | ( n8689 & ~n8690 ) ;
  assign n8692 = n2565 & n8680 ;
  assign n8693 = n8691 | n8692 ;
  assign n8694 = n8693 ^ x35 ^ 1'b0 ;
  assign n8695 = ( n8413 & n8586 ) | ( n8413 & n8694 ) | ( n8586 & n8694 ) ;
  assign n8696 = n8694 ^ n8586 ^ n8413 ;
  assign n8697 = x107 & n4616 ;
  assign n8698 = ( x109 & n4606 ) | ( x109 & n8697 ) | ( n4606 & n8697 ) ;
  assign n8699 = n8697 | n8698 ;
  assign n8700 = n8686 ^ n8576 ^ n8341 ;
  assign n8701 = ( n8341 & n8576 ) | ( n8341 & n8686 ) | ( n8576 & n8686 ) ;
  assign n8702 = n4608 & n8680 ;
  assign n8703 = x108 & ~n4605 ;
  assign n8704 = ( x108 & n8699 ) | ( x108 & ~n8703 ) | ( n8699 & ~n8703 ) ;
  assign n8705 = x107 & n3025 ;
  assign n8706 = n8702 | n8704 ;
  assign n8707 = n8706 ^ x23 ^ 1'b0 ;
  assign n8708 = ( x109 & n3015 ) | ( x109 & n8705 ) | ( n3015 & n8705 ) ;
  assign n8709 = n8705 | n8708 ;
  assign n8710 = n8707 ^ n8383 ^ n8201 ;
  assign n8711 = ( n8201 & n8383 ) | ( n8201 & n8707 ) | ( n8383 & n8707 ) ;
  assign n8712 = x108 & ~n3014 ;
  assign n8713 = ( x108 & n8709 ) | ( x108 & ~n8712 ) | ( n8709 & ~n8712 ) ;
  assign n8714 = x107 & n3734 ;
  assign n8715 = ( x109 & n3732 ) | ( x109 & n8714 ) | ( n3732 & n8714 ) ;
  assign n8716 = n8714 | n8715 ;
  assign n8717 = x108 & ~n3737 ;
  assign n8718 = ( x108 & n8716 ) | ( x108 & ~n8717 ) | ( n8716 & ~n8717 ) ;
  assign n8719 = n3017 & n8680 ;
  assign n8720 = n8713 | n8719 ;
  assign n8721 = n8720 ^ x32 ^ 1'b0 ;
  assign n8722 = n8721 ^ n8597 ^ n8322 ;
  assign n8723 = ( n8322 & n8597 ) | ( n8322 & n8721 ) | ( n8597 & n8721 ) ;
  assign n8724 = n3736 & n8680 ;
  assign n8725 = n8718 | n8724 ;
  assign n8726 = x106 & n3344 ;
  assign n8727 = ( x108 & n3342 ) | ( x108 & n8726 ) | ( n3342 & n8726 ) ;
  assign n8728 = n8726 | n8727 ;
  assign n8729 = x107 & ~n3347 ;
  assign n8730 = ( x107 & n8728 ) | ( x107 & ~n8729 ) | ( n8728 & ~n8729 ) ;
  assign n8731 = ( n3346 & n8557 ) | ( n3346 & n8730 ) | ( n8557 & n8730 ) ;
  assign n8732 = n8730 | n8731 ;
  assign n8733 = n8725 ^ x26 ^ 1'b0 ;
  assign n8734 = n8732 ^ x29 ^ 1'b0 ;
  assign n8735 = n8734 ^ n8260 ^ n8150 ;
  assign n8736 = ( n8150 & n8260 ) | ( n8150 & n8734 ) | ( n8260 & n8734 ) ;
  assign n8737 = ( n8373 & n8677 ) | ( n8373 & n8733 ) | ( n8677 & n8733 ) ;
  assign n8738 = n8733 ^ n8677 ^ n8373 ;
  assign n8739 = x107 & n4790 ;
  assign n8740 = ( x109 & n4792 ) | ( x109 & n8739 ) | ( n4792 & n8739 ) ;
  assign n8741 = x108 & ~n4786 ;
  assign n8742 = n8739 | n8740 ;
  assign n8743 = ( x108 & ~n8741 ) | ( x108 & n8742 ) | ( ~n8741 & n8742 ) ;
  assign n8744 = x107 & n5979 ;
  assign n8745 = ( x109 & n5969 ) | ( x109 & n8744 ) | ( n5969 & n8744 ) ;
  assign n8746 = n8744 | n8745 ;
  assign n8747 = x108 & ~n5970 ;
  assign n8748 = ( x108 & n8746 ) | ( x108 & ~n8747 ) | ( n8746 & ~n8747 ) ;
  assign n8749 = n5968 & n8680 ;
  assign n8750 = n8748 | n8749 ;
  assign n8751 = n4787 & n8680 ;
  assign n8752 = n8743 | n8751 ;
  assign n8753 = n8752 ^ x20 ^ 1'b0 ;
  assign n8754 = ( n8423 & n8646 ) | ( n8423 & n8753 ) | ( n8646 & n8753 ) ;
  assign n8755 = n8753 ^ n8646 ^ n8423 ;
  assign n8756 = x107 & n5011 ;
  assign n8757 = ( x109 & n5012 ) | ( x109 & n8756 ) | ( n5012 & n8756 ) ;
  assign n8758 = n8756 | n8757 ;
  assign n8759 = x108 & ~n5008 ;
  assign n8760 = ( x108 & n8758 ) | ( x108 & ~n8759 ) | ( n8758 & ~n8759 ) ;
  assign n8761 = n5020 & n8680 ;
  assign n8762 = n8760 | n8761 ;
  assign n8763 = n8762 ^ x17 ^ 1'b0 ;
  assign n8764 = n8763 ^ n8616 ^ n8353 ;
  assign n8765 = ( n8353 & n8616 ) | ( n8353 & n8763 ) | ( n8616 & n8763 ) ;
  assign n8766 = x107 & n4972 ;
  assign n8767 = ( x109 & n4985 ) | ( x109 & n8766 ) | ( n4985 & n8766 ) ;
  assign n8768 = n8766 | n8767 ;
  assign n8769 = x108 & ~n4980 ;
  assign n8770 = ( x108 & n8768 ) | ( x108 & ~n8769 ) | ( n8768 & ~n8769 ) ;
  assign n8771 = n4987 & n8680 ;
  assign n8772 = n8770 | n8771 ;
  assign n8773 = n8772 ^ x14 ^ 1'b0 ;
  assign n8774 = n8750 ^ x5 ^ 1'b0 ;
  assign n8775 = n8774 ^ n8636 ^ n8432 ;
  assign n8776 = ( n8432 & n8636 ) | ( n8432 & n8774 ) | ( n8636 & n8774 ) ;
  assign n8777 = x107 & n3344 ;
  assign n8778 = ( x109 & n3342 ) | ( x109 & n8777 ) | ( n3342 & n8777 ) ;
  assign n8779 = n8777 | n8778 ;
  assign n8780 = x108 & ~n3347 ;
  assign n8781 = ( x108 & n8779 ) | ( x108 & ~n8780 ) | ( n8779 & ~n8780 ) ;
  assign n8782 = n8773 ^ n8656 ^ n8362 ;
  assign n8783 = ( n8362 & n8656 ) | ( n8362 & n8773 ) | ( n8656 & n8773 ) ;
  assign n8784 = x107 & n5499 ;
  assign n8785 = ( x109 & n5497 ) | ( x109 & n8784 ) | ( n5497 & n8784 ) ;
  assign n8786 = n8784 | n8785 ;
  assign n8787 = x108 & ~n5502 ;
  assign n8788 = ( x108 & n8786 ) | ( x108 & ~n8787 ) | ( n8786 & ~n8787 ) ;
  assign n8789 = n5501 & n8680 ;
  assign n8790 = n8788 | n8789 ;
  assign n8791 = n3346 & n8680 ;
  assign n8792 = n8781 | n8791 ;
  assign n8793 = n8790 ^ x11 ^ 1'b0 ;
  assign n8794 = n8792 ^ x29 ^ 1'b0 ;
  assign n8795 = ( n8311 & n8736 ) | ( n8311 & n8794 ) | ( n8736 & n8794 ) ;
  assign n8796 = n8794 ^ n8736 ^ n8311 ;
  assign n8797 = x107 & n5718 ;
  assign n8798 = ( x109 & n5720 ) | ( x109 & n8797 ) | ( n5720 & n8797 ) ;
  assign n8799 = n8797 | n8798 ;
  assign n8800 = n8793 ^ n8626 ^ n8393 ;
  assign n8801 = ( n8393 & n8626 ) | ( n8393 & n8793 ) | ( n8626 & n8793 ) ;
  assign n8802 = x108 & ~n5727 ;
  assign n8803 = n5726 & n8680 ;
  assign n8804 = ( x108 & n8799 ) | ( x108 & ~n8802 ) | ( n8799 & ~n8802 ) ;
  assign n8805 = n8803 | n8804 ;
  assign n8806 = n8805 ^ x8 ^ 1'b0 ;
  assign n8807 = ( n8332 & n8667 ) | ( n8332 & n8806 ) | ( n8667 & n8806 ) ;
  assign n8808 = n8806 ^ n8667 ^ n8332 ;
  assign n8809 = x109 & ~n5008 ;
  assign n8810 = x108 & n5011 ;
  assign n8811 = ( x110 & n5012 ) | ( x110 & n8810 ) | ( n5012 & n8810 ) ;
  assign n8812 = n8810 | n8811 ;
  assign n8813 = x108 & n2560 ;
  assign n8814 = ( x109 & ~n8809 ) | ( x109 & n8812 ) | ( ~n8809 & n8812 ) ;
  assign n8815 = ( x110 & n2567 ) | ( x110 & n8813 ) | ( n2567 & n8813 ) ;
  assign n8816 = n8813 | n8815 ;
  assign n8817 = x109 & ~n2562 ;
  assign n8818 = ( x108 & x109 ) | ( x108 & n8585 ) | ( x109 & n8585 ) ;
  assign n8819 = ( x109 & n8816 ) | ( x109 & ~n8817 ) | ( n8816 & ~n8817 ) ;
  assign n8820 = n8818 ^ x110 ^ x109 ;
  assign n8821 = n5020 & n8820 ;
  assign n8822 = n8814 | n8821 ;
  assign n8823 = n2565 & n8820 ;
  assign n8824 = n8819 | n8823 ;
  assign n8825 = n8824 ^ x35 ^ 1'b0 ;
  assign n8826 = n8825 ^ n8463 ^ n8412 ;
  assign n8827 = ( n8412 & n8463 ) | ( n8412 & n8825 ) | ( n8463 & n8825 ) ;
  assign n8828 = x108 & n4972 ;
  assign n8829 = ( x110 & n4985 ) | ( x110 & n8828 ) | ( n4985 & n8828 ) ;
  assign n8830 = n8828 | n8829 ;
  assign n8831 = n8822 ^ x17 ^ 1'b0 ;
  assign n8832 = x109 & ~n4980 ;
  assign n8833 = ( x109 & n8830 ) | ( x109 & ~n8832 ) | ( n8830 & ~n8832 ) ;
  assign n8834 = n4987 & n8820 ;
  assign n8835 = n8833 | n8834 ;
  assign n8836 = n8835 ^ x14 ^ 1'b0 ;
  assign n8837 = n8836 ^ n8783 ^ n8461 ;
  assign n8838 = ( n8461 & n8783 ) | ( n8461 & n8836 ) | ( n8783 & n8836 ) ;
  assign n8839 = x108 & n3344 ;
  assign n8840 = ( x110 & n3342 ) | ( x110 & n8839 ) | ( n3342 & n8839 ) ;
  assign n8841 = n8839 | n8840 ;
  assign n8842 = x109 & ~n3347 ;
  assign n8843 = ( x109 & n8841 ) | ( x109 & ~n8842 ) | ( n8841 & ~n8842 ) ;
  assign n8844 = n8831 ^ n8765 ^ n8545 ;
  assign n8845 = ( x109 & x110 ) | ( x109 & n8818 ) | ( x110 & n8818 ) ;
  assign n8846 = ( n8545 & n8765 ) | ( n8545 & n8831 ) | ( n8765 & n8831 ) ;
  assign n8847 = x108 & n3025 ;
  assign n8848 = ( x110 & n3015 ) | ( x110 & n8847 ) | ( n3015 & n8847 ) ;
  assign n8849 = n8847 | n8848 ;
  assign n8850 = x109 & ~n3014 ;
  assign n8851 = ( x109 & n8849 ) | ( x109 & ~n8850 ) | ( n8849 & ~n8850 ) ;
  assign n8852 = ( n3017 & n8820 ) | ( n3017 & n8851 ) | ( n8820 & n8851 ) ;
  assign n8853 = n8851 | n8852 ;
  assign n8854 = n8853 ^ x32 ^ 1'b0 ;
  assign n8855 = ( n8321 & n8606 ) | ( n8321 & n8854 ) | ( n8606 & n8854 ) ;
  assign n8856 = n8854 ^ n8606 ^ n8321 ;
  assign n8857 = x108 & n4616 ;
  assign n8858 = ( x110 & n4606 ) | ( x110 & n8857 ) | ( n4606 & n8857 ) ;
  assign n8859 = n8857 | n8858 ;
  assign n8860 = x109 & ~n4605 ;
  assign n8861 = ( x109 & n8859 ) | ( x109 & ~n8860 ) | ( n8859 & ~n8860 ) ;
  assign n8862 = n4608 & n8820 ;
  assign n8863 = n8861 | n8862 ;
  assign n8864 = ( n3346 & n8820 ) | ( n3346 & n8843 ) | ( n8820 & n8843 ) ;
  assign n8865 = n8843 | n8864 ;
  assign n8866 = n8865 ^ x29 ^ 1'b0 ;
  assign n8867 = n8866 ^ n8494 ^ n8312 ;
  assign n8868 = ( n8312 & n8494 ) | ( n8312 & n8866 ) | ( n8494 & n8866 ) ;
  assign n8869 = x108 & n3734 ;
  assign n8870 = ( x110 & n3732 ) | ( x110 & n8869 ) | ( n3732 & n8869 ) ;
  assign n8871 = n8869 | n8870 ;
  assign n8872 = x109 & ~n3737 ;
  assign n8873 = ( x109 & n8871 ) | ( x109 & ~n8872 ) | ( n8871 & ~n8872 ) ;
  assign n8874 = ( n3736 & n8820 ) | ( n3736 & n8873 ) | ( n8820 & n8873 ) ;
  assign n8875 = n8863 ^ x23 ^ 1'b0 ;
  assign n8876 = n8873 | n8874 ;
  assign n8877 = n8875 ^ n8535 ^ n8382 ;
  assign n8878 = n8876 ^ x26 ^ 1'b0 ;
  assign n8879 = ( n8382 & n8535 ) | ( n8382 & n8875 ) | ( n8535 & n8875 ) ;
  assign n8880 = ( n8372 & n8451 ) | ( n8372 & n8878 ) | ( n8451 & n8878 ) ;
  assign n8881 = n8878 ^ n8451 ^ n8372 ;
  assign n8882 = x108 & n5499 ;
  assign n8883 = ( x110 & n5497 ) | ( x110 & n8882 ) | ( n5497 & n8882 ) ;
  assign n8884 = n8882 | n8883 ;
  assign n8885 = x109 & ~n5502 ;
  assign n8886 = ( x109 & n8884 ) | ( x109 & ~n8885 ) | ( n8884 & ~n8885 ) ;
  assign n8887 = n5501 & n8820 ;
  assign n8888 = n8886 | n8887 ;
  assign n8889 = n8888 ^ x11 ^ 1'b0 ;
  assign n8890 = n8889 ^ n8801 ^ n8515 ;
  assign n8891 = ( n8515 & n8801 ) | ( n8515 & n8889 ) | ( n8801 & n8889 ) ;
  assign n8892 = x106 & n2156 ;
  assign n8893 = ( x108 & n2163 ) | ( x108 & n8892 ) | ( n2163 & n8892 ) ;
  assign n8894 = n8892 | n8893 ;
  assign n8895 = x107 & ~n2158 ;
  assign n8896 = ( x107 & n8894 ) | ( x107 & ~n8895 ) | ( n8894 & ~n8895 ) ;
  assign n8897 = n2161 & n8557 ;
  assign n8898 = n8896 | n8897 ;
  assign n8899 = n8898 ^ x38 ^ 1'b0 ;
  assign n8900 = ( n8110 & n8285 ) | ( n8110 & n8899 ) | ( n8285 & n8899 ) ;
  assign n8901 = n8899 ^ n8285 ^ n8110 ;
  assign n8902 = x108 & n5979 ;
  assign n8903 = ( x110 & n5969 ) | ( x110 & n8902 ) | ( n5969 & n8902 ) ;
  assign n8904 = n8902 | n8903 ;
  assign n8905 = x109 & ~n5970 ;
  assign n8906 = ( x109 & n8904 ) | ( x109 & ~n8905 ) | ( n8904 & ~n8905 ) ;
  assign n8907 = n5968 & n8820 ;
  assign n8908 = n8906 | n8907 ;
  assign n8909 = n8908 ^ x5 ^ 1'b0 ;
  assign n8910 = ( n8492 & n8776 ) | ( n8492 & n8909 ) | ( n8776 & n8909 ) ;
  assign n8911 = n8909 ^ n8776 ^ n8492 ;
  assign n8912 = x107 & n2156 ;
  assign n8913 = ( x109 & n2163 ) | ( x109 & n8912 ) | ( n2163 & n8912 ) ;
  assign n8914 = n8912 | n8913 ;
  assign n8915 = x108 & ~n2158 ;
  assign n8916 = ( x108 & n8914 ) | ( x108 & ~n8915 ) | ( n8914 & ~n8915 ) ;
  assign n8917 = n2161 & n8680 ;
  assign n8918 = n8916 | n8917 ;
  assign n8919 = n8918 ^ x38 ^ 1'b0 ;
  assign n8920 = n8919 ^ n8900 ^ n8291 ;
  assign n8921 = ( n8291 & n8900 ) | ( n8291 & n8919 ) | ( n8900 & n8919 ) ;
  assign n8922 = x108 & n6104 ;
  assign n8923 = ( x110 & n6105 ) | ( x110 & n8922 ) | ( n6105 & n8922 ) ;
  assign n8924 = n8922 | n8923 ;
  assign n8925 = x109 & ~n6107 ;
  assign n8926 = ( x109 & n8924 ) | ( x109 & ~n8925 ) | ( n8924 & ~n8925 ) ;
  assign n8927 = ~n6108 & n8820 ;
  assign n8928 = ( n8820 & n8926 ) | ( n8820 & ~n8927 ) | ( n8926 & ~n8927 ) ;
  assign n8929 = n8928 ^ x2 ^ 1'b0 ;
  assign n8930 = ( n8525 & n8701 ) | ( n8525 & n8929 ) | ( n8701 & n8929 ) ;
  assign n8931 = n8929 ^ n8701 ^ n8525 ;
  assign n8932 = x108 & n4790 ;
  assign n8933 = ( x110 & n4792 ) | ( x110 & n8932 ) | ( n4792 & n8932 ) ;
  assign n8934 = n8932 | n8933 ;
  assign n8935 = x109 & ~n4786 ;
  assign n8936 = ( x109 & n8934 ) | ( x109 & ~n8935 ) | ( n8934 & ~n8935 ) ;
  assign n8937 = n4787 & n8820 ;
  assign n8938 = n8936 | n8937 ;
  assign n8939 = n8938 ^ x20 ^ 1'b0 ;
  assign n8940 = n8939 ^ n8754 ^ n8505 ;
  assign n8941 = ( n8505 & n8754 ) | ( n8505 & n8939 ) | ( n8754 & n8939 ) ;
  assign n8942 = x109 & n4616 ;
  assign n8943 = ( x111 & n4606 ) | ( x111 & n8942 ) | ( n4606 & n8942 ) ;
  assign n8944 = n8942 | n8943 ;
  assign n8945 = x110 & ~n4605 ;
  assign n8946 = n8845 ^ x111 ^ x110 ;
  assign n8947 = ( x110 & n8944 ) | ( x110 & ~n8945 ) | ( n8944 & ~n8945 ) ;
  assign n8948 = n4608 & n8946 ;
  assign n8949 = n8947 | n8948 ;
  assign n8950 = n8949 ^ x23 ^ 1'b0 ;
  assign n8951 = n8950 ^ n8679 ^ n8534 ;
  assign n8952 = ( n8534 & n8679 ) | ( n8534 & n8950 ) | ( n8679 & n8950 ) ;
  assign n8953 = x109 & n2560 ;
  assign n8954 = ( x111 & n2567 ) | ( x111 & n8953 ) | ( n2567 & n8953 ) ;
  assign n8955 = n8953 | n8954 ;
  assign n8956 = x110 & ~n2562 ;
  assign n8957 = ( x110 & n8955 ) | ( x110 & ~n8956 ) | ( n8955 & ~n8956 ) ;
  assign n8958 = x108 & n5718 ;
  assign n8959 = n2565 & n8946 ;
  assign n8960 = n8957 | n8959 ;
  assign n8961 = ( x110 & n5720 ) | ( x110 & n8958 ) | ( n5720 & n8958 ) ;
  assign n8962 = n8958 | n8961 ;
  assign n8963 = x109 & ~n5727 ;
  assign n8964 = ( x109 & n8962 ) | ( x109 & ~n8963 ) | ( n8962 & ~n8963 ) ;
  assign n8965 = n5726 & n8820 ;
  assign n8966 = n8964 | n8965 ;
  assign n8967 = n8966 ^ x8 ^ 1'b0 ;
  assign n8968 = ( n8554 & n8807 ) | ( n8554 & n8967 ) | ( n8807 & n8967 ) ;
  assign n8969 = n8967 ^ n8807 ^ n8554 ;
  assign n8970 = x109 & n6104 ;
  assign n8971 = n8960 ^ x35 ^ 1'b0 ;
  assign n8972 = ( x111 & n6105 ) | ( x111 & n8970 ) | ( n6105 & n8970 ) ;
  assign n8973 = n8970 | n8972 ;
  assign n8974 = n8971 ^ n8901 ^ n8465 ;
  assign n8975 = ( n8465 & n8901 ) | ( n8465 & n8971 ) | ( n8901 & n8971 ) ;
  assign n8976 = x110 & ~n6107 ;
  assign n8977 = x109 & n3734 ;
  assign n8978 = ( x110 & n8973 ) | ( x110 & ~n8976 ) | ( n8973 & ~n8976 ) ;
  assign n8979 = ( x111 & n3732 ) | ( x111 & n8977 ) | ( n3732 & n8977 ) ;
  assign n8980 = n8977 | n8979 ;
  assign n8981 = ~n6108 & n8946 ;
  assign n8982 = ( n8946 & n8978 ) | ( n8946 & ~n8981 ) | ( n8978 & ~n8981 ) ;
  assign n8983 = n8982 ^ x2 ^ 1'b0 ;
  assign n8984 = x110 & ~n3737 ;
  assign n8985 = ( x110 & n8980 ) | ( x110 & ~n8984 ) | ( n8980 & ~n8984 ) ;
  assign n8986 = n8983 ^ n8930 ^ n8637 ;
  assign n8987 = ( n8637 & n8930 ) | ( n8637 & n8983 ) | ( n8930 & n8983 ) ;
  assign n8988 = n3736 & n8946 ;
  assign n8989 = x109 & n3025 ;
  assign n8990 = n8985 | n8988 ;
  assign n8991 = ( x111 & n3015 ) | ( x111 & n8989 ) | ( n3015 & n8989 ) ;
  assign n8992 = n8989 | n8991 ;
  assign n8993 = n8990 ^ x26 ^ 1'b0 ;
  assign n8994 = n8993 ^ n8735 ^ n8450 ;
  assign n8995 = ( n8450 & n8735 ) | ( n8450 & n8993 ) | ( n8735 & n8993 ) ;
  assign n8996 = x110 & ~n3014 ;
  assign n8997 = ( x110 & n8992 ) | ( x110 & ~n8996 ) | ( n8992 & ~n8996 ) ;
  assign n8998 = ( n3017 & n8946 ) | ( n3017 & n8997 ) | ( n8946 & n8997 ) ;
  assign n8999 = n8997 | n8998 ;
  assign n9000 = n8999 ^ x32 ^ 1'b0 ;
  assign n9001 = ( n8587 & n8607 ) | ( n8587 & n9000 ) | ( n8607 & n9000 ) ;
  assign n9002 = n9000 ^ n8607 ^ n8587 ;
  assign n9003 = ( x110 & x111 ) | ( x110 & n8845 ) | ( x111 & n8845 ) ;
  assign n9004 = x109 & n4790 ;
  assign n9005 = ( x111 & n4792 ) | ( x111 & n9004 ) | ( n4792 & n9004 ) ;
  assign n9006 = x110 & ~n4786 ;
  assign n9007 = n9004 | n9005 ;
  assign n9008 = ( x110 & ~n9006 ) | ( x110 & n9007 ) | ( ~n9006 & n9007 ) ;
  assign n9009 = x109 & n5979 ;
  assign n9010 = ( x111 & n5969 ) | ( x111 & n9009 ) | ( n5969 & n9009 ) ;
  assign n9011 = n9009 | n9010 ;
  assign n9012 = x110 & ~n5970 ;
  assign n9013 = ( x110 & n9011 ) | ( x110 & ~n9012 ) | ( n9011 & ~n9012 ) ;
  assign n9014 = n5968 & n8946 ;
  assign n9015 = n9013 | n9014 ;
  assign n9016 = n4787 & n8946 ;
  assign n9017 = n9008 | n9016 ;
  assign n9018 = n9017 ^ x20 ^ 1'b0 ;
  assign n9019 = ( n8565 & n8941 ) | ( n8565 & n9018 ) | ( n8941 & n9018 ) ;
  assign n9020 = n9018 ^ n8941 ^ n8565 ;
  assign n9021 = x109 & n5011 ;
  assign n9022 = ( x111 & n5012 ) | ( x111 & n9021 ) | ( n5012 & n9021 ) ;
  assign n9023 = n9021 | n9022 ;
  assign n9024 = x110 & ~n5008 ;
  assign n9025 = ( x110 & n9023 ) | ( x110 & ~n9024 ) | ( n9023 & ~n9024 ) ;
  assign n9026 = n5020 & n8946 ;
  assign n9027 = n9025 | n9026 ;
  assign n9028 = n9027 ^ x17 ^ 1'b0 ;
  assign n9029 = n9028 ^ n8846 ^ n8647 ;
  assign n9030 = ( n8647 & n8846 ) | ( n8647 & n9028 ) | ( n8846 & n9028 ) ;
  assign n9031 = x109 & n4972 ;
  assign n9032 = ( x111 & n4985 ) | ( x111 & n9031 ) | ( n4985 & n9031 ) ;
  assign n9033 = n9031 | n9032 ;
  assign n9034 = x110 & ~n4980 ;
  assign n9035 = ( x110 & n9033 ) | ( x110 & ~n9034 ) | ( n9033 & ~n9034 ) ;
  assign n9036 = n4987 & n8946 ;
  assign n9037 = n9035 | n9036 ;
  assign n9038 = n9037 ^ x14 ^ 1'b0 ;
  assign n9039 = n9015 ^ x5 ^ 1'b0 ;
  assign n9040 = n9039 ^ n8910 ^ n8666 ;
  assign n9041 = ( n8666 & n8910 ) | ( n8666 & n9039 ) | ( n8910 & n9039 ) ;
  assign n9042 = x109 & n3344 ;
  assign n9043 = ( x111 & n3342 ) | ( x111 & n9042 ) | ( n3342 & n9042 ) ;
  assign n9044 = n9042 | n9043 ;
  assign n9045 = x110 & ~n3347 ;
  assign n9046 = ( x110 & n9044 ) | ( x110 & ~n9045 ) | ( n9044 & ~n9045 ) ;
  assign n9047 = n9038 ^ n8838 ^ n8617 ;
  assign n9048 = ( n8617 & n8838 ) | ( n8617 & n9038 ) | ( n8838 & n9038 ) ;
  assign n9049 = x109 & n5499 ;
  assign n9050 = ( x111 & n5497 ) | ( x111 & n9049 ) | ( n5497 & n9049 ) ;
  assign n9051 = n9049 | n9050 ;
  assign n9052 = x110 & ~n5502 ;
  assign n9053 = ( x110 & n9051 ) | ( x110 & ~n9052 ) | ( n9051 & ~n9052 ) ;
  assign n9054 = n5501 & n8946 ;
  assign n9055 = n9053 | n9054 ;
  assign n9056 = n3346 & n8946 ;
  assign n9057 = n9046 | n9056 ;
  assign n9058 = n9055 ^ x11 ^ 1'b0 ;
  assign n9059 = n9057 ^ x29 ^ 1'b0 ;
  assign n9060 = ( n8495 & n8596 ) | ( n8495 & n9059 ) | ( n8596 & n9059 ) ;
  assign n9061 = n9059 ^ n8596 ^ n8495 ;
  assign n9062 = x109 & n5718 ;
  assign n9063 = ( x111 & n5720 ) | ( x111 & n9062 ) | ( n5720 & n9062 ) ;
  assign n9064 = n9062 | n9063 ;
  assign n9065 = n9058 ^ n8891 ^ n8657 ;
  assign n9066 = ( n8657 & n8891 ) | ( n8657 & n9058 ) | ( n8891 & n9058 ) ;
  assign n9067 = x110 & ~n5727 ;
  assign n9068 = n5726 & n8946 ;
  assign n9069 = ( x110 & n9064 ) | ( x110 & ~n9067 ) | ( n9064 & ~n9067 ) ;
  assign n9070 = n9068 | n9069 ;
  assign n9071 = n9070 ^ x8 ^ 1'b0 ;
  assign n9072 = ( n8627 & n8968 ) | ( n8627 & n9071 ) | ( n8968 & n9071 ) ;
  assign n9073 = n9071 ^ n8968 ^ n8627 ;
  assign n9074 = x110 & n2560 ;
  assign n9075 = ( x112 & n2567 ) | ( x112 & n9074 ) | ( n2567 & n9074 ) ;
  assign n9076 = x110 & n3344 ;
  assign n9077 = ( x112 & n3342 ) | ( x112 & n9076 ) | ( n3342 & n9076 ) ;
  assign n9078 = n9074 | n9075 ;
  assign n9079 = n9076 | n9077 ;
  assign n9080 = n9003 ^ x112 ^ x111 ;
  assign n9081 = x111 & ~n2562 ;
  assign n9082 = ( x111 & n9078 ) | ( x111 & ~n9081 ) | ( n9078 & ~n9081 ) ;
  assign n9083 = x111 & ~n3347 ;
  assign n9084 = ( x111 & n9079 ) | ( x111 & ~n9083 ) | ( n9079 & ~n9083 ) ;
  assign n9085 = n2565 & n9080 ;
  assign n9086 = n9082 | n9085 ;
  assign n9087 = n3346 & n9080 ;
  assign n9088 = n9084 | n9087 ;
  assign n9089 = n9088 ^ x29 ^ 1'b0 ;
  assign n9090 = ( n8722 & n9060 ) | ( n8722 & n9089 ) | ( n9060 & n9089 ) ;
  assign n9091 = n9089 ^ n9060 ^ n8722 ;
  assign n9092 = x110 & n5011 ;
  assign n9093 = ( x112 & n5012 ) | ( x112 & n9092 ) | ( n5012 & n9092 ) ;
  assign n9094 = n9092 | n9093 ;
  assign n9095 = x111 & ~n5008 ;
  assign n9096 = ( x111 & n9094 ) | ( x111 & ~n9095 ) | ( n9094 & ~n9095 ) ;
  assign n9097 = n5020 & n9080 ;
  assign n9098 = n9096 | n9097 ;
  assign n9099 = n9098 ^ x17 ^ 1'b0 ;
  assign n9100 = n9086 ^ x35 ^ 1'b0 ;
  assign n9101 = n9099 ^ n9030 ^ n8755 ;
  assign n9102 = ( n8755 & n9030 ) | ( n8755 & n9099 ) | ( n9030 & n9099 ) ;
  assign n9103 = n9100 ^ n8975 ^ n8920 ;
  assign n9104 = x110 & n6104 ;
  assign n9105 = ( n8920 & n8975 ) | ( n8920 & n9100 ) | ( n8975 & n9100 ) ;
  assign n9106 = ( x112 & n6105 ) | ( x112 & n9104 ) | ( n6105 & n9104 ) ;
  assign n9107 = n9104 | n9106 ;
  assign n9108 = ( x111 & x112 ) | ( x111 & n9003 ) | ( x112 & n9003 ) ;
  assign n9109 = x111 & ~n6107 ;
  assign n9110 = ( x111 & n9107 ) | ( x111 & ~n9109 ) | ( n9107 & ~n9109 ) ;
  assign n9111 = ~n6108 & n9080 ;
  assign n9112 = ( n9080 & n9110 ) | ( n9080 & ~n9111 ) | ( n9110 & ~n9111 ) ;
  assign n9113 = n9112 ^ x2 ^ 1'b0 ;
  assign n9114 = ( n8775 & n8987 ) | ( n8775 & n9113 ) | ( n8987 & n9113 ) ;
  assign n9115 = n9113 ^ n8987 ^ n8775 ;
  assign n9116 = x110 & n5718 ;
  assign n9117 = ( x112 & n5720 ) | ( x112 & n9116 ) | ( n5720 & n9116 ) ;
  assign n9118 = x111 & ~n5727 ;
  assign n9119 = n9116 | n9117 ;
  assign n9120 = x110 & n3025 ;
  assign n9121 = ( x111 & ~n9118 ) | ( x111 & n9119 ) | ( ~n9118 & n9119 ) ;
  assign n9122 = n5726 & n9080 ;
  assign n9123 = n9121 | n9122 ;
  assign n9124 = ( x112 & n3015 ) | ( x112 & n9120 ) | ( n3015 & n9120 ) ;
  assign n9125 = n9120 | n9124 ;
  assign n9126 = x111 & ~n3014 ;
  assign n9127 = ( x111 & n9125 ) | ( x111 & ~n9126 ) | ( n9125 & ~n9126 ) ;
  assign n9128 = n9123 ^ x8 ^ 1'b0 ;
  assign n9129 = n3017 & n9080 ;
  assign n9130 = n9127 | n9129 ;
  assign n9131 = n9130 ^ x32 ^ 1'b0 ;
  assign n9132 = n9128 ^ n9072 ^ n8800 ;
  assign n9133 = ( n8800 & n9072 ) | ( n8800 & n9128 ) | ( n9072 & n9128 ) ;
  assign n9134 = n9131 ^ n9001 ^ n8696 ;
  assign n9135 = ( n8696 & n9001 ) | ( n8696 & n9131 ) | ( n9001 & n9131 ) ;
  assign n9136 = x110 & n4616 ;
  assign n9137 = ( x112 & n4606 ) | ( x112 & n9136 ) | ( n4606 & n9136 ) ;
  assign n9138 = n9136 | n9137 ;
  assign n9139 = x111 & ~n4605 ;
  assign n9140 = ( x111 & n9138 ) | ( x111 & ~n9139 ) | ( n9138 & ~n9139 ) ;
  assign n9141 = n4608 & n9080 ;
  assign n9142 = n9140 | n9141 ;
  assign n9143 = n9142 ^ x23 ^ 1'b0 ;
  assign n9144 = ( n8738 & n8952 ) | ( n8738 & n9143 ) | ( n8952 & n9143 ) ;
  assign n9145 = n9143 ^ n8952 ^ n8738 ;
  assign n9146 = x110 & n4972 ;
  assign n9147 = ( x112 & n4985 ) | ( x112 & n9146 ) | ( n4985 & n9146 ) ;
  assign n9148 = n9146 | n9147 ;
  assign n9149 = x111 & ~n4980 ;
  assign n9150 = ( x111 & n9148 ) | ( x111 & ~n9149 ) | ( n9148 & ~n9149 ) ;
  assign n9151 = n4987 & n9080 ;
  assign n9152 = n9150 | n9151 ;
  assign n9153 = n9152 ^ x14 ^ 1'b0 ;
  assign n9154 = ( n8764 & n9048 ) | ( n8764 & n9153 ) | ( n9048 & n9153 ) ;
  assign n9155 = n9153 ^ n9048 ^ n8764 ;
  assign n9156 = x110 & n5979 ;
  assign n9157 = ( x112 & n5969 ) | ( x112 & n9156 ) | ( n5969 & n9156 ) ;
  assign n9158 = n9156 | n9157 ;
  assign n9159 = x111 & ~n5970 ;
  assign n9160 = ( x111 & n9158 ) | ( x111 & ~n9159 ) | ( n9158 & ~n9159 ) ;
  assign n9161 = n5968 & n9080 ;
  assign n9162 = n9160 | n9161 ;
  assign n9163 = n9162 ^ x5 ^ 1'b0 ;
  assign n9164 = ( n8808 & n9041 ) | ( n8808 & n9163 ) | ( n9041 & n9163 ) ;
  assign n9165 = n9163 ^ n9041 ^ n8808 ;
  assign n9166 = x110 & n3734 ;
  assign n9167 = ( x112 & n3732 ) | ( x112 & n9166 ) | ( n3732 & n9166 ) ;
  assign n9168 = n9166 | n9167 ;
  assign n9169 = x111 & ~n3737 ;
  assign n9170 = ( x111 & n9168 ) | ( x111 & ~n9169 ) | ( n9168 & ~n9169 ) ;
  assign n9171 = n3736 & n9080 ;
  assign n9172 = n9170 | n9171 ;
  assign n9173 = n9172 ^ x26 ^ 1'b0 ;
  assign n9174 = ( n8796 & n8995 ) | ( n8796 & n9173 ) | ( n8995 & n9173 ) ;
  assign n9175 = n9173 ^ n8995 ^ n8796 ;
  assign n9176 = x110 & n4790 ;
  assign n9177 = ( x112 & n4792 ) | ( x112 & n9176 ) | ( n4792 & n9176 ) ;
  assign n9178 = n9176 | n9177 ;
  assign n9179 = x111 & ~n4786 ;
  assign n9180 = ( x111 & n9178 ) | ( x111 & ~n9179 ) | ( n9178 & ~n9179 ) ;
  assign n9181 = n4787 & n9080 ;
  assign n9182 = n9180 | n9181 ;
  assign n9183 = n9182 ^ x20 ^ 1'b0 ;
  assign n9184 = ( n8566 & n8710 ) | ( n8566 & n9183 ) | ( n8710 & n9183 ) ;
  assign n9185 = n9183 ^ n8710 ^ n8566 ;
  assign n9186 = x110 & n5499 ;
  assign n9187 = ( x112 & n5497 ) | ( x112 & n9186 ) | ( n5497 & n9186 ) ;
  assign n9188 = n9186 | n9187 ;
  assign n9189 = x111 & ~n5502 ;
  assign n9190 = ( x111 & n9188 ) | ( x111 & ~n9189 ) | ( n9188 & ~n9189 ) ;
  assign n9191 = n5501 & n9080 ;
  assign n9192 = n9190 | n9191 ;
  assign n9193 = n9192 ^ x11 ^ 1'b0 ;
  assign n9194 = n9193 ^ n9066 ^ n8782 ;
  assign n9195 = ( n8782 & n9066 ) | ( n8782 & n9193 ) | ( n9066 & n9193 ) ;
  assign n9196 = x111 & n5011 ;
  assign n9197 = ( x113 & n5012 ) | ( x113 & n9196 ) | ( n5012 & n9196 ) ;
  assign n9198 = n9196 | n9197 ;
  assign n9199 = n9108 ^ x113 ^ x112 ;
  assign n9200 = x112 & ~n5008 ;
  assign n9201 = ( x112 & n9198 ) | ( x112 & ~n9200 ) | ( n9198 & ~n9200 ) ;
  assign n9202 = n5020 & n9199 ;
  assign n9203 = n9201 | n9202 ;
  assign n9204 = n9203 ^ x17 ^ 1'b0 ;
  assign n9205 = n9204 ^ n9102 ^ n8940 ;
  assign n9206 = ( n8940 & n9102 ) | ( n8940 & n9204 ) | ( n9102 & n9204 ) ;
  assign n9207 = x111 & n6104 ;
  assign n9208 = ( x113 & n6105 ) | ( x113 & n9207 ) | ( n6105 & n9207 ) ;
  assign n9209 = n9207 | n9208 ;
  assign n9210 = x112 & ~n6107 ;
  assign n9211 = ( x112 & n9209 ) | ( x112 & ~n9210 ) | ( n9209 & ~n9210 ) ;
  assign n9212 = ~n6108 & n9199 ;
  assign n9213 = ( n9199 & n9211 ) | ( n9199 & ~n9212 ) | ( n9211 & ~n9212 ) ;
  assign n9214 = n9213 ^ x2 ^ 1'b0 ;
  assign n9215 = ( n8911 & n9114 ) | ( n8911 & n9214 ) | ( n9114 & n9214 ) ;
  assign n9216 = n9214 ^ n9114 ^ n8911 ;
  assign n9217 = x111 & n5718 ;
  assign n9218 = ( x113 & n5720 ) | ( x113 & n9217 ) | ( n5720 & n9217 ) ;
  assign n9219 = n9217 | n9218 ;
  assign n9220 = x112 & ~n5727 ;
  assign n9221 = ( x112 & n9219 ) | ( x112 & ~n9220 ) | ( n9219 & ~n9220 ) ;
  assign n9222 = n5726 & n9199 ;
  assign n9223 = n9221 | n9222 ;
  assign n9224 = n9223 ^ x8 ^ 1'b0 ;
  assign n9225 = ( n8890 & n9133 ) | ( n8890 & n9224 ) | ( n9133 & n9224 ) ;
  assign n9226 = n9224 ^ n9133 ^ n8890 ;
  assign n9227 = x111 & n5979 ;
  assign n9228 = ( x113 & n5969 ) | ( x113 & n9227 ) | ( n5969 & n9227 ) ;
  assign n9229 = n9227 | n9228 ;
  assign n9230 = x112 & ~n5970 ;
  assign n9231 = ( x112 & n9229 ) | ( x112 & ~n9230 ) | ( n9229 & ~n9230 ) ;
  assign n9232 = n5968 & n9199 ;
  assign n9233 = n9231 | n9232 ;
  assign n9234 = n9233 ^ x5 ^ 1'b0 ;
  assign n9235 = ( n8969 & n9164 ) | ( n8969 & n9234 ) | ( n9164 & n9234 ) ;
  assign n9236 = n9234 ^ n9164 ^ n8969 ;
  assign n9237 = x111 & n4790 ;
  assign n9238 = ( x113 & n4792 ) | ( x113 & n9237 ) | ( n4792 & n9237 ) ;
  assign n9239 = n9237 | n9238 ;
  assign n9240 = x112 & ~n4786 ;
  assign n9241 = ( x112 & n9239 ) | ( x112 & ~n9240 ) | ( n9239 & ~n9240 ) ;
  assign n9242 = n4787 & n9199 ;
  assign n9243 = n9241 | n9242 ;
  assign n9244 = n9243 ^ x20 ^ 1'b0 ;
  assign n9245 = n9244 ^ n8877 ^ n8711 ;
  assign n9246 = ( n8711 & n8877 ) | ( n8711 & n9244 ) | ( n8877 & n9244 ) ;
  assign n9247 = x111 & n4972 ;
  assign n9248 = ( x113 & n4985 ) | ( x113 & n9247 ) | ( n4985 & n9247 ) ;
  assign n9249 = n9247 | n9248 ;
  assign n9250 = x112 & ~n4980 ;
  assign n9251 = ( x112 & n9249 ) | ( x112 & ~n9250 ) | ( n9249 & ~n9250 ) ;
  assign n9252 = n4987 & n9199 ;
  assign n9253 = n9251 | n9252 ;
  assign n9254 = n9253 ^ x14 ^ 1'b0 ;
  assign n9255 = n9254 ^ n9154 ^ n8844 ;
  assign n9256 = ( n8844 & n9154 ) | ( n8844 & n9254 ) | ( n9154 & n9254 ) ;
  assign n9257 = x111 & n5499 ;
  assign n9258 = ( x113 & n5497 ) | ( x113 & n9257 ) | ( n5497 & n9257 ) ;
  assign n9259 = n9257 | n9258 ;
  assign n9260 = ( x112 & x113 ) | ( x112 & n9108 ) | ( x113 & n9108 ) ;
  assign n9261 = x112 & ~n5502 ;
  assign n9262 = ( x112 & n9259 ) | ( x112 & ~n9261 ) | ( n9259 & ~n9261 ) ;
  assign n9263 = n5501 & n9199 ;
  assign n9264 = n9262 | n9263 ;
  assign n9265 = n9264 ^ x11 ^ 1'b0 ;
  assign n9266 = ( n8837 & n9195 ) | ( n8837 & n9265 ) | ( n9195 & n9265 ) ;
  assign n9267 = n9265 ^ n9195 ^ n8837 ;
  assign n9268 = x111 & n3344 ;
  assign n9269 = ( x113 & n3342 ) | ( x113 & n9268 ) | ( n3342 & n9268 ) ;
  assign n9270 = n9268 | n9269 ;
  assign n9271 = x112 & ~n3347 ;
  assign n9272 = ( x112 & n9270 ) | ( x112 & ~n9271 ) | ( n9270 & ~n9271 ) ;
  assign n9273 = n3346 & n9199 ;
  assign n9274 = x112 & n5499 ;
  assign n9275 = n9272 | n9273 ;
  assign n9276 = n9275 ^ x29 ^ 1'b0 ;
  assign n9277 = ( n8723 & n8856 ) | ( n8723 & n9276 ) | ( n8856 & n9276 ) ;
  assign n9278 = n9276 ^ n8856 ^ n8723 ;
  assign n9279 = n9260 ^ x114 ^ x113 ;
  assign n9280 = ( x114 & n5497 ) | ( x114 & n9274 ) | ( n5497 & n9274 ) ;
  assign n9281 = n9274 | n9280 ;
  assign n9282 = ( x113 & x114 ) | ( x113 & n9260 ) | ( x114 & n9260 ) ;
  assign n9283 = x113 & ~n5502 ;
  assign n9284 = ( x113 & n9281 ) | ( x113 & ~n9283 ) | ( n9281 & ~n9283 ) ;
  assign n9285 = n5501 & n9279 ;
  assign n9286 = n9284 | n9285 ;
  assign n9287 = n9286 ^ x11 ^ 1'b0 ;
  assign n9288 = n9287 ^ n9266 ^ n9047 ;
  assign n9289 = ( n9047 & n9266 ) | ( n9047 & n9287 ) | ( n9266 & n9287 ) ;
  assign n9290 = x111 & n4616 ;
  assign n9291 = ( x113 & n4606 ) | ( x113 & n9290 ) | ( n4606 & n9290 ) ;
  assign n9292 = n9290 | n9291 ;
  assign n9293 = x112 & ~n4605 ;
  assign n9294 = ( x112 & n9292 ) | ( x112 & ~n9293 ) | ( n9292 & ~n9293 ) ;
  assign n9295 = n4608 & n9199 ;
  assign n9296 = n9294 | n9295 ;
  assign n9297 = n9296 ^ x23 ^ 1'b0 ;
  assign n9298 = ( n8737 & n8881 ) | ( n8737 & n9297 ) | ( n8881 & n9297 ) ;
  assign n9299 = n9297 ^ n8881 ^ n8737 ;
  assign n9300 = x112 & n5011 ;
  assign n9301 = ( x114 & n5012 ) | ( x114 & n9300 ) | ( n5012 & n9300 ) ;
  assign n9302 = n9300 | n9301 ;
  assign n9303 = x113 & ~n5008 ;
  assign n9304 = ( x113 & n9302 ) | ( x113 & ~n9303 ) | ( n9302 & ~n9303 ) ;
  assign n9305 = n5020 & n9279 ;
  assign n9306 = n9304 | n9305 ;
  assign n9307 = n9306 ^ x17 ^ 1'b0 ;
  assign n9308 = ( n9020 & n9206 ) | ( n9020 & n9307 ) | ( n9206 & n9307 ) ;
  assign n9309 = n9307 ^ n9206 ^ n9020 ;
  assign n9310 = x111 & n3734 ;
  assign n9311 = ( x113 & n3732 ) | ( x113 & n9310 ) | ( n3732 & n9310 ) ;
  assign n9312 = n9310 | n9311 ;
  assign n9313 = x112 & ~n3737 ;
  assign n9314 = ( x112 & n9312 ) | ( x112 & ~n9313 ) | ( n9312 & ~n9313 ) ;
  assign n9315 = n3736 & n9199 ;
  assign n9316 = n9314 | n9315 ;
  assign n9317 = n9316 ^ x26 ^ 1'b0 ;
  assign n9318 = n9317 ^ n8867 ^ n8795 ;
  assign n9319 = ( n8795 & n8867 ) | ( n8795 & n9317 ) | ( n8867 & n9317 ) ;
  assign n9320 = x111 & n3025 ;
  assign n9321 = ( x113 & n3015 ) | ( x113 & n9320 ) | ( n3015 & n9320 ) ;
  assign n9322 = n9320 | n9321 ;
  assign n9323 = x112 & ~n3014 ;
  assign n9324 = ( x112 & n9322 ) | ( x112 & ~n9323 ) | ( n9322 & ~n9323 ) ;
  assign n9325 = n3017 & n9199 ;
  assign n9326 = n9324 | n9325 ;
  assign n9327 = n9326 ^ x32 ^ 1'b0 ;
  assign n9328 = n9327 ^ n8826 ^ n8695 ;
  assign n9329 = ( n8695 & n8826 ) | ( n8695 & n9327 ) | ( n8826 & n9327 ) ;
  assign n9330 = x112 & n3344 ;
  assign n9331 = ( x114 & n3342 ) | ( x114 & n9330 ) | ( n3342 & n9330 ) ;
  assign n9332 = n9330 | n9331 ;
  assign n9333 = x113 & ~n3347 ;
  assign n9334 = ( x113 & n9332 ) | ( x113 & ~n9333 ) | ( n9332 & ~n9333 ) ;
  assign n9335 = ( n3346 & n9279 ) | ( n3346 & n9334 ) | ( n9279 & n9334 ) ;
  assign n9336 = n9334 | n9335 ;
  assign n9337 = n9336 ^ x29 ^ 1'b0 ;
  assign n9338 = ( n8855 & n9002 ) | ( n8855 & n9337 ) | ( n9002 & n9337 ) ;
  assign n9339 = n9337 ^ n9002 ^ n8855 ;
  assign n9340 = x112 & n5979 ;
  assign n9341 = x112 & n4790 ;
  assign n9342 = ( x114 & n4792 ) | ( x114 & n9341 ) | ( n4792 & n9341 ) ;
  assign n9343 = n9341 | n9342 ;
  assign n9344 = ( x114 & n5969 ) | ( x114 & n9340 ) | ( n5969 & n9340 ) ;
  assign n9345 = n9340 | n9344 ;
  assign n9346 = x113 & ~n5970 ;
  assign n9347 = ( x113 & n9345 ) | ( x113 & ~n9346 ) | ( n9345 & ~n9346 ) ;
  assign n9348 = n5968 & n9279 ;
  assign n9349 = n9347 | n9348 ;
  assign n9350 = x113 & ~n4786 ;
  assign n9351 = ( x113 & n9343 ) | ( x113 & ~n9350 ) | ( n9343 & ~n9350 ) ;
  assign n9352 = n4787 & n9279 ;
  assign n9353 = n9351 | n9352 ;
  assign n9354 = n9349 ^ x5 ^ 1'b0 ;
  assign n9355 = n9353 ^ x20 ^ 1'b0 ;
  assign n9356 = ( n8879 & n8951 ) | ( n8879 & n9355 ) | ( n8951 & n9355 ) ;
  assign n9357 = n9355 ^ n8951 ^ n8879 ;
  assign n9358 = n9354 ^ n9235 ^ n9073 ;
  assign n9359 = ( n9073 & n9235 ) | ( n9073 & n9354 ) | ( n9235 & n9354 ) ;
  assign n9360 = x113 & ~n5727 ;
  assign n9361 = x112 & n5718 ;
  assign n9362 = ( x114 & n5720 ) | ( x114 & n9361 ) | ( n5720 & n9361 ) ;
  assign n9363 = n9361 | n9362 ;
  assign n9364 = ( x113 & ~n9360 ) | ( x113 & n9363 ) | ( ~n9360 & n9363 ) ;
  assign n9365 = n5726 & n9279 ;
  assign n9366 = n9364 | n9365 ;
  assign n9367 = n9366 ^ x8 ^ 1'b0 ;
  assign n9368 = n9367 ^ n9225 ^ n9065 ;
  assign n9369 = x112 & n3734 ;
  assign n9370 = ( n9065 & n9225 ) | ( n9065 & n9367 ) | ( n9225 & n9367 ) ;
  assign n9371 = ( x114 & n3732 ) | ( x114 & n9369 ) | ( n3732 & n9369 ) ;
  assign n9372 = n9369 | n9371 ;
  assign n9373 = x113 & ~n3737 ;
  assign n9374 = ( x113 & n9372 ) | ( x113 & ~n9373 ) | ( n9372 & ~n9373 ) ;
  assign n9375 = ( n3736 & n9279 ) | ( n3736 & n9374 ) | ( n9279 & n9374 ) ;
  assign n9376 = n9374 | n9375 ;
  assign n9377 = n9376 ^ x26 ^ 1'b0 ;
  assign n9378 = n9377 ^ n9061 ^ n8868 ;
  assign n9379 = ( n8868 & n9061 ) | ( n8868 & n9377 ) | ( n9061 & n9377 ) ;
  assign n9380 = n4987 & n9279 ;
  assign n9381 = x112 & n4972 ;
  assign n9382 = ( x114 & n4985 ) | ( x114 & n9381 ) | ( n4985 & n9381 ) ;
  assign n9383 = n9381 | n9382 ;
  assign n9384 = x113 & ~n4980 ;
  assign n9385 = ( x113 & n9383 ) | ( x113 & ~n9384 ) | ( n9383 & ~n9384 ) ;
  assign n9386 = x112 & n3025 ;
  assign n9387 = n9380 | n9385 ;
  assign n9388 = n9387 ^ x14 ^ 1'b0 ;
  assign n9389 = ( x114 & n3015 ) | ( x114 & n9386 ) | ( n3015 & n9386 ) ;
  assign n9390 = n9386 | n9389 ;
  assign n9391 = x113 & ~n3014 ;
  assign n9392 = ( x113 & n9390 ) | ( x113 & ~n9391 ) | ( n9390 & ~n9391 ) ;
  assign n9393 = ( n9029 & n9256 ) | ( n9029 & n9388 ) | ( n9256 & n9388 ) ;
  assign n9394 = n9388 ^ n9256 ^ n9029 ;
  assign n9395 = n4608 & n9279 ;
  assign n9396 = n3017 & n9279 ;
  assign n9397 = n9392 | n9396 ;
  assign n9398 = n9397 ^ x32 ^ 1'b0 ;
  assign n9399 = ( n8827 & n8974 ) | ( n8827 & n9398 ) | ( n8974 & n9398 ) ;
  assign n9400 = n9398 ^ n8974 ^ n8827 ;
  assign n9401 = x112 & n4616 ;
  assign n9402 = ( x114 & n4606 ) | ( x114 & n9401 ) | ( n4606 & n9401 ) ;
  assign n9403 = n9401 | n9402 ;
  assign n9404 = x113 & ~n4605 ;
  assign n9405 = ( x113 & n9403 ) | ( x113 & ~n9404 ) | ( n9403 & ~n9404 ) ;
  assign n9406 = n9395 | n9405 ;
  assign n9407 = n9406 ^ x23 ^ 1'b0 ;
  assign n9408 = ( n8880 & n8994 ) | ( n8880 & n9407 ) | ( n8994 & n9407 ) ;
  assign n9409 = n9407 ^ n8994 ^ n8880 ;
  assign n9410 = x114 & ~n3347 ;
  assign n9411 = x113 & n3344 ;
  assign n9412 = ( x115 & n3342 ) | ( x115 & n9411 ) | ( n3342 & n9411 ) ;
  assign n9413 = n9411 | n9412 ;
  assign n9414 = n9282 ^ x115 ^ x114 ;
  assign n9415 = ( x114 & ~n9410 ) | ( x114 & n9413 ) | ( ~n9410 & n9413 ) ;
  assign n9416 = n3346 & n9414 ;
  assign n9417 = n9415 | n9416 ;
  assign n9418 = n9417 ^ x29 ^ 1'b0 ;
  assign n9419 = ( n9134 & n9338 ) | ( n9134 & n9418 ) | ( n9338 & n9418 ) ;
  assign n9420 = n9418 ^ n9338 ^ n9134 ;
  assign n9421 = x113 & n3025 ;
  assign n9422 = ( x115 & n3015 ) | ( x115 & n9421 ) | ( n3015 & n9421 ) ;
  assign n9423 = ( x114 & x115 ) | ( x114 & n9282 ) | ( x115 & n9282 ) ;
  assign n9424 = n9421 | n9422 ;
  assign n9425 = x114 & ~n3014 ;
  assign n9426 = ( x114 & n9424 ) | ( x114 & ~n9425 ) | ( n9424 & ~n9425 ) ;
  assign n9427 = n3017 & n9414 ;
  assign n9428 = n9426 | n9427 ;
  assign n9429 = n9428 ^ x32 ^ 1'b0 ;
  assign n9430 = ( n9103 & n9399 ) | ( n9103 & n9429 ) | ( n9399 & n9429 ) ;
  assign n9431 = n9429 ^ n9399 ^ n9103 ;
  assign n9432 = x113 & n4616 ;
  assign n9433 = ( x115 & n4606 ) | ( x115 & n9432 ) | ( n4606 & n9432 ) ;
  assign n9434 = n9432 | n9433 ;
  assign n9435 = x114 & ~n4605 ;
  assign n9436 = ( x114 & n9434 ) | ( x114 & ~n9435 ) | ( n9434 & ~n9435 ) ;
  assign n9437 = n4608 & n9414 ;
  assign n9438 = n9436 | n9437 ;
  assign n9439 = n9438 ^ x23 ^ 1'b0 ;
  assign n9440 = ( n9175 & n9408 ) | ( n9175 & n9439 ) | ( n9408 & n9439 ) ;
  assign n9441 = n9439 ^ n9408 ^ n9175 ;
  assign n9442 = x113 & n3734 ;
  assign n9443 = ( x115 & n3732 ) | ( x115 & n9442 ) | ( n3732 & n9442 ) ;
  assign n9444 = n9442 | n9443 ;
  assign n9445 = x114 & ~n3737 ;
  assign n9446 = ( x114 & n9444 ) | ( x114 & ~n9445 ) | ( n9444 & ~n9445 ) ;
  assign n9447 = n3736 & n9414 ;
  assign n9448 = n9446 | n9447 ;
  assign n9449 = n9448 ^ x26 ^ 1'b0 ;
  assign n9450 = n9449 ^ n9379 ^ n9091 ;
  assign n9451 = ( n9091 & n9379 ) | ( n9091 & n9449 ) | ( n9379 & n9449 ) ;
  assign n9452 = x113 & n5979 ;
  assign n9453 = ( x115 & n5969 ) | ( x115 & n9452 ) | ( n5969 & n9452 ) ;
  assign n9454 = n9452 | n9453 ;
  assign n9455 = x114 & ~n5970 ;
  assign n9456 = ( x114 & n9454 ) | ( x114 & ~n9455 ) | ( n9454 & ~n9455 ) ;
  assign n9457 = n5968 & n9414 ;
  assign n9458 = n9456 | n9457 ;
  assign n9459 = n9458 ^ x5 ^ 1'b0 ;
  assign n9460 = n9459 ^ n9359 ^ n9132 ;
  assign n9461 = ( n9132 & n9359 ) | ( n9132 & n9459 ) | ( n9359 & n9459 ) ;
  assign n9462 = x113 & n5011 ;
  assign n9463 = ( x115 & n5012 ) | ( x115 & n9462 ) | ( n5012 & n9462 ) ;
  assign n9464 = n9462 | n9463 ;
  assign n9465 = x114 & ~n5008 ;
  assign n9466 = ( x114 & n9464 ) | ( x114 & ~n9465 ) | ( n9464 & ~n9465 ) ;
  assign n9467 = n5020 & n9414 ;
  assign n9468 = n9466 | n9467 ;
  assign n9469 = n9468 ^ x17 ^ 1'b0 ;
  assign n9470 = n9469 ^ n9185 ^ n9019 ;
  assign n9471 = ( n9019 & n9185 ) | ( n9019 & n9469 ) | ( n9185 & n9469 ) ;
  assign n9472 = x113 & n4790 ;
  assign n9473 = ( x115 & n4792 ) | ( x115 & n9472 ) | ( n4792 & n9472 ) ;
  assign n9474 = n9472 | n9473 ;
  assign n9475 = x114 & ~n4786 ;
  assign n9476 = ( x114 & n9474 ) | ( x114 & ~n9475 ) | ( n9474 & ~n9475 ) ;
  assign n9477 = n4787 & n9414 ;
  assign n9478 = n9476 | n9477 ;
  assign n9479 = n9478 ^ x20 ^ 1'b0 ;
  assign n9480 = n9479 ^ n9356 ^ n9145 ;
  assign n9481 = ( n9145 & n9356 ) | ( n9145 & n9479 ) | ( n9356 & n9479 ) ;
  assign n9482 = x113 & n5718 ;
  assign n9483 = ( x115 & n5720 ) | ( x115 & n9482 ) | ( n5720 & n9482 ) ;
  assign n9484 = n9482 | n9483 ;
  assign n9485 = x114 & ~n5727 ;
  assign n9486 = ( x114 & n9484 ) | ( x114 & ~n9485 ) | ( n9484 & ~n9485 ) ;
  assign n9487 = n5726 & n9414 ;
  assign n9488 = n9486 | n9487 ;
  assign n9489 = n9488 ^ x8 ^ 1'b0 ;
  assign n9490 = n9489 ^ n9370 ^ n9194 ;
  assign n9491 = ( n9194 & n9370 ) | ( n9194 & n9489 ) | ( n9370 & n9489 ) ;
  assign n9492 = x113 & n4972 ;
  assign n9493 = x112 & n6104 ;
  assign n9494 = ( x114 & n6105 ) | ( x114 & n9493 ) | ( n6105 & n9493 ) ;
  assign n9495 = n9493 | n9494 ;
  assign n9496 = ( x115 & n4985 ) | ( x115 & n9492 ) | ( n4985 & n9492 ) ;
  assign n9497 = n9492 | n9496 ;
  assign n9498 = x114 & ~n4980 ;
  assign n9499 = ( x114 & n9497 ) | ( x114 & ~n9498 ) | ( n9497 & ~n9498 ) ;
  assign n9500 = n4987 & n9414 ;
  assign n9501 = n9499 | n9500 ;
  assign n9502 = x113 & ~n6107 ;
  assign n9503 = ( x113 & n9495 ) | ( x113 & ~n9502 ) | ( n9495 & ~n9502 ) ;
  assign n9504 = ~n6108 & n9279 ;
  assign n9505 = ( n9279 & n9503 ) | ( n9279 & ~n9504 ) | ( n9503 & ~n9504 ) ;
  assign n9506 = n9501 ^ x14 ^ 1'b0 ;
  assign n9507 = ( n9101 & n9393 ) | ( n9101 & n9506 ) | ( n9393 & n9506 ) ;
  assign n9508 = n9505 ^ x2 ^ 1'b0 ;
  assign n9509 = n9506 ^ n9393 ^ n9101 ;
  assign n9510 = ( n9040 & n9215 ) | ( n9040 & n9508 ) | ( n9215 & n9508 ) ;
  assign n9511 = n9508 ^ n9215 ^ n9040 ;
  assign n9512 = x114 & n4972 ;
  assign n9513 = n9423 ^ x116 ^ x115 ;
  assign n9514 = ( x116 & n4985 ) | ( x116 & n9512 ) | ( n4985 & n9512 ) ;
  assign n9515 = n9512 | n9514 ;
  assign n9516 = x115 & ~n4980 ;
  assign n9517 = ( x115 & n9515 ) | ( x115 & ~n9516 ) | ( n9515 & ~n9516 ) ;
  assign n9518 = n4987 & n9513 ;
  assign n9519 = n9517 | n9518 ;
  assign n9520 = n9519 ^ x14 ^ 1'b0 ;
  assign n9521 = ( n9205 & n9507 ) | ( n9205 & n9520 ) | ( n9507 & n9520 ) ;
  assign n9522 = n9520 ^ n9507 ^ n9205 ;
  assign n9523 = x113 & n6104 ;
  assign n9524 = ( x115 & n6105 ) | ( x115 & n9523 ) | ( n6105 & n9523 ) ;
  assign n9525 = n9523 | n9524 ;
  assign n9526 = x114 & ~n6107 ;
  assign n9527 = ( x114 & n9525 ) | ( x114 & ~n9526 ) | ( n9525 & ~n9526 ) ;
  assign n9528 = ~n6108 & n9414 ;
  assign n9529 = ( n9414 & n9527 ) | ( n9414 & ~n9528 ) | ( n9527 & ~n9528 ) ;
  assign n9530 = n9529 ^ x2 ^ 1'b0 ;
  assign n9531 = n9530 ^ n9510 ^ n9165 ;
  assign n9532 = ( n9165 & n9510 ) | ( n9165 & n9530 ) | ( n9510 & n9530 ) ;
  assign n9533 = x114 & n5979 ;
  assign n9534 = ( x116 & n5969 ) | ( x116 & n9533 ) | ( n5969 & n9533 ) ;
  assign n9535 = n9533 | n9534 ;
  assign n9536 = x115 & ~n5970 ;
  assign n9537 = ( x115 & n9535 ) | ( x115 & ~n9536 ) | ( n9535 & ~n9536 ) ;
  assign n9538 = n5968 & n9513 ;
  assign n9539 = n9537 | n9538 ;
  assign n9540 = n9539 ^ x5 ^ 1'b0 ;
  assign n9541 = ( n9226 & n9461 ) | ( n9226 & n9540 ) | ( n9461 & n9540 ) ;
  assign n9542 = ( x115 & x116 ) | ( x115 & n9423 ) | ( x116 & n9423 ) ;
  assign n9543 = n9540 ^ n9461 ^ n9226 ;
  assign n9544 = x113 & n5499 ;
  assign n9545 = ( x115 & n5497 ) | ( x115 & n9544 ) | ( n5497 & n9544 ) ;
  assign n9546 = n9544 | n9545 ;
  assign n9547 = x114 & ~n5502 ;
  assign n9548 = ( x114 & n9546 ) | ( x114 & ~n9547 ) | ( n9546 & ~n9547 ) ;
  assign n9549 = n5501 & n9414 ;
  assign n9550 = n9548 | n9549 ;
  assign n9551 = n9550 ^ x11 ^ 1'b0 ;
  assign n9552 = n9551 ^ n9289 ^ n9155 ;
  assign n9553 = ( n9155 & n9289 ) | ( n9155 & n9551 ) | ( n9289 & n9551 ) ;
  assign n9554 = x114 & n6104 ;
  assign n9555 = ( x116 & n6105 ) | ( x116 & n9554 ) | ( n6105 & n9554 ) ;
  assign n9556 = n9554 | n9555 ;
  assign n9557 = x115 & ~n6107 ;
  assign n9558 = ( x115 & n9556 ) | ( x115 & ~n9557 ) | ( n9556 & ~n9557 ) ;
  assign n9559 = ~n6108 & n9513 ;
  assign n9560 = ( n9513 & n9558 ) | ( n9513 & ~n9559 ) | ( n9558 & ~n9559 ) ;
  assign n9561 = n9560 ^ x2 ^ 1'b0 ;
  assign n9562 = n9561 ^ n9532 ^ n9236 ;
  assign n9563 = ( n9236 & n9532 ) | ( n9236 & n9561 ) | ( n9532 & n9561 ) ;
  assign n9564 = x116 & ~n6107 ;
  assign n9565 = x115 & n6104 ;
  assign n9566 = ( x117 & n6105 ) | ( x117 & n9565 ) | ( n6105 & n9565 ) ;
  assign n9567 = n9565 | n9566 ;
  assign n9568 = ( x116 & ~n9564 ) | ( x116 & n9567 ) | ( ~n9564 & n9567 ) ;
  assign n9569 = n9542 ^ x117 ^ x116 ;
  assign n9570 = ~n6108 & n9569 ;
  assign n9571 = ( n9568 & n9569 ) | ( n9568 & ~n9570 ) | ( n9569 & ~n9570 ) ;
  assign n9572 = n9571 ^ x2 ^ 1'b0 ;
  assign n9573 = ( n9358 & n9563 ) | ( n9358 & n9572 ) | ( n9563 & n9572 ) ;
  assign n9574 = n9572 ^ n9563 ^ n9358 ;
  assign n9575 = x115 & n5979 ;
  assign n9576 = ( x117 & n5969 ) | ( x117 & n9575 ) | ( n5969 & n9575 ) ;
  assign n9577 = n9575 | n9576 ;
  assign n9578 = x116 & ~n5970 ;
  assign n9579 = ( x116 & n9577 ) | ( x116 & ~n9578 ) | ( n9577 & ~n9578 ) ;
  assign n9580 = n5968 & n9569 ;
  assign n9581 = n9579 | n9580 ;
  assign n9582 = ( x116 & x117 ) | ( x116 & n9542 ) | ( x117 & n9542 ) ;
  assign n9583 = n9581 ^ x5 ^ 1'b0 ;
  assign n9584 = n9583 ^ n9541 ^ n9368 ;
  assign n9585 = ( n9368 & n9541 ) | ( n9368 & n9583 ) | ( n9541 & n9583 ) ;
  assign n9586 = x114 & n5011 ;
  assign n9587 = ( x116 & n5012 ) | ( x116 & n9586 ) | ( n5012 & n9586 ) ;
  assign n9588 = n9586 | n9587 ;
  assign n9589 = x115 & ~n5008 ;
  assign n9590 = ( x115 & n9588 ) | ( x115 & ~n9589 ) | ( n9588 & ~n9589 ) ;
  assign n9591 = n5020 & n9513 ;
  assign n9592 = n9590 | n9591 ;
  assign n9593 = n9592 ^ x17 ^ 1'b0 ;
  assign n9594 = ( n9184 & n9245 ) | ( n9184 & n9593 ) | ( n9245 & n9593 ) ;
  assign n9595 = n9593 ^ n9245 ^ n9184 ;
  assign n9596 = x114 & n5499 ;
  assign n9597 = ( x116 & n5497 ) | ( x116 & n9596 ) | ( n5497 & n9596 ) ;
  assign n9598 = n9596 | n9597 ;
  assign n9599 = x115 & ~n5502 ;
  assign n9600 = ( x115 & n9598 ) | ( x115 & ~n9599 ) | ( n9598 & ~n9599 ) ;
  assign n9601 = n5501 & n9513 ;
  assign n9602 = n9600 | n9601 ;
  assign n9603 = n9602 ^ x11 ^ 1'b0 ;
  assign n9604 = ( n9255 & n9553 ) | ( n9255 & n9603 ) | ( n9553 & n9603 ) ;
  assign n9605 = n9603 ^ n9553 ^ n9255 ;
  assign n9606 = x115 & n5011 ;
  assign n9607 = ( x117 & n5012 ) | ( x117 & n9606 ) | ( n5012 & n9606 ) ;
  assign n9608 = n9606 | n9607 ;
  assign n9609 = x116 & ~n5008 ;
  assign n9610 = ( x116 & n9608 ) | ( x116 & ~n9609 ) | ( n9608 & ~n9609 ) ;
  assign n9611 = ( n5020 & n9569 ) | ( n5020 & n9610 ) | ( n9569 & n9610 ) ;
  assign n9612 = n9610 | n9611 ;
  assign n9613 = n9612 ^ x17 ^ 1'b0 ;
  assign n9614 = ( n9246 & n9357 ) | ( n9246 & n9613 ) | ( n9357 & n9613 ) ;
  assign n9615 = n9613 ^ n9357 ^ n9246 ;
  assign n9616 = x115 & n5499 ;
  assign n9617 = ( x117 & n5497 ) | ( x117 & n9616 ) | ( n5497 & n9616 ) ;
  assign n9618 = n9616 | n9617 ;
  assign n9619 = x116 & ~n5502 ;
  assign n9620 = ( x116 & n9618 ) | ( x116 & ~n9619 ) | ( n9618 & ~n9619 ) ;
  assign n9621 = n5501 & n9569 ;
  assign n9622 = n9620 | n9621 ;
  assign n9623 = n9622 ^ x11 ^ 1'b0 ;
  assign n9624 = n9623 ^ n9604 ^ n9394 ;
  assign n9625 = ( n9394 & n9604 ) | ( n9394 & n9623 ) | ( n9604 & n9623 ) ;
  assign n9626 = x115 & n3734 ;
  assign n9627 = ( x117 & n3732 ) | ( x117 & n9626 ) | ( n3732 & n9626 ) ;
  assign n9628 = n9626 | n9627 ;
  assign n9629 = x116 & ~n3737 ;
  assign n9630 = ( x116 & n9628 ) | ( x116 & ~n9629 ) | ( n9628 & ~n9629 ) ;
  assign n9631 = n3736 & n9569 ;
  assign n9632 = n9630 | n9631 ;
  assign n9633 = n9632 ^ x26 ^ 1'b0 ;
  assign n9634 = n9633 ^ n9339 ^ n9277 ;
  assign n9635 = ( n9277 & n9339 ) | ( n9277 & n9633 ) | ( n9339 & n9633 ) ;
  assign n9636 = x115 & n4972 ;
  assign n9637 = ( x117 & n4985 ) | ( x117 & n9636 ) | ( n4985 & n9636 ) ;
  assign n9638 = n9636 | n9637 ;
  assign n9639 = x116 & ~n4980 ;
  assign n9640 = ( x116 & n9638 ) | ( x116 & ~n9639 ) | ( n9638 & ~n9639 ) ;
  assign n9641 = n4987 & n9569 ;
  assign n9642 = n9640 | n9641 ;
  assign n9643 = n9642 ^ x14 ^ 1'b0 ;
  assign n9644 = ( n9309 & n9521 ) | ( n9309 & n9643 ) | ( n9521 & n9643 ) ;
  assign n9645 = n9643 ^ n9521 ^ n9309 ;
  assign n9646 = x114 & n5718 ;
  assign n9647 = x115 & ~n5727 ;
  assign n9648 = ( x116 & n5720 ) | ( x116 & n9646 ) | ( n5720 & n9646 ) ;
  assign n9649 = n9646 | n9648 ;
  assign n9650 = n5726 & n9513 ;
  assign n9651 = ( x115 & ~n9647 ) | ( x115 & n9649 ) | ( ~n9647 & n9649 ) ;
  assign n9652 = n9650 | n9651 ;
  assign n9653 = n9652 ^ x8 ^ 1'b0 ;
  assign n9654 = ( n9267 & n9491 ) | ( n9267 & n9653 ) | ( n9491 & n9653 ) ;
  assign n9655 = x115 & n5718 ;
  assign n9656 = n9653 ^ n9491 ^ n9267 ;
  assign n9657 = ( x117 & n5720 ) | ( x117 & n9655 ) | ( n5720 & n9655 ) ;
  assign n9658 = x116 & ~n5727 ;
  assign n9659 = n9655 | n9657 ;
  assign n9660 = ( x116 & ~n9658 ) | ( x116 & n9659 ) | ( ~n9658 & n9659 ) ;
  assign n9661 = x116 & n5718 ;
  assign n9662 = n5726 & n9569 ;
  assign n9663 = n9660 | n9662 ;
  assign n9664 = ( x118 & n5720 ) | ( x118 & n9661 ) | ( n5720 & n9661 ) ;
  assign n9665 = n9661 | n9664 ;
  assign n9666 = n9663 ^ x8 ^ 1'b0 ;
  assign n9667 = ( n9288 & n9654 ) | ( n9288 & n9666 ) | ( n9654 & n9666 ) ;
  assign n9668 = n9666 ^ n9654 ^ n9288 ;
  assign n9669 = x117 & ~n5727 ;
  assign n9670 = ( x117 & n9665 ) | ( x117 & ~n9669 ) | ( n9665 & ~n9669 ) ;
  assign n9671 = n9582 ^ x118 ^ x117 ;
  assign n9672 = n5726 & n9671 ;
  assign n9673 = n9670 | n9672 ;
  assign n9674 = n9673 ^ x8 ^ 1'b0 ;
  assign n9675 = ( x117 & x118 ) | ( x117 & n9582 ) | ( x118 & n9582 ) ;
  assign n9676 = ( n9552 & n9667 ) | ( n9552 & n9674 ) | ( n9667 & n9674 ) ;
  assign n9677 = n9674 ^ n9667 ^ n9552 ;
  assign n9678 = x116 & n5979 ;
  assign n9679 = ( x118 & n5969 ) | ( x118 & n9678 ) | ( n5969 & n9678 ) ;
  assign n9680 = n9678 | n9679 ;
  assign n9681 = x117 & ~n5970 ;
  assign n9682 = ( x117 & n9680 ) | ( x117 & ~n9681 ) | ( n9680 & ~n9681 ) ;
  assign n9683 = n5968 & n9671 ;
  assign n9684 = n9682 | n9683 ;
  assign n9685 = n9684 ^ x5 ^ 1'b0 ;
  assign n9686 = ( n9490 & n9585 ) | ( n9490 & n9685 ) | ( n9585 & n9685 ) ;
  assign n9687 = n9685 ^ n9585 ^ n9490 ;
  assign n9688 = x116 & n4972 ;
  assign n9689 = ( x118 & n4985 ) | ( x118 & n9688 ) | ( n4985 & n9688 ) ;
  assign n9690 = n9688 | n9689 ;
  assign n9691 = x117 & ~n4980 ;
  assign n9692 = ( x117 & n9690 ) | ( x117 & ~n9691 ) | ( n9690 & ~n9691 ) ;
  assign n9693 = ( n4987 & n9671 ) | ( n4987 & n9692 ) | ( n9671 & n9692 ) ;
  assign n9694 = n9692 | n9693 ;
  assign n9695 = n9694 ^ x14 ^ 1'b0 ;
  assign n9696 = ( n9308 & n9470 ) | ( n9308 & n9695 ) | ( n9470 & n9695 ) ;
  assign n9697 = n9695 ^ n9470 ^ n9308 ;
  assign n9698 = x116 & n6104 ;
  assign n9699 = ( x118 & n6105 ) | ( x118 & n9698 ) | ( n6105 & n9698 ) ;
  assign n9700 = n9698 | n9699 ;
  assign n9701 = x117 & ~n6107 ;
  assign n9702 = ( x117 & n9700 ) | ( x117 & ~n9701 ) | ( n9700 & ~n9701 ) ;
  assign n9703 = ~n6108 & n9671 ;
  assign n9704 = ( n9671 & n9702 ) | ( n9671 & ~n9703 ) | ( n9702 & ~n9703 ) ;
  assign n9705 = n9704 ^ x2 ^ 1'b0 ;
  assign n9706 = n9705 ^ n9573 ^ n9460 ;
  assign n9707 = ( n9460 & n9573 ) | ( n9460 & n9705 ) | ( n9573 & n9705 ) ;
  assign n9708 = x116 & n5011 ;
  assign n9709 = ( x118 & n5012 ) | ( x118 & n9708 ) | ( n5012 & n9708 ) ;
  assign n9710 = n9708 | n9709 ;
  assign n9711 = x117 & ~n5008 ;
  assign n9712 = ( x117 & n9710 ) | ( x117 & ~n9711 ) | ( n9710 & ~n9711 ) ;
  assign n9713 = n5020 & n9671 ;
  assign n9714 = n9712 | n9713 ;
  assign n9715 = n9714 ^ x17 ^ 1'b0 ;
  assign n9716 = n9715 ^ n9614 ^ n9480 ;
  assign n9717 = ( n9480 & n9614 ) | ( n9480 & n9715 ) | ( n9614 & n9715 ) ;
  assign n9718 = x116 & n5499 ;
  assign n9719 = ( x118 & n5497 ) | ( x118 & n9718 ) | ( n5497 & n9718 ) ;
  assign n9720 = n9718 | n9719 ;
  assign n9721 = x117 & ~n5502 ;
  assign n9722 = ( x117 & n9720 ) | ( x117 & ~n9721 ) | ( n9720 & ~n9721 ) ;
  assign n9723 = n5501 & n9671 ;
  assign n9724 = n9722 | n9723 ;
  assign n9725 = n9724 ^ x11 ^ 1'b0 ;
  assign n9726 = ( n9509 & n9625 ) | ( n9509 & n9725 ) | ( n9625 & n9725 ) ;
  assign n9727 = n9725 ^ n9625 ^ n9509 ;
  assign n9728 = x117 & n5718 ;
  assign n9729 = ( x119 & n5720 ) | ( x119 & n9728 ) | ( n5720 & n9728 ) ;
  assign n9730 = n9728 | n9729 ;
  assign n9731 = x118 & ~n5727 ;
  assign n9732 = ( x118 & n9730 ) | ( x118 & ~n9731 ) | ( n9730 & ~n9731 ) ;
  assign n9733 = n9675 ^ x119 ^ x118 ;
  assign n9734 = n5726 & n9733 ;
  assign n9735 = n9732 | n9734 ;
  assign n9736 = x118 & ~n6107 ;
  assign n9737 = x117 & n6104 ;
  assign n9738 = x118 & n6104 ;
  assign n9739 = ( x119 & n6105 ) | ( x119 & n9737 ) | ( n6105 & n9737 ) ;
  assign n9740 = n9737 | n9739 ;
  assign n9741 = ( x118 & ~n9736 ) | ( x118 & n9740 ) | ( ~n9736 & n9740 ) ;
  assign n9742 = ( x120 & n6105 ) | ( x120 & n9738 ) | ( n6105 & n9738 ) ;
  assign n9743 = x117 & n4972 ;
  assign n9744 = n9738 | n9742 ;
  assign n9745 = ~n6108 & n9733 ;
  assign n9746 = ( n9733 & n9741 ) | ( n9733 & ~n9745 ) | ( n9741 & ~n9745 ) ;
  assign n9747 = x119 & ~n6107 ;
  assign n9748 = n9746 ^ x2 ^ 1'b0 ;
  assign n9749 = ( x119 & n9744 ) | ( x119 & ~n9747 ) | ( n9744 & ~n9747 ) ;
  assign n9750 = ( x118 & x119 ) | ( x118 & n9675 ) | ( x119 & n9675 ) ;
  assign n9751 = ( x119 & n4985 ) | ( x119 & n9743 ) | ( n4985 & n9743 ) ;
  assign n9752 = n9743 | n9751 ;
  assign n9753 = n9735 ^ x8 ^ 1'b0 ;
  assign n9754 = ( n9543 & n9707 ) | ( n9543 & n9748 ) | ( n9707 & n9748 ) ;
  assign n9755 = n9748 ^ n9707 ^ n9543 ;
  assign n9756 = n9750 ^ x120 ^ x119 ;
  assign n9757 = ~n6108 & n9756 ;
  assign n9758 = ( n9749 & n9756 ) | ( n9749 & ~n9757 ) | ( n9756 & ~n9757 ) ;
  assign n9759 = n9758 ^ x2 ^ 1'b0 ;
  assign n9760 = ( n9584 & n9754 ) | ( n9584 & n9759 ) | ( n9754 & n9759 ) ;
  assign n9761 = n9759 ^ n9754 ^ n9584 ;
  assign n9762 = n4987 & n9733 ;
  assign n9763 = x118 & ~n4980 ;
  assign n9764 = ( x118 & n9752 ) | ( x118 & ~n9763 ) | ( n9752 & ~n9763 ) ;
  assign n9765 = n9753 ^ n9676 ^ n9605 ;
  assign n9766 = n9762 | n9764 ;
  assign n9767 = ( n9605 & n9676 ) | ( n9605 & n9753 ) | ( n9676 & n9753 ) ;
  assign n9768 = x118 & ~n5502 ;
  assign n9769 = n9766 ^ x14 ^ 1'b0 ;
  assign n9770 = x117 & n5499 ;
  assign n9771 = ( x119 & n5497 ) | ( x119 & n9770 ) | ( n5497 & n9770 ) ;
  assign n9772 = n9770 | n9771 ;
  assign n9773 = ( n9471 & n9595 ) | ( n9471 & n9769 ) | ( n9595 & n9769 ) ;
  assign n9774 = ( x118 & ~n9768 ) | ( x118 & n9772 ) | ( ~n9768 & n9772 ) ;
  assign n9775 = n9769 ^ n9595 ^ n9471 ;
  assign n9776 = x117 & n5979 ;
  assign n9777 = x119 & ~n4980 ;
  assign n9778 = n5501 & n9733 ;
  assign n9779 = n9774 | n9778 ;
  assign n9780 = n9779 ^ x11 ^ 1'b0 ;
  assign n9781 = n9780 ^ n9726 ^ n9522 ;
  assign n9782 = ( n9522 & n9726 ) | ( n9522 & n9780 ) | ( n9726 & n9780 ) ;
  assign n9783 = ( x119 & x120 ) | ( x119 & n9750 ) | ( x120 & n9750 ) ;
  assign n9784 = x118 & n4972 ;
  assign n9785 = ( x120 & n4985 ) | ( x120 & n9784 ) | ( n4985 & n9784 ) ;
  assign n9786 = n9784 | n9785 ;
  assign n9787 = ( x119 & ~n9777 ) | ( x119 & n9786 ) | ( ~n9777 & n9786 ) ;
  assign n9788 = n5968 & n9733 ;
  assign n9789 = ( x119 & n5969 ) | ( x119 & n9776 ) | ( n5969 & n9776 ) ;
  assign n9790 = n9776 | n9789 ;
  assign n9791 = x118 & ~n5970 ;
  assign n9792 = ( x118 & n9790 ) | ( x118 & ~n9791 ) | ( n9790 & ~n9791 ) ;
  assign n9793 = n4987 & n9756 ;
  assign n9794 = n9788 | n9792 ;
  assign n9795 = n9794 ^ x5 ^ 1'b0 ;
  assign n9796 = n9787 | n9793 ;
  assign n9797 = n9796 ^ x14 ^ 1'b0 ;
  assign n9798 = ( n9656 & n9686 ) | ( n9656 & n9795 ) | ( n9686 & n9795 ) ;
  assign n9799 = n9795 ^ n9686 ^ n9656 ;
  assign n9800 = n9797 ^ n9615 ^ n9594 ;
  assign n9801 = ( n9594 & n9615 ) | ( n9594 & n9797 ) | ( n9615 & n9797 ) ;
  assign n9802 = ( x120 & x121 ) | ( x120 & n9783 ) | ( x121 & n9783 ) ;
  assign n9803 = x120 & n6104 ;
  assign n9804 = x121 & ~n6107 ;
  assign n9805 = ( x122 & n6105 ) | ( x122 & n9803 ) | ( n6105 & n9803 ) ;
  assign n9806 = n9802 ^ x122 ^ x121 ;
  assign n9807 = n9803 | n9805 ;
  assign n9808 = n9783 ^ x121 ^ x120 ;
  assign n9809 = ( x121 & ~n9804 ) | ( x121 & n9807 ) | ( ~n9804 & n9807 ) ;
  assign n9810 = ~n6108 & n9806 ;
  assign n9811 = ( x121 & x122 ) | ( x121 & n9802 ) | ( x122 & n9802 ) ;
  assign n9812 = ( n9806 & n9809 ) | ( n9806 & ~n9810 ) | ( n9809 & ~n9810 ) ;
  assign n9813 = x119 & n6104 ;
  assign n9814 = n9812 ^ x2 ^ 1'b0 ;
  assign n9815 = ( x121 & n6105 ) | ( x121 & n9813 ) | ( n6105 & n9813 ) ;
  assign n9816 = x120 & ~n6107 ;
  assign n9817 = n9813 | n9815 ;
  assign n9818 = ( x120 & ~n9816 ) | ( x120 & n9817 ) | ( ~n9816 & n9817 ) ;
  assign n9819 = ~n6108 & n9808 ;
  assign n9820 = ( n9808 & n9818 ) | ( n9808 & ~n9819 ) | ( n9818 & ~n9819 ) ;
  assign n9821 = n9820 ^ x2 ^ 1'b0 ;
  assign n9822 = n9821 ^ n9760 ^ n9687 ;
  assign n9823 = ( n9687 & n9760 ) | ( n9687 & n9821 ) | ( n9760 & n9821 ) ;
  assign n9824 = ( n9799 & n9814 ) | ( n9799 & n9823 ) | ( n9814 & n9823 ) ;
  assign n9825 = x121 & n6104 ;
  assign n9826 = n9823 ^ n9814 ^ n9799 ;
  assign n9827 = ( x123 & n6105 ) | ( x123 & n9825 ) | ( n6105 & n9825 ) ;
  assign n9828 = n9811 ^ x123 ^ x122 ;
  assign n9829 = n9825 | n9827 ;
  assign n9830 = x122 & ~n6107 ;
  assign n9831 = ( x122 & n9829 ) | ( x122 & ~n9830 ) | ( n9829 & ~n9830 ) ;
  assign n9832 = ~n6108 & n9828 ;
  assign n9833 = ( n9828 & n9831 ) | ( n9828 & ~n9832 ) | ( n9831 & ~n9832 ) ;
  assign n9834 = n9833 ^ x2 ^ 1'b0 ;
  assign n9835 = ( x122 & x123 ) | ( x122 & n9811 ) | ( x123 & n9811 ) ;
  assign n9836 = x118 & n5979 ;
  assign n9837 = ( x120 & n5969 ) | ( x120 & n9836 ) | ( n5969 & n9836 ) ;
  assign n9838 = n9836 | n9837 ;
  assign n9839 = x119 & ~n5970 ;
  assign n9840 = ( x119 & n9838 ) | ( x119 & ~n9839 ) | ( n9838 & ~n9839 ) ;
  assign n9841 = n5968 & n9756 ;
  assign n9842 = n9840 | n9841 ;
  assign n9843 = n9842 ^ x5 ^ 1'b0 ;
  assign n9844 = ( n9668 & n9834 ) | ( n9668 & n9843 ) | ( n9834 & n9843 ) ;
  assign n9845 = n9843 ^ n9834 ^ n9668 ;
  assign n9846 = n9845 ^ n9824 ^ n9798 ;
  assign n9847 = ( n9798 & n9824 ) | ( n9798 & n9845 ) | ( n9824 & n9845 ) ;
  assign n9848 = x119 & n5979 ;
  assign n9849 = x120 & ~n5970 ;
  assign n9850 = ( x121 & n5969 ) | ( x121 & n9848 ) | ( n5969 & n9848 ) ;
  assign n9851 = n9848 | n9850 ;
  assign n9852 = x120 & n5979 ;
  assign n9853 = n5968 & n9808 ;
  assign n9854 = ( x122 & n5969 ) | ( x122 & n9852 ) | ( n5969 & n9852 ) ;
  assign n9855 = n9852 | n9854 ;
  assign n9856 = x121 & ~n5970 ;
  assign n9857 = ( x121 & n9855 ) | ( x121 & ~n9856 ) | ( n9855 & ~n9856 ) ;
  assign n9858 = n9835 ^ x124 ^ x123 ;
  assign n9859 = ( x120 & ~n9849 ) | ( x120 & n9851 ) | ( ~n9849 & n9851 ) ;
  assign n9860 = x122 & n6104 ;
  assign n9861 = n9853 | n9859 ;
  assign n9862 = ( x124 & n6105 ) | ( x124 & n9860 ) | ( n6105 & n9860 ) ;
  assign n9863 = n9860 | n9862 ;
  assign n9864 = x123 & ~n6107 ;
  assign n9865 = ( x123 & n9863 ) | ( x123 & ~n9864 ) | ( n9863 & ~n9864 ) ;
  assign n9866 = ~n6108 & n9858 ;
  assign n9867 = ( n9858 & n9865 ) | ( n9858 & ~n9866 ) | ( n9865 & ~n9866 ) ;
  assign n9868 = n9861 ^ x5 ^ 1'b0 ;
  assign n9869 = n9867 ^ x2 ^ 1'b0 ;
  assign n9870 = ( n9677 & n9868 ) | ( n9677 & n9869 ) | ( n9868 & n9869 ) ;
  assign n9871 = n9869 ^ n9868 ^ n9677 ;
  assign n9872 = n5968 & n9806 ;
  assign n9873 = x123 & n6104 ;
  assign n9874 = n9857 | n9872 ;
  assign n9875 = ( x125 & n6105 ) | ( x125 & n9873 ) | ( n6105 & n9873 ) ;
  assign n9876 = n9873 | n9875 ;
  assign n9877 = x124 & ~n6107 ;
  assign n9878 = ( x124 & n9876 ) | ( x124 & ~n9877 ) | ( n9876 & ~n9877 ) ;
  assign n9879 = n9874 ^ x5 ^ 1'b0 ;
  assign n9880 = ( x123 & x124 ) | ( x123 & n9835 ) | ( x124 & n9835 ) ;
  assign n9881 = n9871 ^ n9847 ^ n9844 ;
  assign n9882 = ( n9844 & n9847 ) | ( n9844 & n9871 ) | ( n9847 & n9871 ) ;
  assign n9883 = n9880 ^ x125 ^ x124 ;
  assign n9884 = ~n6108 & n9883 ;
  assign n9885 = ( x124 & x125 ) | ( x124 & n9880 ) | ( x125 & n9880 ) ;
  assign n9886 = ( n9878 & n9883 ) | ( n9878 & ~n9884 ) | ( n9883 & ~n9884 ) ;
  assign n9887 = n9886 ^ x2 ^ 1'b0 ;
  assign n9888 = n9887 ^ n9879 ^ n9765 ;
  assign n9889 = ( n9765 & n9879 ) | ( n9765 & n9887 ) | ( n9879 & n9887 ) ;
  assign n9890 = n9888 ^ n9882 ^ n9870 ;
  assign n9891 = ( n9870 & n9882 ) | ( n9870 & n9888 ) | ( n9882 & n9888 ) ;
  assign n9892 = x121 & n5979 ;
  assign n9893 = ( x123 & n5969 ) | ( x123 & n9892 ) | ( n5969 & n9892 ) ;
  assign n9894 = n9892 | n9893 ;
  assign n9895 = x122 & ~n5970 ;
  assign n9896 = ( x122 & n9894 ) | ( x122 & ~n9895 ) | ( n9894 & ~n9895 ) ;
  assign n9897 = n5968 & n9828 ;
  assign n9898 = n9896 | n9897 ;
  assign n9899 = x118 & n5718 ;
  assign n9900 = ( x120 & n5720 ) | ( x120 & n9899 ) | ( n5720 & n9899 ) ;
  assign n9901 = n9899 | n9900 ;
  assign n9902 = x119 & ~n5727 ;
  assign n9903 = ( x119 & n9901 ) | ( x119 & ~n9902 ) | ( n9901 & ~n9902 ) ;
  assign n9904 = n5726 & n9756 ;
  assign n9905 = n9903 | n9904 ;
  assign n9906 = n9905 ^ x8 ^ 1'b0 ;
  assign n9907 = n9898 ^ x5 ^ 1'b0 ;
  assign n9908 = n9907 ^ n9906 ^ n9624 ;
  assign n9909 = x125 & n6104 ;
  assign n9910 = ( n9624 & n9906 ) | ( n9624 & n9907 ) | ( n9906 & n9907 ) ;
  assign n9911 = ( x127 & n6105 ) | ( x127 & n9909 ) | ( n6105 & n9909 ) ;
  assign n9912 = n9909 | n9911 ;
  assign n9913 = x126 & ~n6107 ;
  assign n9914 = ( x126 & n9912 ) | ( x126 & ~n9913 ) | ( n9912 & ~n9913 ) ;
  assign n9915 = ( x125 & x126 ) | ( x125 & n9885 ) | ( x126 & n9885 ) ;
  assign n9916 = x124 & n6104 ;
  assign n9917 = n9885 ^ x126 ^ x125 ;
  assign n9918 = ( x126 & n6105 ) | ( x126 & n9916 ) | ( n6105 & n9916 ) ;
  assign n9919 = n9916 | n9918 ;
  assign n9920 = x125 & ~n6107 ;
  assign n9921 = ( x125 & n9919 ) | ( x125 & ~n9920 ) | ( n9919 & ~n9920 ) ;
  assign n9922 = ~n6108 & n9917 ;
  assign n9923 = ( n9917 & n9921 ) | ( n9917 & ~n9922 ) | ( n9921 & ~n9922 ) ;
  assign n9924 = n9923 ^ x2 ^ 1'b0 ;
  assign n9925 = ( n9767 & n9908 ) | ( n9767 & n9924 ) | ( n9908 & n9924 ) ;
  assign n9926 = x127 & ~n6107 ;
  assign n9927 = n9924 ^ n9908 ^ n9767 ;
  assign n9928 = ( n9889 & n9891 ) | ( n9889 & n9927 ) | ( n9891 & n9927 ) ;
  assign n9929 = n9927 ^ n9891 ^ n9889 ;
  assign n9930 = x119 & n5718 ;
  assign n9931 = ( x121 & n5720 ) | ( x121 & n9930 ) | ( n5720 & n9930 ) ;
  assign n9932 = n9930 | n9931 ;
  assign n9933 = n5726 & n9808 ;
  assign n9934 = x120 & ~n5727 ;
  assign n9935 = ( x120 & n9932 ) | ( x120 & ~n9934 ) | ( n9932 & ~n9934 ) ;
  assign n9936 = n9933 | n9935 ;
  assign n9937 = n9936 ^ x8 ^ 1'b0 ;
  assign n9938 = x122 & n5979 ;
  assign n9939 = ( x124 & n5969 ) | ( x124 & n9938 ) | ( n5969 & n9938 ) ;
  assign n9940 = x123 & ~n5970 ;
  assign n9941 = n9938 | n9939 ;
  assign n9942 = ( x123 & ~n9940 ) | ( x123 & n9941 ) | ( ~n9940 & n9941 ) ;
  assign n9943 = n5968 & n9858 ;
  assign n9944 = x127 ^ x126 ^ 1'b0 ;
  assign n9945 = n9942 | n9943 ;
  assign n9946 = n9945 ^ x5 ^ 1'b0 ;
  assign n9947 = n9946 ^ n9937 ^ n9727 ;
  assign n9948 = ( n9727 & n9937 ) | ( n9727 & n9946 ) | ( n9937 & n9946 ) ;
  assign n9949 = n9944 ^ n9915 ^ 1'b0 ;
  assign n9950 = ~n6108 & n9949 ;
  assign n9951 = ( n9914 & n9949 ) | ( n9914 & ~n9950 ) | ( n9949 & ~n9950 ) ;
  assign n9952 = n9951 ^ x2 ^ 1'b0 ;
  assign n9953 = n9952 ^ n9947 ^ n9910 ;
  assign n9954 = ( n9910 & n9947 ) | ( n9910 & n9952 ) | ( n9947 & n9952 ) ;
  assign n9955 = x120 & n5718 ;
  assign n9956 = ( x122 & n5720 ) | ( x122 & n9955 ) | ( n5720 & n9955 ) ;
  assign n9957 = ( x126 & x127 ) | ( x126 & n9915 ) | ( x127 & n9915 ) ;
  assign n9958 = n9957 ^ n9944 ^ x126 ;
  assign n9959 = n9955 | n9956 ;
  assign n9960 = x121 & ~n5727 ;
  assign n9961 = ( x121 & n9959 ) | ( x121 & ~n9960 ) | ( n9959 & ~n9960 ) ;
  assign n9962 = ( n9925 & n9928 ) | ( n9925 & n9953 ) | ( n9928 & n9953 ) ;
  assign n9963 = n9953 ^ n9928 ^ n9925 ;
  assign n9964 = n5726 & n9806 ;
  assign n9965 = n9961 | n9964 ;
  assign n9966 = x126 & n6104 ;
  assign n9967 = ( x127 & ~n9926 ) | ( x127 & n9966 ) | ( ~n9926 & n9966 ) ;
  assign n9968 = x127 & n9957 ;
  assign n9969 = n6108 & n9968 ;
  assign n9970 = ( n6108 & n9958 ) | ( n6108 & n9966 ) | ( n9958 & n9966 ) ;
  assign n9971 = n9965 ^ x8 ^ 1'b0 ;
  assign n9972 = x127 & n6104 ;
  assign n9973 = n9969 ^ x2 ^ 1'b0 ;
  assign n9974 = ( x2 & n9969 ) | ( x2 & n9972 ) | ( n9969 & n9972 ) ;
  assign n9975 = n9967 | n9970 ;
  assign n9976 = x124 & ~n5970 ;
  assign n9977 = n9975 ^ x2 ^ 1'b0 ;
  assign n9978 = ( n9969 & n9973 ) | ( n9969 & ~n9974 ) | ( n9973 & ~n9974 ) ;
  assign n9979 = x123 & n5979 ;
  assign n9980 = ( x125 & n5969 ) | ( x125 & n9979 ) | ( n5969 & n9979 ) ;
  assign n9981 = n9979 | n9980 ;
  assign n9982 = ( x124 & ~n9976 ) | ( x124 & n9981 ) | ( ~n9976 & n9981 ) ;
  assign n9983 = n5968 & n9883 ;
  assign n9984 = n9982 | n9983 ;
  assign n9985 = n9984 ^ x5 ^ 1'b0 ;
  assign n9986 = n9985 ^ n9971 ^ n9781 ;
  assign n9987 = n9986 ^ n9977 ^ n9948 ;
  assign n9988 = ( n9781 & n9971 ) | ( n9781 & n9985 ) | ( n9971 & n9985 ) ;
  assign n9989 = n9987 ^ n9962 ^ n9954 ;
  assign n9990 = ( n9948 & n9977 ) | ( n9948 & n9986 ) | ( n9977 & n9986 ) ;
  assign n9991 = ( n9954 & n9962 ) | ( n9954 & n9987 ) | ( n9962 & n9987 ) ;
  assign n9992 = x118 & n5499 ;
  assign n9993 = ( x120 & n5497 ) | ( x120 & n9992 ) | ( n5497 & n9992 ) ;
  assign n9994 = n9992 | n9993 ;
  assign n9995 = x121 & n5718 ;
  assign n9996 = x119 & ~n5502 ;
  assign n9997 = ( x119 & n9994 ) | ( x119 & ~n9996 ) | ( n9994 & ~n9996 ) ;
  assign n9998 = ( x123 & n5720 ) | ( x123 & n9995 ) | ( n5720 & n9995 ) ;
  assign n9999 = n9995 | n9998 ;
  assign n10000 = n5501 & n9756 ;
  assign n10001 = n9997 | n10000 ;
  assign n10002 = x122 & ~n5727 ;
  assign n10003 = n10001 ^ x11 ^ 1'b0 ;
  assign n10004 = ( x122 & n9999 ) | ( x122 & ~n10002 ) | ( n9999 & ~n10002 ) ;
  assign n10005 = n5726 & n9828 ;
  assign n10006 = n10004 | n10005 ;
  assign n10007 = n10006 ^ x8 ^ 1'b0 ;
  assign n10008 = n10007 ^ n10003 ^ n9645 ;
  assign n10009 = ( n9645 & n10003 ) | ( n9645 & n10007 ) | ( n10003 & n10007 ) ;
  assign n10010 = x124 & n5979 ;
  assign n10011 = ( x126 & n5969 ) | ( x126 & n10010 ) | ( n5969 & n10010 ) ;
  assign n10012 = n10010 | n10011 ;
  assign n10013 = x125 & n5979 ;
  assign n10014 = ( x127 & n5969 ) | ( x127 & n10013 ) | ( n5969 & n10013 ) ;
  assign n10015 = n10013 | n10014 ;
  assign n10016 = x125 & ~n5970 ;
  assign n10017 = ( x125 & n10012 ) | ( x125 & ~n10016 ) | ( n10012 & ~n10016 ) ;
  assign n10018 = n5968 & n9917 ;
  assign n10019 = n10017 | n10018 ;
  assign n10020 = x126 & ~n5970 ;
  assign n10021 = n10019 ^ x5 ^ 1'b0 ;
  assign n10022 = x127 & ~n5970 ;
  assign n10023 = ( x126 & n10015 ) | ( x126 & ~n10020 ) | ( n10015 & ~n10020 ) ;
  assign n10024 = n5968 & n9949 ;
  assign n10025 = n10023 | n10024 ;
  assign n10026 = x127 & n5979 ;
  assign n10027 = x126 & n5979 ;
  assign n10028 = ( x127 & ~n10022 ) | ( x127 & n10027 ) | ( ~n10022 & n10027 ) ;
  assign n10029 = ( n5968 & n9958 ) | ( n5968 & n10027 ) | ( n9958 & n10027 ) ;
  assign n10030 = n10028 | n10029 ;
  assign n10031 = n10021 ^ n10008 ^ n9782 ;
  assign n10032 = ( n9782 & n10008 ) | ( n9782 & n10021 ) | ( n10008 & n10021 ) ;
  assign n10033 = ( n9978 & n9988 ) | ( n9978 & n10031 ) | ( n9988 & n10031 ) ;
  assign n10034 = n10031 ^ n9988 ^ n9978 ;
  assign n10035 = ( n9990 & n9991 ) | ( n9990 & n10034 ) | ( n9991 & n10034 ) ;
  assign n10036 = n10034 ^ n9991 ^ n9990 ;
  assign n10037 = x120 & n5499 ;
  assign n10038 = ( n5968 & n9968 ) | ( n5968 & n10026 ) | ( n9968 & n10026 ) ;
  assign n10039 = n10026 | n10038 ;
  assign n10040 = ( x122 & n5497 ) | ( x122 & n10037 ) | ( n5497 & n10037 ) ;
  assign n10041 = n10037 | n10040 ;
  assign n10042 = x121 & ~n5502 ;
  assign n10043 = ( x121 & n10041 ) | ( x121 & ~n10042 ) | ( n10041 & ~n10042 ) ;
  assign n10044 = ( n5501 & n9806 ) | ( n5501 & n10043 ) | ( n9806 & n10043 ) ;
  assign n10045 = n10043 | n10044 ;
  assign n10046 = n10045 ^ x11 ^ 1'b0 ;
  assign n10047 = n10046 ^ n9775 ^ n9696 ;
  assign n10048 = n10025 ^ x5 ^ 1'b0 ;
  assign n10049 = ( n9696 & n9775 ) | ( n9696 & n10046 ) | ( n9775 & n10046 ) ;
  assign n10050 = x119 & n5499 ;
  assign n10051 = ( x121 & n5497 ) | ( x121 & n10050 ) | ( n5497 & n10050 ) ;
  assign n10052 = n10050 | n10051 ;
  assign n10053 = x120 & ~n5502 ;
  assign n10054 = ( x120 & n10052 ) | ( x120 & ~n10053 ) | ( n10052 & ~n10053 ) ;
  assign n10055 = n5501 & n9808 ;
  assign n10056 = n10054 | n10055 ;
  assign n10057 = n10056 ^ x11 ^ 1'b0 ;
  assign n10058 = ( n9644 & n9697 ) | ( n9644 & n10057 ) | ( n9697 & n10057 ) ;
  assign n10059 = n10057 ^ n9697 ^ n9644 ;
  assign n10060 = x122 & n5718 ;
  assign n10061 = ( x124 & n5720 ) | ( x124 & n10060 ) | ( n5720 & n10060 ) ;
  assign n10062 = n10060 | n10061 ;
  assign n10063 = x123 & ~n5727 ;
  assign n10064 = ( x123 & n10062 ) | ( x123 & ~n10063 ) | ( n10062 & ~n10063 ) ;
  assign n10065 = n5726 & n9858 ;
  assign n10066 = n10064 | n10065 ;
  assign n10067 = n10066 ^ x8 ^ 1'b0 ;
  assign n10068 = n10067 ^ n10059 ^ n10009 ;
  assign n10069 = ( n10009 & n10059 ) | ( n10009 & n10067 ) | ( n10059 & n10067 ) ;
  assign n10070 = ( n10032 & n10048 ) | ( n10032 & n10068 ) | ( n10048 & n10068 ) ;
  assign n10071 = n10068 ^ n10048 ^ n10032 ;
  assign n10072 = ( n10033 & n10035 ) | ( n10033 & n10071 ) | ( n10035 & n10071 ) ;
  assign n10073 = n10071 ^ n10035 ^ n10033 ;
  assign n10074 = x121 & n5499 ;
  assign n10075 = ( x123 & n5497 ) | ( x123 & n10074 ) | ( n5497 & n10074 ) ;
  assign n10076 = n10074 | n10075 ;
  assign n10077 = x122 & ~n5502 ;
  assign n10078 = ( x122 & n10076 ) | ( x122 & ~n10077 ) | ( n10076 & ~n10077 ) ;
  assign n10079 = n5501 & n9828 ;
  assign n10080 = n10078 | n10079 ;
  assign n10081 = n10080 ^ x11 ^ 1'b0 ;
  assign n10082 = n10030 ^ x5 ^ 1'b0 ;
  assign n10083 = ( n9773 & n9800 ) | ( n9773 & n10081 ) | ( n9800 & n10081 ) ;
  assign n10084 = n10081 ^ n9800 ^ n9773 ;
  assign n10085 = x123 & n5718 ;
  assign n10086 = ( x125 & n5720 ) | ( x125 & n10085 ) | ( n5720 & n10085 ) ;
  assign n10087 = n10085 | n10086 ;
  assign n10088 = x124 & ~n5727 ;
  assign n10089 = ( x124 & n10087 ) | ( x124 & ~n10088 ) | ( n10087 & ~n10088 ) ;
  assign n10090 = ( n5726 & n9883 ) | ( n5726 & n10089 ) | ( n9883 & n10089 ) ;
  assign n10091 = n10089 | n10090 ;
  assign n10092 = n10091 ^ x8 ^ 1'b0 ;
  assign n10093 = ( n10047 & n10058 ) | ( n10047 & n10092 ) | ( n10058 & n10092 ) ;
  assign n10094 = n10092 ^ n10058 ^ n10047 ;
  assign n10095 = n10094 ^ n10082 ^ n10069 ;
  assign n10096 = n10095 ^ n10072 ^ n10070 ;
  assign n10097 = ( n10070 & n10072 ) | ( n10070 & n10095 ) | ( n10072 & n10095 ) ;
  assign n10098 = x119 & n4972 ;
  assign n10099 = ( x121 & n4985 ) | ( x121 & n10098 ) | ( n4985 & n10098 ) ;
  assign n10100 = n10098 | n10099 ;
  assign n10101 = ( n10069 & n10082 ) | ( n10069 & n10094 ) | ( n10082 & n10094 ) ;
  assign n10102 = x120 & ~n4980 ;
  assign n10103 = ( x120 & n10100 ) | ( x120 & ~n10102 ) | ( n10100 & ~n10102 ) ;
  assign n10104 = n4987 & n9808 ;
  assign n10105 = x124 & n5718 ;
  assign n10106 = ( x126 & n5720 ) | ( x126 & n10105 ) | ( n5720 & n10105 ) ;
  assign n10107 = n10105 | n10106 ;
  assign n10108 = n10103 | n10104 ;
  assign n10109 = x126 & ~n5727 ;
  assign n10110 = n10108 ^ x14 ^ 1'b0 ;
  assign n10111 = n10110 ^ n9801 ^ n9716 ;
  assign n10112 = ( n9716 & n9801 ) | ( n9716 & n10110 ) | ( n9801 & n10110 ) ;
  assign n10113 = n5726 & n9949 ;
  assign n10114 = x125 & n5718 ;
  assign n10115 = ( x127 & n5720 ) | ( x127 & n10114 ) | ( n5720 & n10114 ) ;
  assign n10116 = n10114 | n10115 ;
  assign n10117 = x127 & ~n5727 ;
  assign n10118 = ( x126 & ~n10109 ) | ( x126 & n10116 ) | ( ~n10109 & n10116 ) ;
  assign n10119 = n10113 | n10118 ;
  assign n10120 = x126 & n5718 ;
  assign n10121 = ( x127 & ~n10117 ) | ( x127 & n10120 ) | ( ~n10117 & n10120 ) ;
  assign n10122 = x125 & ~n5727 ;
  assign n10123 = x127 & n5718 ;
  assign n10124 = ( n5726 & n9968 ) | ( n5726 & n10123 ) | ( n9968 & n10123 ) ;
  assign n10125 = n10039 ^ x5 ^ 1'b0 ;
  assign n10126 = n10123 | n10124 ;
  assign n10127 = ( x125 & n10107 ) | ( x125 & ~n10122 ) | ( n10107 & ~n10122 ) ;
  assign n10128 = n5501 & n9858 ;
  assign n10129 = ( n5726 & n9917 ) | ( n5726 & n10127 ) | ( n9917 & n10127 ) ;
  assign n10130 = ( n5726 & n9958 ) | ( n5726 & n10120 ) | ( n9958 & n10120 ) ;
  assign n10131 = x123 & ~n5502 ;
  assign n10132 = n10127 | n10129 ;
  assign n10133 = n10121 | n10130 ;
  assign n10134 = n10132 ^ x8 ^ 1'b0 ;
  assign n10135 = x122 & n5499 ;
  assign n10136 = ( x124 & n5497 ) | ( x124 & n10135 ) | ( n5497 & n10135 ) ;
  assign n10137 = n10135 | n10136 ;
  assign n10138 = ( x123 & ~n10131 ) | ( x123 & n10137 ) | ( ~n10131 & n10137 ) ;
  assign n10139 = ( n10049 & n10084 ) | ( n10049 & n10134 ) | ( n10084 & n10134 ) ;
  assign n10140 = n10128 | n10138 ;
  assign n10141 = n10140 ^ x11 ^ 1'b0 ;
  assign n10142 = n10119 ^ x8 ^ 1'b0 ;
  assign n10143 = n10141 ^ n10111 ^ n10083 ;
  assign n10144 = n10143 ^ n10142 ^ n10139 ;
  assign n10145 = n10134 ^ n10084 ^ n10049 ;
  assign n10146 = ( n10083 & n10111 ) | ( n10083 & n10141 ) | ( n10111 & n10141 ) ;
  assign n10147 = n10145 ^ n10125 ^ n10093 ;
  assign n10148 = n10147 ^ n10101 ^ n10097 ;
  assign n10149 = ( n10097 & n10101 ) | ( n10097 & n10147 ) | ( n10101 & n10147 ) ;
  assign n10150 = ( n10093 & n10125 ) | ( n10093 & n10145 ) | ( n10125 & n10145 ) ;
  assign n10151 = ( n10139 & n10142 ) | ( n10139 & n10143 ) | ( n10142 & n10143 ) ;
  assign n10152 = n10150 ^ n10149 ^ n10144 ;
  assign n10153 = ( n10144 & n10149 ) | ( n10144 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10154 = x114 & n4790 ;
  assign n10155 = ( x116 & n4792 ) | ( x116 & n10154 ) | ( n4792 & n10154 ) ;
  assign n10156 = n10154 | n10155 ;
  assign n10157 = x115 & ~n4786 ;
  assign n10158 = ( x115 & n10156 ) | ( x115 & ~n10157 ) | ( n10156 & ~n10157 ) ;
  assign n10159 = n4787 & n9513 ;
  assign n10160 = n10158 | n10159 ;
  assign n10161 = n10160 ^ x20 ^ 1'b0 ;
  assign n10162 = n10161 ^ n9299 ^ n9144 ;
  assign n10163 = ( n9144 & n9299 ) | ( n9144 & n10161 ) | ( n9299 & n10161 ) ;
  assign n10164 = x117 & n5011 ;
  assign n10165 = ( x119 & n5012 ) | ( x119 & n10164 ) | ( n5012 & n10164 ) ;
  assign n10166 = n10164 | n10165 ;
  assign n10167 = x118 & ~n5008 ;
  assign n10168 = ( x118 & n10166 ) | ( x118 & ~n10167 ) | ( n10166 & ~n10167 ) ;
  assign n10169 = n5020 & n9733 ;
  assign n10170 = n10133 ^ x8 ^ 1'b0 ;
  assign n10171 = n10168 | n10169 ;
  assign n10172 = n10171 ^ x17 ^ 1'b0 ;
  assign n10173 = n10172 ^ n10162 ^ n9481 ;
  assign n10174 = ( n9481 & n10162 ) | ( n9481 & n10172 ) | ( n10162 & n10172 ) ;
  assign n10175 = x120 & n4972 ;
  assign n10176 = ( x122 & n4985 ) | ( x122 & n10175 ) | ( n4985 & n10175 ) ;
  assign n10177 = n10175 | n10176 ;
  assign n10178 = x121 & ~n4980 ;
  assign n10179 = ( x121 & n10177 ) | ( x121 & ~n10178 ) | ( n10177 & ~n10178 ) ;
  assign n10180 = ( n4987 & n9806 ) | ( n4987 & n10179 ) | ( n9806 & n10179 ) ;
  assign n10181 = n10179 | n10180 ;
  assign n10182 = n10181 ^ x14 ^ 1'b0 ;
  assign n10183 = n10182 ^ n10173 ^ n9717 ;
  assign n10184 = ( n9717 & n10173 ) | ( n9717 & n10182 ) | ( n10173 & n10182 ) ;
  assign n10185 = x123 & n5499 ;
  assign n10186 = ( x125 & n5497 ) | ( x125 & n10185 ) | ( n5497 & n10185 ) ;
  assign n10187 = n10185 | n10186 ;
  assign n10188 = x124 & ~n5502 ;
  assign n10189 = ( x124 & n10187 ) | ( x124 & ~n10188 ) | ( n10187 & ~n10188 ) ;
  assign n10190 = n5501 & n9883 ;
  assign n10191 = n10189 | n10190 ;
  assign n10192 = n10191 ^ x11 ^ 1'b0 ;
  assign n10193 = ( n10112 & n10183 ) | ( n10112 & n10192 ) | ( n10183 & n10192 ) ;
  assign n10194 = n10192 ^ n10183 ^ n10112 ;
  assign n10195 = x115 & n4790 ;
  assign n10196 = ( x117 & n4792 ) | ( x117 & n10195 ) | ( n4792 & n10195 ) ;
  assign n10197 = n10195 | n10196 ;
  assign n10198 = x116 & ~n4786 ;
  assign n10199 = ( x116 & n10197 ) | ( x116 & ~n10198 ) | ( n10197 & ~n10198 ) ;
  assign n10200 = ( n4787 & n9569 ) | ( n4787 & n10199 ) | ( n9569 & n10199 ) ;
  assign n10201 = n10199 | n10200 ;
  assign n10202 = ( n10146 & n10170 ) | ( n10146 & n10194 ) | ( n10170 & n10194 ) ;
  assign n10203 = n10194 ^ n10170 ^ n10146 ;
  assign n10204 = x118 & n5011 ;
  assign n10205 = ( n10151 & n10153 ) | ( n10151 & n10203 ) | ( n10153 & n10203 ) ;
  assign n10206 = n10203 ^ n10153 ^ n10151 ;
  assign n10207 = ( x120 & n5012 ) | ( x120 & n10204 ) | ( n5012 & n10204 ) ;
  assign n10208 = n10204 | n10207 ;
  assign n10209 = x119 & ~n5008 ;
  assign n10210 = n5020 & n9756 ;
  assign n10211 = n10201 ^ x20 ^ 1'b0 ;
  assign n10212 = ( x119 & n10208 ) | ( x119 & ~n10209 ) | ( n10208 & ~n10209 ) ;
  assign n10213 = n10211 ^ n9409 ^ n9298 ;
  assign n10214 = n10210 | n10212 ;
  assign n10215 = n10214 ^ x17 ^ 1'b0 ;
  assign n10216 = ( n10163 & n10213 ) | ( n10163 & n10215 ) | ( n10213 & n10215 ) ;
  assign n10217 = ( n9298 & n9409 ) | ( n9298 & n10211 ) | ( n9409 & n10211 ) ;
  assign n10218 = n10215 ^ n10213 ^ n10163 ;
  assign n10219 = x121 & n4972 ;
  assign n10220 = ( x123 & n4985 ) | ( x123 & n10219 ) | ( n4985 & n10219 ) ;
  assign n10221 = x122 & ~n4980 ;
  assign n10222 = n10219 | n10220 ;
  assign n10223 = ( x122 & ~n10221 ) | ( x122 & n10222 ) | ( ~n10221 & n10222 ) ;
  assign n10224 = n4987 & n9828 ;
  assign n10225 = n10223 | n10224 ;
  assign n10226 = n10225 ^ x14 ^ 1'b0 ;
  assign n10227 = n10226 ^ n10218 ^ n10174 ;
  assign n10228 = ( n10174 & n10218 ) | ( n10174 & n10226 ) | ( n10218 & n10226 ) ;
  assign n10229 = x116 & n4790 ;
  assign n10230 = ( x118 & n4792 ) | ( x118 & n10229 ) | ( n4792 & n10229 ) ;
  assign n10231 = n10229 | n10230 ;
  assign n10232 = x117 & ~n4786 ;
  assign n10233 = ( x117 & n10231 ) | ( x117 & ~n10232 ) | ( n10231 & ~n10232 ) ;
  assign n10234 = n4787 & n9671 ;
  assign n10235 = n10233 | n10234 ;
  assign n10236 = n10235 ^ x20 ^ 1'b0 ;
  assign n10237 = n10236 ^ n10217 ^ n9441 ;
  assign n10238 = ( n9441 & n10217 ) | ( n9441 & n10236 ) | ( n10217 & n10236 ) ;
  assign n10239 = x124 & n5499 ;
  assign n10240 = ( x126 & n5497 ) | ( x126 & n10239 ) | ( n5497 & n10239 ) ;
  assign n10241 = n10239 | n10240 ;
  assign n10242 = x125 & ~n5502 ;
  assign n10243 = n10126 ^ x8 ^ 1'b0 ;
  assign n10244 = ( x125 & n10241 ) | ( x125 & ~n10242 ) | ( n10241 & ~n10242 ) ;
  assign n10245 = ( n5501 & n9917 ) | ( n5501 & n10244 ) | ( n9917 & n10244 ) ;
  assign n10246 = n10244 | n10245 ;
  assign n10247 = n10246 ^ x11 ^ 1'b0 ;
  assign n10248 = ( n10184 & n10227 ) | ( n10184 & n10247 ) | ( n10227 & n10247 ) ;
  assign n10249 = n10247 ^ n10227 ^ n10184 ;
  assign n10250 = x119 & n5011 ;
  assign n10251 = ( x121 & n5012 ) | ( x121 & n10250 ) | ( n5012 & n10250 ) ;
  assign n10252 = n10250 | n10251 ;
  assign n10253 = x120 & ~n5008 ;
  assign n10254 = ( x120 & n10252 ) | ( x120 & ~n10253 ) | ( n10252 & ~n10253 ) ;
  assign n10255 = n5020 & n9808 ;
  assign n10256 = n10254 | n10255 ;
  assign n10257 = x125 & n5499 ;
  assign n10258 = ( x127 & n5497 ) | ( x127 & n10257 ) | ( n5497 & n10257 ) ;
  assign n10259 = n10257 | n10258 ;
  assign n10260 = n10249 ^ n10243 ^ n10193 ;
  assign n10261 = ( n10193 & n10243 ) | ( n10193 & n10249 ) | ( n10243 & n10249 ) ;
  assign n10262 = x126 & ~n5502 ;
  assign n10263 = ( x126 & n10259 ) | ( x126 & ~n10262 ) | ( n10259 & ~n10262 ) ;
  assign n10264 = n5501 & n9949 ;
  assign n10265 = n10263 | n10264 ;
  assign n10266 = x122 & n4972 ;
  assign n10267 = ( x124 & n4985 ) | ( x124 & n10266 ) | ( n4985 & n10266 ) ;
  assign n10268 = n10266 | n10267 ;
  assign n10269 = x123 & ~n4980 ;
  assign n10270 = ( x123 & n10268 ) | ( x123 & ~n10269 ) | ( n10268 & ~n10269 ) ;
  assign n10271 = n4987 & n9858 ;
  assign n10272 = n10265 ^ x11 ^ 1'b0 ;
  assign n10273 = x127 & ~n5502 ;
  assign n10274 = n10270 | n10271 ;
  assign n10275 = x127 & n5499 ;
  assign n10276 = n10274 ^ x14 ^ 1'b0 ;
  assign n10277 = x126 & n5499 ;
  assign n10278 = ( x127 & ~n10273 ) | ( x127 & n10277 ) | ( ~n10273 & n10277 ) ;
  assign n10279 = ( n5501 & n9958 ) | ( n5501 & n10277 ) | ( n9958 & n10277 ) ;
  assign n10280 = n10256 ^ x17 ^ 1'b0 ;
  assign n10281 = ( n5501 & n9968 ) | ( n5501 & n10275 ) | ( n9968 & n10275 ) ;
  assign n10282 = n10278 | n10279 ;
  assign n10283 = ( n10216 & n10237 ) | ( n10216 & n10280 ) | ( n10237 & n10280 ) ;
  assign n10284 = n10280 ^ n10237 ^ n10216 ;
  assign n10285 = ( n10202 & n10205 ) | ( n10202 & n10260 ) | ( n10205 & n10260 ) ;
  assign n10286 = n10260 ^ n10205 ^ n10202 ;
  assign n10287 = n10275 | n10281 ;
  assign n10288 = ( n10228 & n10276 ) | ( n10228 & n10284 ) | ( n10276 & n10284 ) ;
  assign n10289 = n10284 ^ n10276 ^ n10228 ;
  assign n10290 = n10289 ^ n10272 ^ n10248 ;
  assign n10291 = ( n10261 & n10285 ) | ( n10261 & n10290 ) | ( n10285 & n10290 ) ;
  assign n10292 = ( n10248 & n10272 ) | ( n10248 & n10289 ) | ( n10272 & n10289 ) ;
  assign n10293 = n10290 ^ n10285 ^ n10261 ;
  assign n10294 = x114 & n4616 ;
  assign n10295 = ( x116 & n4606 ) | ( x116 & n10294 ) | ( n4606 & n10294 ) ;
  assign n10296 = n10294 | n10295 ;
  assign n10297 = x115 & ~n4605 ;
  assign n10298 = ( x115 & n10296 ) | ( x115 & ~n10297 ) | ( n10296 & ~n10297 ) ;
  assign n10299 = n4608 & n9513 ;
  assign n10300 = n10298 | n10299 ;
  assign n10301 = n10300 ^ x23 ^ 1'b0 ;
  assign n10302 = ( n9174 & n9318 ) | ( n9174 & n10301 ) | ( n9318 & n10301 ) ;
  assign n10303 = n10301 ^ n9318 ^ n9174 ;
  assign n10304 = x117 & n4790 ;
  assign n10305 = ( x119 & n4792 ) | ( x119 & n10304 ) | ( n4792 & n10304 ) ;
  assign n10306 = n10304 | n10305 ;
  assign n10307 = x118 & ~n4786 ;
  assign n10308 = ( x118 & n10306 ) | ( x118 & ~n10307 ) | ( n10306 & ~n10307 ) ;
  assign n10309 = n4787 & n9733 ;
  assign n10310 = n10308 | n10309 ;
  assign n10311 = n10310 ^ x20 ^ 1'b0 ;
  assign n10312 = ( n9440 & n10303 ) | ( n9440 & n10311 ) | ( n10303 & n10311 ) ;
  assign n10313 = n10311 ^ n10303 ^ n9440 ;
  assign n10314 = x120 & n5011 ;
  assign n10315 = ( x122 & n5012 ) | ( x122 & n10314 ) | ( n5012 & n10314 ) ;
  assign n10316 = n10314 | n10315 ;
  assign n10317 = x121 & ~n5008 ;
  assign n10318 = ( x121 & n10316 ) | ( x121 & ~n10317 ) | ( n10316 & ~n10317 ) ;
  assign n10319 = ( n5020 & n9806 ) | ( n5020 & n10318 ) | ( n9806 & n10318 ) ;
  assign n10320 = n10318 | n10319 ;
  assign n10321 = n10320 ^ x17 ^ 1'b0 ;
  assign n10322 = n10321 ^ n10313 ^ n10238 ;
  assign n10323 = ( n10238 & n10313 ) | ( n10238 & n10321 ) | ( n10313 & n10321 ) ;
  assign n10324 = x123 & n4972 ;
  assign n10325 = ( x125 & n4985 ) | ( x125 & n10324 ) | ( n4985 & n10324 ) ;
  assign n10326 = n10324 | n10325 ;
  assign n10327 = n10282 ^ x11 ^ 1'b0 ;
  assign n10328 = x124 & ~n4980 ;
  assign n10329 = ( x124 & n10326 ) | ( x124 & ~n10328 ) | ( n10326 & ~n10328 ) ;
  assign n10330 = n4987 & n9883 ;
  assign n10331 = n10329 | n10330 ;
  assign n10332 = n10331 ^ x14 ^ 1'b0 ;
  assign n10333 = n10332 ^ n10322 ^ n10283 ;
  assign n10334 = ( n10283 & n10322 ) | ( n10283 & n10332 ) | ( n10322 & n10332 ) ;
  assign n10335 = x126 & ~n4980 ;
  assign n10336 = n10333 ^ n10327 ^ n10288 ;
  assign n10337 = ( n10288 & n10327 ) | ( n10288 & n10333 ) | ( n10327 & n10333 ) ;
  assign n10338 = x125 & n4972 ;
  assign n10339 = ( n10291 & n10292 ) | ( n10291 & n10336 ) | ( n10292 & n10336 ) ;
  assign n10340 = n10336 ^ n10292 ^ n10291 ;
  assign n10341 = ( x127 & n4985 ) | ( x127 & n10338 ) | ( n4985 & n10338 ) ;
  assign n10342 = n4987 & n9949 ;
  assign n10343 = n10338 | n10341 ;
  assign n10344 = ( x126 & ~n10335 ) | ( x126 & n10343 ) | ( ~n10335 & n10343 ) ;
  assign n10345 = n10342 | n10344 ;
  assign n10346 = x116 & ~n4605 ;
  assign n10347 = x115 & n4616 ;
  assign n10348 = ( x117 & n4606 ) | ( x117 & n10347 ) | ( n4606 & n10347 ) ;
  assign n10349 = n10347 | n10348 ;
  assign n10350 = x127 & ~n4980 ;
  assign n10351 = ( x116 & ~n10346 ) | ( x116 & n10349 ) | ( ~n10346 & n10349 ) ;
  assign n10352 = x125 & ~n4980 ;
  assign n10353 = x126 & n4972 ;
  assign n10354 = ( x127 & ~n10350 ) | ( x127 & n10353 ) | ( ~n10350 & n10353 ) ;
  assign n10355 = ( n4987 & n9958 ) | ( n4987 & n10353 ) | ( n9958 & n10353 ) ;
  assign n10356 = n10354 | n10355 ;
  assign n10357 = ( n4608 & n9569 ) | ( n4608 & n10351 ) | ( n9569 & n10351 ) ;
  assign n10358 = n10351 | n10357 ;
  assign n10359 = n10358 ^ x23 ^ 1'b0 ;
  assign n10360 = x124 & n4972 ;
  assign n10361 = ( x126 & n4985 ) | ( x126 & n10360 ) | ( n4985 & n10360 ) ;
  assign n10362 = x127 & n4972 ;
  assign n10363 = n10360 | n10361 ;
  assign n10364 = ( x125 & ~n10352 ) | ( x125 & n10363 ) | ( ~n10352 & n10363 ) ;
  assign n10365 = ( n4987 & n9968 ) | ( n4987 & n10362 ) | ( n9968 & n10362 ) ;
  assign n10366 = ( n4987 & n9917 ) | ( n4987 & n10364 ) | ( n9917 & n10364 ) ;
  assign n10367 = ( n9319 & n9378 ) | ( n9319 & n10359 ) | ( n9378 & n10359 ) ;
  assign n10368 = n10362 | n10365 ;
  assign n10369 = n10359 ^ n9378 ^ n9319 ;
  assign n10370 = n10364 | n10366 ;
  assign n10371 = x118 & n4790 ;
  assign n10372 = ( x120 & n4792 ) | ( x120 & n10371 ) | ( n4792 & n10371 ) ;
  assign n10373 = n10371 | n10372 ;
  assign n10374 = x119 & ~n4786 ;
  assign n10375 = ( x119 & n10373 ) | ( x119 & ~n10374 ) | ( n10373 & ~n10374 ) ;
  assign n10376 = n4787 & n9756 ;
  assign n10377 = n10375 | n10376 ;
  assign n10378 = n10377 ^ x20 ^ 1'b0 ;
  assign n10379 = n10378 ^ n10369 ^ n10302 ;
  assign n10380 = ( n10302 & n10369 ) | ( n10302 & n10378 ) | ( n10369 & n10378 ) ;
  assign n10381 = x121 & n5011 ;
  assign n10382 = ( x123 & n5012 ) | ( x123 & n10381 ) | ( n5012 & n10381 ) ;
  assign n10383 = n10381 | n10382 ;
  assign n10384 = x122 & ~n5008 ;
  assign n10385 = ( x122 & n10383 ) | ( x122 & ~n10384 ) | ( n10383 & ~n10384 ) ;
  assign n10386 = n5020 & n9828 ;
  assign n10387 = n10385 | n10386 ;
  assign n10388 = n10370 ^ x14 ^ 1'b0 ;
  assign n10389 = n10387 ^ x17 ^ 1'b0 ;
  assign n10390 = n10287 ^ x11 ^ 1'b0 ;
  assign n10391 = ( n10312 & n10379 ) | ( n10312 & n10389 ) | ( n10379 & n10389 ) ;
  assign n10392 = n10389 ^ n10379 ^ n10312 ;
  assign n10393 = n10392 ^ n10388 ^ n10323 ;
  assign n10394 = ( n10334 & n10390 ) | ( n10334 & n10393 ) | ( n10390 & n10393 ) ;
  assign n10395 = n10393 ^ n10390 ^ n10334 ;
  assign n10396 = x117 & ~n4605 ;
  assign n10397 = ( n10323 & n10388 ) | ( n10323 & n10392 ) | ( n10388 & n10392 ) ;
  assign n10398 = x119 & n4790 ;
  assign n10399 = ( x121 & n4792 ) | ( x121 & n10398 ) | ( n4792 & n10398 ) ;
  assign n10400 = x116 & n4616 ;
  assign n10401 = n10398 | n10399 ;
  assign n10402 = ( x118 & n4606 ) | ( x118 & n10400 ) | ( n4606 & n10400 ) ;
  assign n10403 = n10400 | n10402 ;
  assign n10404 = n10395 ^ n10339 ^ n10337 ;
  assign n10405 = ( n10337 & n10339 ) | ( n10337 & n10395 ) | ( n10339 & n10395 ) ;
  assign n10406 = n4787 & n9808 ;
  assign n10407 = ( x117 & ~n10396 ) | ( x117 & n10403 ) | ( ~n10396 & n10403 ) ;
  assign n10408 = x123 & ~n5008 ;
  assign n10409 = n4608 & n9671 ;
  assign n10410 = n10345 ^ x14 ^ 1'b0 ;
  assign n10411 = n10407 | n10409 ;
  assign n10412 = n10411 ^ x23 ^ 1'b0 ;
  assign n10413 = x120 & ~n4786 ;
  assign n10414 = ( x120 & n10401 ) | ( x120 & ~n10413 ) | ( n10401 & ~n10413 ) ;
  assign n10415 = n10412 ^ n10367 ^ n9450 ;
  assign n10416 = n10406 | n10414 ;
  assign n10417 = n10416 ^ x20 ^ 1'b0 ;
  assign n10418 = ( n10380 & n10415 ) | ( n10380 & n10417 ) | ( n10415 & n10417 ) ;
  assign n10419 = ( n9450 & n10367 ) | ( n9450 & n10412 ) | ( n10367 & n10412 ) ;
  assign n10420 = n10417 ^ n10415 ^ n10380 ;
  assign n10421 = x122 & n5011 ;
  assign n10422 = ( x124 & n5012 ) | ( x124 & n10421 ) | ( n5012 & n10421 ) ;
  assign n10423 = n10421 | n10422 ;
  assign n10424 = ( x123 & ~n10408 ) | ( x123 & n10423 ) | ( ~n10408 & n10423 ) ;
  assign n10425 = n5020 & n9858 ;
  assign n10426 = n10424 | n10425 ;
  assign n10427 = n10426 ^ x17 ^ 1'b0 ;
  assign n10428 = n10427 ^ n10420 ^ n10391 ;
  assign n10429 = n10428 ^ n10410 ^ n10397 ;
  assign n10430 = ( n10397 & n10410 ) | ( n10397 & n10428 ) | ( n10410 & n10428 ) ;
  assign n10431 = n10429 ^ n10405 ^ n10394 ;
  assign n10432 = ( n10394 & n10405 ) | ( n10394 & n10429 ) | ( n10405 & n10429 ) ;
  assign n10433 = ( n10391 & n10420 ) | ( n10391 & n10427 ) | ( n10420 & n10427 ) ;
  assign n10434 = x114 & n3734 ;
  assign n10435 = ( x116 & n3732 ) | ( x116 & n10434 ) | ( n3732 & n10434 ) ;
  assign n10436 = n10434 | n10435 ;
  assign n10437 = x125 & n5011 ;
  assign n10438 = ( x127 & n5012 ) | ( x127 & n10437 ) | ( n5012 & n10437 ) ;
  assign n10439 = x115 & ~n3737 ;
  assign n10440 = ( x115 & n10436 ) | ( x115 & ~n10439 ) | ( n10436 & ~n10439 ) ;
  assign n10441 = ( n3736 & n9513 ) | ( n3736 & n10440 ) | ( n9513 & n10440 ) ;
  assign n10442 = n10440 | n10441 ;
  assign n10443 = n10442 ^ x26 ^ 1'b0 ;
  assign n10444 = x124 & ~n5008 ;
  assign n10445 = n10443 ^ n9278 ^ n9090 ;
  assign n10446 = n10437 | n10438 ;
  assign n10447 = x126 & ~n5008 ;
  assign n10448 = ( x126 & n10446 ) | ( x126 & ~n10447 ) | ( n10446 & ~n10447 ) ;
  assign n10449 = x123 & n5011 ;
  assign n10450 = ( n9090 & n9278 ) | ( n9090 & n10443 ) | ( n9278 & n10443 ) ;
  assign n10451 = ( x125 & n5012 ) | ( x125 & n10449 ) | ( n5012 & n10449 ) ;
  assign n10452 = x127 & n5011 ;
  assign n10453 = n10449 | n10451 ;
  assign n10454 = x127 & ~n5008 ;
  assign n10455 = ( x124 & ~n10444 ) | ( x124 & n10453 ) | ( ~n10444 & n10453 ) ;
  assign n10456 = x124 & n5011 ;
  assign n10457 = x126 & n5011 ;
  assign n10458 = n10368 ^ x14 ^ 1'b0 ;
  assign n10459 = n10356 ^ x14 ^ 1'b0 ;
  assign n10460 = x125 & ~n5008 ;
  assign n10461 = ( x126 & n5012 ) | ( x126 & n10456 ) | ( n5012 & n10456 ) ;
  assign n10462 = n10456 | n10461 ;
  assign n10463 = n5020 & n9949 ;
  assign n10464 = ( x125 & ~n10460 ) | ( x125 & n10462 ) | ( ~n10460 & n10462 ) ;
  assign n10465 = ( n5020 & n9917 ) | ( n5020 & n10464 ) | ( n9917 & n10464 ) ;
  assign n10466 = ( x127 & ~n10454 ) | ( x127 & n10457 ) | ( ~n10454 & n10457 ) ;
  assign n10467 = n10464 | n10465 ;
  assign n10468 = ( n5020 & n9968 ) | ( n5020 & n10452 ) | ( n9968 & n10452 ) ;
  assign n10469 = ( n5020 & n9958 ) | ( n5020 & n10457 ) | ( n9958 & n10457 ) ;
  assign n10470 = n5020 & n9883 ;
  assign n10471 = n10455 | n10470 ;
  assign n10472 = n10452 | n10468 ;
  assign n10473 = x117 & n4616 ;
  assign n10474 = ( x119 & n4606 ) | ( x119 & n10473 ) | ( n4606 & n10473 ) ;
  assign n10475 = n10473 | n10474 ;
  assign n10476 = n10448 | n10463 ;
  assign n10477 = x120 & n4790 ;
  assign n10478 = ( x122 & n4792 ) | ( x122 & n10477 ) | ( n4792 & n10477 ) ;
  assign n10479 = n10477 | n10478 ;
  assign n10480 = x118 & ~n4605 ;
  assign n10481 = ( x118 & n10475 ) | ( x118 & ~n10480 ) | ( n10475 & ~n10480 ) ;
  assign n10482 = n10466 | n10469 ;
  assign n10483 = x121 & ~n4786 ;
  assign n10484 = ( x121 & n10479 ) | ( x121 & ~n10483 ) | ( n10479 & ~n10483 ) ;
  assign n10485 = ( n4787 & n9806 ) | ( n4787 & n10484 ) | ( n9806 & n10484 ) ;
  assign n10486 = n10484 | n10485 ;
  assign n10487 = n4608 & n9733 ;
  assign n10488 = n10481 | n10487 ;
  assign n10489 = n10488 ^ x23 ^ 1'b0 ;
  assign n10490 = n10486 ^ x20 ^ 1'b0 ;
  assign n10491 = n10489 ^ n10445 ^ n9451 ;
  assign n10492 = n10471 ^ x17 ^ 1'b0 ;
  assign n10493 = ( n10419 & n10490 ) | ( n10419 & n10491 ) | ( n10490 & n10491 ) ;
  assign n10494 = n10491 ^ n10490 ^ n10419 ;
  assign n10495 = ( n9451 & n10445 ) | ( n9451 & n10489 ) | ( n10445 & n10489 ) ;
  assign n10496 = ( n10418 & n10492 ) | ( n10418 & n10494 ) | ( n10492 & n10494 ) ;
  assign n10497 = n10494 ^ n10492 ^ n10418 ;
  assign n10498 = n10497 ^ n10459 ^ n10433 ;
  assign n10499 = ( n10430 & n10432 ) | ( n10430 & n10498 ) | ( n10432 & n10498 ) ;
  assign n10500 = ( n10433 & n10459 ) | ( n10433 & n10497 ) | ( n10459 & n10497 ) ;
  assign n10501 = n10498 ^ n10432 ^ n10430 ;
  assign n10502 = x118 & n4616 ;
  assign n10503 = ( x120 & n4606 ) | ( x120 & n10502 ) | ( n4606 & n10502 ) ;
  assign n10504 = n10502 | n10503 ;
  assign n10505 = x119 & ~n4605 ;
  assign n10506 = ( x119 & n10504 ) | ( x119 & ~n10505 ) | ( n10504 & ~n10505 ) ;
  assign n10507 = n4608 & n9756 ;
  assign n10508 = n10506 | n10507 ;
  assign n10509 = n10508 ^ x23 ^ 1'b0 ;
  assign n10510 = n10509 ^ n10450 ^ n9634 ;
  assign n10511 = ( n9634 & n10450 ) | ( n9634 & n10509 ) | ( n10450 & n10509 ) ;
  assign n10512 = x121 & n4790 ;
  assign n10513 = ( x123 & n4792 ) | ( x123 & n10512 ) | ( n4792 & n10512 ) ;
  assign n10514 = n10512 | n10513 ;
  assign n10515 = x122 & ~n4786 ;
  assign n10516 = ( x122 & n10514 ) | ( x122 & ~n10515 ) | ( n10514 & ~n10515 ) ;
  assign n10517 = n4787 & n9828 ;
  assign n10518 = n10516 | n10517 ;
  assign n10519 = n10518 ^ x20 ^ 1'b0 ;
  assign n10520 = ( n10495 & n10510 ) | ( n10495 & n10519 ) | ( n10510 & n10519 ) ;
  assign n10521 = n10519 ^ n10510 ^ n10495 ;
  assign n10522 = n10467 ^ x17 ^ 1'b0 ;
  assign n10523 = n10522 ^ n10521 ^ n10493 ;
  assign n10524 = ( n10493 & n10521 ) | ( n10493 & n10522 ) | ( n10521 & n10522 ) ;
  assign n10525 = x116 & n3734 ;
  assign n10526 = ( x118 & n3732 ) | ( x118 & n10525 ) | ( n3732 & n10525 ) ;
  assign n10527 = n10525 | n10526 ;
  assign n10528 = x117 & ~n3737 ;
  assign n10529 = ( x117 & n10527 ) | ( x117 & ~n10528 ) | ( n10527 & ~n10528 ) ;
  assign n10530 = n3736 & n9671 ;
  assign n10531 = n10529 | n10530 ;
  assign n10532 = n10531 ^ x26 ^ 1'b0 ;
  assign n10533 = ( n9420 & n9635 ) | ( n9420 & n10532 ) | ( n9635 & n10532 ) ;
  assign n10534 = n10532 ^ n9635 ^ n9420 ;
  assign n10535 = n10523 ^ n10496 ^ n10458 ;
  assign n10536 = x122 & n4790 ;
  assign n10537 = ( x124 & n4792 ) | ( x124 & n10536 ) | ( n4792 & n10536 ) ;
  assign n10538 = n10536 | n10537 ;
  assign n10539 = x123 & ~n4786 ;
  assign n10540 = ( x123 & n10538 ) | ( x123 & ~n10539 ) | ( n10538 & ~n10539 ) ;
  assign n10541 = n10535 ^ n10500 ^ n10499 ;
  assign n10542 = ( n10499 & n10500 ) | ( n10499 & n10535 ) | ( n10500 & n10535 ) ;
  assign n10543 = n4787 & n9858 ;
  assign n10544 = n10476 ^ x17 ^ 1'b0 ;
  assign n10545 = x120 & ~n4605 ;
  assign n10546 = n10540 | n10543 ;
  assign n10547 = ( n10458 & n10496 ) | ( n10458 & n10523 ) | ( n10496 & n10523 ) ;
  assign n10548 = n4608 & n9808 ;
  assign n10549 = x119 & n4616 ;
  assign n10550 = n10546 ^ x20 ^ 1'b0 ;
  assign n10551 = ( x121 & n4606 ) | ( x121 & n10549 ) | ( n4606 & n10549 ) ;
  assign n10552 = n10549 | n10551 ;
  assign n10553 = ( x120 & ~n10545 ) | ( x120 & n10552 ) | ( ~n10545 & n10552 ) ;
  assign n10554 = n10548 | n10553 ;
  assign n10555 = n10554 ^ x23 ^ 1'b0 ;
  assign n10556 = n10555 ^ n10534 ^ n10511 ;
  assign n10557 = n10556 ^ n10550 ^ n10520 ;
  assign n10558 = ( n10524 & n10544 ) | ( n10524 & n10557 ) | ( n10544 & n10557 ) ;
  assign n10559 = n10557 ^ n10544 ^ n10524 ;
  assign n10560 = ( n10511 & n10534 ) | ( n10511 & n10555 ) | ( n10534 & n10555 ) ;
  assign n10561 = ( n10520 & n10550 ) | ( n10520 & n10556 ) | ( n10550 & n10556 ) ;
  assign n10562 = ( n10542 & n10547 ) | ( n10542 & n10559 ) | ( n10547 & n10559 ) ;
  assign n10563 = n10559 ^ n10547 ^ n10542 ;
  assign n10564 = x114 & n3344 ;
  assign n10565 = n3346 & n9513 ;
  assign n10566 = x115 & n3344 ;
  assign n10567 = ( x116 & n3342 ) | ( x116 & n10564 ) | ( n3342 & n10564 ) ;
  assign n10568 = n10564 | n10567 ;
  assign n10569 = x115 & ~n3347 ;
  assign n10570 = ( x115 & n10568 ) | ( x115 & ~n10569 ) | ( n10568 & ~n10569 ) ;
  assign n10571 = ( x117 & n3342 ) | ( x117 & n10566 ) | ( n3342 & n10566 ) ;
  assign n10572 = n10566 | n10571 ;
  assign n10573 = x117 & n3734 ;
  assign n10574 = n10565 | n10570 ;
  assign n10575 = ( x119 & n3732 ) | ( x119 & n10573 ) | ( n3732 & n10573 ) ;
  assign n10576 = n10573 | n10575 ;
  assign n10577 = x116 & ~n3347 ;
  assign n10578 = n10574 ^ x29 ^ 1'b0 ;
  assign n10579 = ( x116 & n10572 ) | ( x116 & ~n10577 ) | ( n10572 & ~n10577 ) ;
  assign n10580 = n10578 ^ n9328 ^ n9135 ;
  assign n10581 = n10482 ^ x17 ^ 1'b0 ;
  assign n10582 = ( n9135 & n9328 ) | ( n9135 & n10578 ) | ( n9328 & n10578 ) ;
  assign n10583 = n3346 & n9569 ;
  assign n10584 = x118 & ~n3737 ;
  assign n10585 = n10579 | n10583 ;
  assign n10586 = ( x118 & n10576 ) | ( x118 & ~n10584 ) | ( n10576 & ~n10584 ) ;
  assign n10587 = n3736 & n9733 ;
  assign n10588 = n10586 | n10587 ;
  assign n10589 = n10585 ^ x29 ^ 1'b0 ;
  assign n10590 = x118 & n3734 ;
  assign n10591 = ( x120 & n3732 ) | ( x120 & n10590 ) | ( n3732 & n10590 ) ;
  assign n10592 = n10590 | n10591 ;
  assign n10593 = ( n9329 & n9400 ) | ( n9329 & n10589 ) | ( n9400 & n10589 ) ;
  assign n10594 = n10589 ^ n9400 ^ n9329 ;
  assign n10595 = x120 & n4616 ;
  assign n10596 = ( x122 & n4606 ) | ( x122 & n10595 ) | ( n4606 & n10595 ) ;
  assign n10597 = n10588 ^ x26 ^ 1'b0 ;
  assign n10598 = n10595 | n10596 ;
  assign n10599 = x119 & ~n3737 ;
  assign n10600 = ( x119 & n10592 ) | ( x119 & ~n10599 ) | ( n10592 & ~n10599 ) ;
  assign n10601 = n3736 & n9756 ;
  assign n10602 = n10600 | n10601 ;
  assign n10603 = ( n9419 & n10580 ) | ( n9419 & n10597 ) | ( n10580 & n10597 ) ;
  assign n10604 = n10602 ^ x26 ^ 1'b0 ;
  assign n10605 = n10597 ^ n10580 ^ n9419 ;
  assign n10606 = ( n10582 & n10594 ) | ( n10582 & n10604 ) | ( n10594 & n10604 ) ;
  assign n10607 = n10604 ^ n10594 ^ n10582 ;
  assign n10608 = x121 & n4616 ;
  assign n10609 = ( x123 & n4606 ) | ( x123 & n10608 ) | ( n4606 & n10608 ) ;
  assign n10610 = n10608 | n10609 ;
  assign n10611 = x122 & ~n4605 ;
  assign n10612 = x121 & ~n4605 ;
  assign n10613 = ( x121 & n10598 ) | ( x121 & ~n10612 ) | ( n10598 & ~n10612 ) ;
  assign n10614 = x123 & n4790 ;
  assign n10615 = ( x122 & n10610 ) | ( x122 & ~n10611 ) | ( n10610 & ~n10611 ) ;
  assign n10616 = ( x125 & n4792 ) | ( x125 & n10614 ) | ( n4792 & n10614 ) ;
  assign n10617 = n10614 | n10616 ;
  assign n10618 = ( n4608 & n9806 ) | ( n4608 & n10613 ) | ( n9806 & n10613 ) ;
  assign n10619 = n10613 | n10618 ;
  assign n10620 = n10619 ^ x23 ^ 1'b0 ;
  assign n10621 = n10620 ^ n10605 ^ n10533 ;
  assign n10622 = ( n10533 & n10605 ) | ( n10533 & n10620 ) | ( n10605 & n10620 ) ;
  assign n10623 = x124 & ~n4786 ;
  assign n10624 = n4787 & n9883 ;
  assign n10625 = ( x124 & n10617 ) | ( x124 & ~n10623 ) | ( n10617 & ~n10623 ) ;
  assign n10626 = n4608 & n9828 ;
  assign n10627 = n10624 | n10625 ;
  assign n10628 = n10615 | n10626 ;
  assign n10629 = n10628 ^ x23 ^ 1'b0 ;
  assign n10630 = n10629 ^ n10607 ^ n10603 ;
  assign n10631 = n10627 ^ x20 ^ 1'b0 ;
  assign n10632 = ( n10560 & n10621 ) | ( n10560 & n10631 ) | ( n10621 & n10631 ) ;
  assign n10633 = n10631 ^ n10621 ^ n10560 ;
  assign n10634 = ( n10561 & n10581 ) | ( n10561 & n10633 ) | ( n10581 & n10633 ) ;
  assign n10635 = n10633 ^ n10581 ^ n10561 ;
  assign n10636 = ( n10558 & n10562 ) | ( n10558 & n10635 ) | ( n10562 & n10635 ) ;
  assign n10637 = ( n10603 & n10607 ) | ( n10603 & n10629 ) | ( n10607 & n10629 ) ;
  assign n10638 = n10635 ^ n10562 ^ n10558 ;
  assign n10639 = x124 & n4790 ;
  assign n10640 = ( x126 & n4792 ) | ( x126 & n10639 ) | ( n4792 & n10639 ) ;
  assign n10641 = n10639 | n10640 ;
  assign n10642 = x125 & ~n4786 ;
  assign n10643 = ( x125 & n10641 ) | ( x125 & ~n10642 ) | ( n10641 & ~n10642 ) ;
  assign n10644 = n4787 & n9917 ;
  assign n10645 = n10643 | n10644 ;
  assign n10646 = n10472 ^ x17 ^ 1'b0 ;
  assign n10647 = n10645 ^ x20 ^ 1'b0 ;
  assign n10648 = ( n10622 & n10630 ) | ( n10622 & n10647 ) | ( n10630 & n10647 ) ;
  assign n10649 = n10647 ^ n10630 ^ n10622 ;
  assign n10650 = n10649 ^ n10646 ^ n10632 ;
  assign n10651 = n10650 ^ n10636 ^ n10634 ;
  assign n10652 = ( n10634 & n10636 ) | ( n10634 & n10650 ) | ( n10636 & n10650 ) ;
  assign n10653 = x119 & n3734 ;
  assign n10654 = ( x121 & n3732 ) | ( x121 & n10653 ) | ( n3732 & n10653 ) ;
  assign n10655 = n10653 | n10654 ;
  assign n10656 = n3736 & n9808 ;
  assign n10657 = ( n10632 & n10646 ) | ( n10632 & n10649 ) | ( n10646 & n10649 ) ;
  assign n10658 = x120 & ~n3737 ;
  assign n10659 = x127 & n4790 ;
  assign n10660 = ( x120 & n10655 ) | ( x120 & ~n10658 ) | ( n10655 & ~n10658 ) ;
  assign n10661 = n10656 | n10660 ;
  assign n10662 = n10661 ^ x26 ^ 1'b0 ;
  assign n10663 = x127 & ~n4786 ;
  assign n10664 = x125 & n4790 ;
  assign n10665 = x126 & ~n4786 ;
  assign n10666 = ( x127 & n4792 ) | ( x127 & n10664 ) | ( n4792 & n10664 ) ;
  assign n10667 = n10664 | n10666 ;
  assign n10668 = ( x126 & ~n10665 ) | ( x126 & n10667 ) | ( ~n10665 & n10667 ) ;
  assign n10669 = ( n4787 & n9968 ) | ( n4787 & n10659 ) | ( n9968 & n10659 ) ;
  assign n10670 = x126 & n4790 ;
  assign n10671 = ( x127 & ~n10663 ) | ( x127 & n10670 ) | ( ~n10663 & n10670 ) ;
  assign n10672 = x122 & n4616 ;
  assign n10673 = n10659 | n10669 ;
  assign n10674 = ( x124 & n4606 ) | ( x124 & n10672 ) | ( n4606 & n10672 ) ;
  assign n10675 = n10672 | n10674 ;
  assign n10676 = x123 & ~n4605 ;
  assign n10677 = ( x123 & n10675 ) | ( x123 & ~n10676 ) | ( n10675 & ~n10676 ) ;
  assign n10678 = n4608 & n9858 ;
  assign n10679 = n10677 | n10678 ;
  assign n10680 = ( n4787 & n9958 ) | ( n4787 & n10670 ) | ( n9958 & n10670 ) ;
  assign n10681 = n10671 | n10680 ;
  assign n10682 = n10681 ^ x20 ^ 1'b0 ;
  assign n10683 = x116 & n3344 ;
  assign n10684 = ( x118 & n3342 ) | ( x118 & n10683 ) | ( n3342 & n10683 ) ;
  assign n10685 = n10679 ^ x23 ^ 1'b0 ;
  assign n10686 = n4787 & n9949 ;
  assign n10687 = n10668 | n10686 ;
  assign n10688 = x117 & ~n3347 ;
  assign n10689 = n10683 | n10684 ;
  assign n10690 = n3346 & n9671 ;
  assign n10691 = ( x117 & ~n10688 ) | ( x117 & n10689 ) | ( ~n10688 & n10689 ) ;
  assign n10692 = n10690 | n10691 ;
  assign n10693 = n10692 ^ x29 ^ 1'b0 ;
  assign n10694 = ( n9431 & n10593 ) | ( n9431 & n10693 ) | ( n10593 & n10693 ) ;
  assign n10695 = n10687 ^ x20 ^ 1'b0 ;
  assign n10696 = n10693 ^ n10593 ^ n9431 ;
  assign n10697 = n10696 ^ n10662 ^ n10606 ;
  assign n10698 = n10697 ^ n10685 ^ n10637 ;
  assign n10699 = ( n10606 & n10662 ) | ( n10606 & n10696 ) | ( n10662 & n10696 ) ;
  assign n10700 = n10698 ^ n10695 ^ n10648 ;
  assign n10701 = ( n10637 & n10685 ) | ( n10637 & n10697 ) | ( n10685 & n10697 ) ;
  assign n10702 = n10700 ^ n10657 ^ n10652 ;
  assign n10703 = ( n10648 & n10695 ) | ( n10648 & n10698 ) | ( n10695 & n10698 ) ;
  assign n10704 = ( n10652 & n10657 ) | ( n10652 & n10700 ) | ( n10657 & n10700 ) ;
  assign n10705 = x87 & n133 ;
  assign n10706 = ( x89 & n142 ) | ( x89 & n10705 ) | ( n142 & n10705 ) ;
  assign n10707 = n10705 | n10706 ;
  assign n10708 = x88 & ~n134 ;
  assign n10709 = ( x88 & n10707 ) | ( x88 & ~n10708 ) | ( n10707 & ~n10708 ) ;
  assign n10710 = x83 & ~n242 ;
  assign n10711 = x82 & n325 ;
  assign n10712 = ( x83 & ~n10710 ) | ( x83 & n10711 ) | ( ~n10710 & n10711 ) ;
  assign n10713 = n140 & n1654 ;
  assign n10714 = n10709 | n10713 ;
  assign n10715 = n10714 ^ x59 ^ 1'b0 ;
  assign n10716 = ( n4551 & n7874 ) | ( n4551 & ~n10712 ) | ( n7874 & ~n10712 ) ;
  assign n10717 = n10712 ^ n7874 ^ n4551 ;
  assign n10718 = n10717 ^ n10715 ^ n4553 ;
  assign n10719 = ( n4553 & n10715 ) | ( n4553 & ~n10717 ) | ( n10715 & ~n10717 ) ;
  assign n10720 = x90 & n263 ;
  assign n10721 = ( x92 & n264 ) | ( x92 & n10720 ) | ( n264 & n10720 ) ;
  assign n10722 = n10720 | n10721 ;
  assign n10723 = x91 & ~n260 ;
  assign n10724 = ( x91 & n10722 ) | ( x91 & ~n10723 ) | ( n10722 & ~n10723 ) ;
  assign n10725 = n272 & n2420 ;
  assign n10726 = n10724 | n10725 ;
  assign n10727 = n10726 ^ x56 ^ 1'b0 ;
  assign n10728 = n10727 ^ n10718 ^ n4563 ;
  assign n10729 = ( n4563 & ~n10718 ) | ( n4563 & n10727 ) | ( ~n10718 & n10727 ) ;
  assign n10730 = x93 & n408 ;
  assign n10731 = ( x95 & n403 ) | ( x95 & n10730 ) | ( n403 & n10730 ) ;
  assign n10732 = n10730 | n10731 ;
  assign n10733 = x94 & ~n410 ;
  assign n10734 = ( x94 & n10732 ) | ( x94 & ~n10733 ) | ( n10732 & ~n10733 ) ;
  assign n10735 = n402 & n2854 ;
  assign n10736 = n10734 | n10735 ;
  assign n10737 = n10736 ^ x53 ^ 1'b0 ;
  assign n10738 = ( n4574 & ~n10728 ) | ( n4574 & n10737 ) | ( ~n10728 & n10737 ) ;
  assign n10739 = n10737 ^ n10728 ^ n4574 ;
  assign n10740 = x96 & n561 ;
  assign n10741 = ( x98 & n551 ) | ( x98 & n10740 ) | ( n551 & n10740 ) ;
  assign n10742 = n10740 | n10741 ;
  assign n10743 = x97 & ~n550 ;
  assign n10744 = ( x97 & n10742 ) | ( x97 & ~n10743 ) | ( n10742 & ~n10743 ) ;
  assign n10745 = n553 & n4052 ;
  assign n10746 = n10744 | n10745 ;
  assign n10747 = n10746 ^ x50 ^ 1'b0 ;
  assign n10748 = ( n4588 & ~n10739 ) | ( n4588 & n10747 ) | ( ~n10739 & n10747 ) ;
  assign n10749 = n10747 ^ n10739 ^ n4588 ;
  assign n10750 = x99 & n744 ;
  assign n10751 = ( x101 & n730 ) | ( x101 & n10750 ) | ( n730 & n10750 ) ;
  assign n10752 = n10750 | n10751 ;
  assign n10753 = x100 & ~n732 ;
  assign n10754 = ( x100 & n10752 ) | ( x100 & ~n10753 ) | ( n10752 & ~n10753 ) ;
  assign n10755 = n731 & n5687 ;
  assign n10756 = n10754 | n10755 ;
  assign n10757 = n10756 ^ x47 ^ 1'b0 ;
  assign n10758 = n10757 ^ n10749 ^ n4599 ;
  assign n10759 = ( n4599 & ~n10749 ) | ( n4599 & n10757 ) | ( ~n10749 & n10757 ) ;
  assign n10760 = x85 & n208 ;
  assign n10761 = ( x87 & n194 ) | ( x87 & n10760 ) | ( n194 & n10760 ) ;
  assign n10762 = n10760 | n10761 ;
  assign n10763 = x86 & ~n192 ;
  assign n10764 = ( x86 & n10762 ) | ( x86 & ~n10763 ) | ( n10762 & ~n10763 ) ;
  assign n10765 = ( n197 & n1484 ) | ( n197 & n10764 ) | ( n1484 & n10764 ) ;
  assign n10766 = x102 & n888 ;
  assign n10767 = n10764 | n10765 ;
  assign n10768 = ( x104 & n878 ) | ( x104 & n10766 ) | ( n878 & n10766 ) ;
  assign n10769 = n10766 | n10768 ;
  assign n10770 = x103 & ~n877 ;
  assign n10771 = n10767 ^ x62 ^ 1'b0 ;
  assign n10772 = ( x103 & n10769 ) | ( x103 & ~n10770 ) | ( n10769 & ~n10770 ) ;
  assign n10773 = n880 & n8012 ;
  assign n10774 = n10772 | n10773 ;
  assign n10775 = n10774 ^ x44 ^ 1'b0 ;
  assign n10776 = ( n4601 & ~n10758 ) | ( n4601 & n10775 ) | ( ~n10758 & n10775 ) ;
  assign n10777 = n10775 ^ n10758 ^ n4601 ;
  assign n10778 = x105 & n1058 ;
  assign n10779 = ( x107 & n1065 ) | ( x107 & n10778 ) | ( n1065 & n10778 ) ;
  assign n10780 = n10778 | n10779 ;
  assign n10781 = x106 & ~n1060 ;
  assign n10782 = ( x106 & n10780 ) | ( x106 & ~n10781 ) | ( n10780 & ~n10781 ) ;
  assign n10783 = n1063 & n8440 ;
  assign n10784 = n10782 | n10783 ;
  assign n10785 = n10784 ^ x41 ^ 1'b0 ;
  assign n10786 = n10785 ^ n10777 ^ n7875 ;
  assign n10787 = ( n7875 & n10777 ) | ( n7875 & ~n10785 ) | ( n10777 & ~n10785 ) ;
  assign n10788 = x108 & n2156 ;
  assign n10789 = ( x110 & n2163 ) | ( x110 & n10788 ) | ( n2163 & n10788 ) ;
  assign n10790 = n10788 | n10789 ;
  assign n10791 = x109 & ~n2158 ;
  assign n10792 = ( x109 & n10790 ) | ( x109 & ~n10791 ) | ( n10790 & ~n10791 ) ;
  assign n10793 = n2161 & n8820 ;
  assign n10794 = n10792 | n10793 ;
  assign n10795 = n10794 ^ x38 ^ 1'b0 ;
  assign n10796 = n10795 ^ n10786 ^ n8292 ;
  assign n10797 = ( n8292 & n10786 ) | ( n8292 & n10795 ) | ( n10786 & n10795 ) ;
  assign n10798 = x111 & n2560 ;
  assign n10799 = ( x113 & n2567 ) | ( x113 & n10798 ) | ( n2567 & n10798 ) ;
  assign n10800 = n10798 | n10799 ;
  assign n10801 = x112 & ~n2562 ;
  assign n10802 = ( x112 & n10800 ) | ( x112 & ~n10801 ) | ( n10800 & ~n10801 ) ;
  assign n10803 = n2565 & n9199 ;
  assign n10804 = n10802 | n10803 ;
  assign n10805 = n10804 ^ x35 ^ 1'b0 ;
  assign n10806 = n10805 ^ n10796 ^ n8921 ;
  assign n10807 = ( n8921 & n10796 ) | ( n8921 & n10805 ) | ( n10796 & n10805 ) ;
  assign n10808 = x114 & n3025 ;
  assign n10809 = ( x116 & n3015 ) | ( x116 & n10808 ) | ( n3015 & n10808 ) ;
  assign n10810 = n10808 | n10809 ;
  assign n10811 = x115 & ~n3014 ;
  assign n10812 = ( x115 & n10810 ) | ( x115 & ~n10811 ) | ( n10810 & ~n10811 ) ;
  assign n10813 = n3017 & n9513 ;
  assign n10814 = n10812 | n10813 ;
  assign n10815 = n10814 ^ x32 ^ 1'b0 ;
  assign n10816 = n10815 ^ n10806 ^ n9105 ;
  assign n10817 = ( n9105 & n10806 ) | ( n9105 & n10815 ) | ( n10806 & n10815 ) ;
  assign n10818 = x117 & n3344 ;
  assign n10819 = ( x119 & n3342 ) | ( x119 & n10818 ) | ( n3342 & n10818 ) ;
  assign n10820 = n10818 | n10819 ;
  assign n10821 = x118 & ~n3347 ;
  assign n10822 = ( x118 & n10820 ) | ( x118 & ~n10821 ) | ( n10820 & ~n10821 ) ;
  assign n10823 = n3346 & n9733 ;
  assign n10824 = n10822 | n10823 ;
  assign n10825 = n10824 ^ x29 ^ 1'b0 ;
  assign n10826 = ( n9430 & n10816 ) | ( n9430 & n10825 ) | ( n10816 & n10825 ) ;
  assign n10827 = n10825 ^ n10816 ^ n9430 ;
  assign n10828 = x120 & n3734 ;
  assign n10829 = ( x122 & n3732 ) | ( x122 & n10828 ) | ( n3732 & n10828 ) ;
  assign n10830 = n10828 | n10829 ;
  assign n10831 = x121 & ~n3737 ;
  assign n10832 = ( x121 & n10830 ) | ( x121 & ~n10831 ) | ( n10830 & ~n10831 ) ;
  assign n10833 = n3736 & n9806 ;
  assign n10834 = n10832 | n10833 ;
  assign n10835 = n10834 ^ x26 ^ 1'b0 ;
  assign n10836 = ( n10694 & n10827 ) | ( n10694 & n10835 ) | ( n10827 & n10835 ) ;
  assign n10837 = n10835 ^ n10827 ^ n10694 ;
  assign n10838 = x123 & n4616 ;
  assign n10839 = ( x125 & n4606 ) | ( x125 & n10838 ) | ( n4606 & n10838 ) ;
  assign n10840 = n10838 | n10839 ;
  assign n10841 = x124 & ~n4605 ;
  assign n10842 = ( x124 & n10840 ) | ( x124 & ~n10841 ) | ( n10840 & ~n10841 ) ;
  assign n10843 = n4608 & n9883 ;
  assign n10844 = n10842 | n10843 ;
  assign n10845 = n10844 ^ x23 ^ 1'b0 ;
  assign n10846 = ( n10699 & n10837 ) | ( n10699 & n10845 ) | ( n10837 & n10845 ) ;
  assign n10847 = n10845 ^ n10837 ^ n10699 ;
  assign n10848 = n10847 ^ n10701 ^ n10682 ;
  assign n10849 = n10848 ^ n10704 ^ n10703 ;
  assign n10850 = ( n10703 & n10704 ) | ( n10703 & n10848 ) | ( n10704 & n10848 ) ;
  assign n10851 = x125 & n4616 ;
  assign n10852 = ( x127 & n4606 ) | ( x127 & n10851 ) | ( n4606 & n10851 ) ;
  assign n10853 = n10851 | n10852 ;
  assign n10854 = x124 & n4616 ;
  assign n10855 = ( n10682 & n10701 ) | ( n10682 & n10847 ) | ( n10701 & n10847 ) ;
  assign n10856 = x127 & ~n4605 ;
  assign n10857 = ( x126 & n4606 ) | ( x126 & n10854 ) | ( n4606 & n10854 ) ;
  assign n10858 = x127 & n4616 ;
  assign n10859 = x126 & n4616 ;
  assign n10860 = ( x127 & ~n10856 ) | ( x127 & n10859 ) | ( ~n10856 & n10859 ) ;
  assign n10861 = ( n4608 & n9958 ) | ( n4608 & n10859 ) | ( n9958 & n10859 ) ;
  assign n10862 = n10860 | n10861 ;
  assign n10863 = ( n4608 & n9968 ) | ( n4608 & n10858 ) | ( n9968 & n10858 ) ;
  assign n10864 = n10858 | n10863 ;
  assign n10865 = x126 & ~n4605 ;
  assign n10866 = x125 & ~n4605 ;
  assign n10867 = n10854 | n10857 ;
  assign n10868 = ( x125 & ~n10866 ) | ( x125 & n10867 ) | ( ~n10866 & n10867 ) ;
  assign n10869 = n4608 & n9917 ;
  assign n10870 = x91 & n263 ;
  assign n10871 = n10868 | n10869 ;
  assign n10872 = n4608 & n9949 ;
  assign n10873 = ( x93 & n264 ) | ( x93 & n10870 ) | ( n264 & n10870 ) ;
  assign n10874 = n10870 | n10873 ;
  assign n10875 = ( x126 & n10853 ) | ( x126 & ~n10865 ) | ( n10853 & ~n10865 ) ;
  assign n10876 = n10872 | n10875 ;
  assign n10877 = n10871 ^ x23 ^ 1'b0 ;
  assign n10878 = x88 & n133 ;
  assign n10879 = ( x90 & n142 ) | ( x90 & n10878 ) | ( n142 & n10878 ) ;
  assign n10880 = x89 & ~n134 ;
  assign n10881 = n10878 | n10879 ;
  assign n10882 = ( x89 & ~n10880 ) | ( x89 & n10881 ) | ( ~n10880 & n10881 ) ;
  assign n10883 = n140 & n1741 ;
  assign n10884 = n10882 | n10883 ;
  assign n10885 = x84 & ~n242 ;
  assign n10886 = x83 & n325 ;
  assign n10887 = ( x84 & ~n10885 ) | ( x84 & n10886 ) | ( ~n10885 & n10886 ) ;
  assign n10888 = ( n10712 & n10771 ) | ( n10712 & ~n10887 ) | ( n10771 & ~n10887 ) ;
  assign n10889 = n10887 ^ n10771 ^ n10712 ;
  assign n10890 = n10884 ^ x59 ^ 1'b0 ;
  assign n10891 = ( n10716 & ~n10889 ) | ( n10716 & n10890 ) | ( ~n10889 & n10890 ) ;
  assign n10892 = n10890 ^ n10889 ^ n10716 ;
  assign n10893 = n272 & n2476 ;
  assign n10894 = x92 & ~n260 ;
  assign n10895 = ( x92 & n10874 ) | ( x92 & ~n10894 ) | ( n10874 & ~n10894 ) ;
  assign n10896 = n10893 | n10895 ;
  assign n10897 = n10896 ^ x56 ^ 1'b0 ;
  assign n10898 = n10897 ^ n10892 ^ n10719 ;
  assign n10899 = x97 & n561 ;
  assign n10900 = ( n10719 & ~n10892 ) | ( n10719 & n10897 ) | ( ~n10892 & n10897 ) ;
  assign n10901 = ( x99 & n551 ) | ( x99 & n10899 ) | ( n551 & n10899 ) ;
  assign n10902 = x94 & n408 ;
  assign n10903 = n10899 | n10901 ;
  assign n10904 = x98 & ~n550 ;
  assign n10905 = ( x98 & n10903 ) | ( x98 & ~n10904 ) | ( n10903 & ~n10904 ) ;
  assign n10906 = ( x96 & n403 ) | ( x96 & n10902 ) | ( n403 & n10902 ) ;
  assign n10907 = n10902 | n10906 ;
  assign n10908 = n553 & n4270 ;
  assign n10909 = n10905 | n10908 ;
  assign n10910 = x95 & ~n410 ;
  assign n10911 = n10909 ^ x50 ^ 1'b0 ;
  assign n10912 = ( x95 & n10907 ) | ( x95 & ~n10910 ) | ( n10907 & ~n10910 ) ;
  assign n10913 = n402 & n2907 ;
  assign n10914 = n10912 | n10913 ;
  assign n10915 = n10914 ^ x53 ^ 1'b0 ;
  assign n10916 = ( n10729 & ~n10898 ) | ( n10729 & n10915 ) | ( ~n10898 & n10915 ) ;
  assign n10917 = n10915 ^ n10898 ^ n10729 ;
  assign n10918 = x106 & n1058 ;
  assign n10919 = ( x108 & n1065 ) | ( x108 & n10918 ) | ( n1065 & n10918 ) ;
  assign n10920 = n10918 | n10919 ;
  assign n10921 = n10917 ^ n10911 ^ n10738 ;
  assign n10922 = ( n10738 & n10911 ) | ( n10738 & ~n10917 ) | ( n10911 & ~n10917 ) ;
  assign n10923 = x107 & ~n1060 ;
  assign n10924 = ( x107 & n10920 ) | ( x107 & ~n10923 ) | ( n10920 & ~n10923 ) ;
  assign n10925 = x100 & n744 ;
  assign n10926 = n1063 & n8557 ;
  assign n10927 = n10924 | n10926 ;
  assign n10928 = n10927 ^ x41 ^ 1'b0 ;
  assign n10929 = ( x102 & n730 ) | ( x102 & n10925 ) | ( n730 & n10925 ) ;
  assign n10930 = n10925 | n10929 ;
  assign n10931 = x101 & ~n732 ;
  assign n10932 = ( x101 & n10930 ) | ( x101 & ~n10931 ) | ( n10930 & ~n10931 ) ;
  assign n10933 = n731 & n5947 ;
  assign n10934 = n10932 | n10933 ;
  assign n10935 = n10934 ^ x47 ^ 1'b0 ;
  assign n10936 = n10935 ^ n10921 ^ n10748 ;
  assign n10937 = ( n10748 & ~n10921 ) | ( n10748 & n10935 ) | ( ~n10921 & n10935 ) ;
  assign n10938 = x103 & n888 ;
  assign n10939 = ( x105 & n878 ) | ( x105 & n10938 ) | ( n878 & n10938 ) ;
  assign n10940 = n10938 | n10939 ;
  assign n10941 = x104 & ~n877 ;
  assign n10942 = ( x104 & n10940 ) | ( x104 & ~n10941 ) | ( n10940 & ~n10941 ) ;
  assign n10943 = n880 & n8105 ;
  assign n10944 = n10942 | n10943 ;
  assign n10945 = n10944 ^ x44 ^ 1'b0 ;
  assign n10946 = n10945 ^ n10936 ^ n10759 ;
  assign n10947 = ( n10759 & ~n10936 ) | ( n10759 & n10945 ) | ( ~n10936 & n10945 ) ;
  assign n10948 = ( n10776 & n10928 ) | ( n10776 & ~n10946 ) | ( n10928 & ~n10946 ) ;
  assign n10949 = n10946 ^ n10928 ^ n10776 ;
  assign n10950 = x109 & n2156 ;
  assign n10951 = ( x111 & n2163 ) | ( x111 & n10950 ) | ( n2163 & n10950 ) ;
  assign n10952 = n10950 | n10951 ;
  assign n10953 = x110 & ~n2158 ;
  assign n10954 = ( x110 & n10952 ) | ( x110 & ~n10953 ) | ( n10952 & ~n10953 ) ;
  assign n10955 = n2161 & n8946 ;
  assign n10956 = n10954 | n10955 ;
  assign n10957 = n10956 ^ x38 ^ 1'b0 ;
  assign n10958 = ( n10787 & n10949 ) | ( n10787 & ~n10957 ) | ( n10949 & ~n10957 ) ;
  assign n10959 = n10957 ^ n10949 ^ n10787 ;
  assign n10960 = x112 & n2560 ;
  assign n10961 = ( x114 & n2567 ) | ( x114 & n10960 ) | ( n2567 & n10960 ) ;
  assign n10962 = n10960 | n10961 ;
  assign n10963 = x113 & ~n2562 ;
  assign n10964 = ( x113 & n10962 ) | ( x113 & ~n10963 ) | ( n10962 & ~n10963 ) ;
  assign n10965 = n2565 & n9279 ;
  assign n10966 = n10964 | n10965 ;
  assign n10967 = n10966 ^ x35 ^ 1'b0 ;
  assign n10968 = ( n10797 & n10959 ) | ( n10797 & n10967 ) | ( n10959 & n10967 ) ;
  assign n10969 = n10967 ^ n10959 ^ n10797 ;
  assign n10970 = x115 & n3025 ;
  assign n10971 = ( x117 & n3015 ) | ( x117 & n10970 ) | ( n3015 & n10970 ) ;
  assign n10972 = n10970 | n10971 ;
  assign n10973 = x116 & ~n3014 ;
  assign n10974 = ( x116 & n10972 ) | ( x116 & ~n10973 ) | ( n10972 & ~n10973 ) ;
  assign n10975 = n3017 & n9569 ;
  assign n10976 = n10673 ^ x20 ^ 1'b0 ;
  assign n10977 = n10974 | n10975 ;
  assign n10978 = n10977 ^ x32 ^ 1'b0 ;
  assign n10979 = ( n10807 & n10969 ) | ( n10807 & n10978 ) | ( n10969 & n10978 ) ;
  assign n10980 = n10978 ^ n10969 ^ n10807 ;
  assign n10981 = x118 & n3344 ;
  assign n10982 = ( x120 & n3342 ) | ( x120 & n10981 ) | ( n3342 & n10981 ) ;
  assign n10983 = n10981 | n10982 ;
  assign n10984 = x119 & ~n3347 ;
  assign n10985 = ( x119 & n10983 ) | ( x119 & ~n10984 ) | ( n10983 & ~n10984 ) ;
  assign n10986 = n3346 & n9756 ;
  assign n10987 = n10985 | n10986 ;
  assign n10988 = n10987 ^ x29 ^ 1'b0 ;
  assign n10989 = ( n10817 & n10980 ) | ( n10817 & n10988 ) | ( n10980 & n10988 ) ;
  assign n10990 = n10988 ^ n10980 ^ n10817 ;
  assign n10991 = x121 & n3734 ;
  assign n10992 = ( x123 & n3732 ) | ( x123 & n10991 ) | ( n3732 & n10991 ) ;
  assign n10993 = n10991 | n10992 ;
  assign n10994 = x122 & ~n3737 ;
  assign n10995 = ( x122 & n10993 ) | ( x122 & ~n10994 ) | ( n10993 & ~n10994 ) ;
  assign n10996 = n3736 & n9828 ;
  assign n10997 = n10995 | n10996 ;
  assign n10998 = n10997 ^ x26 ^ 1'b0 ;
  assign n10999 = ( n10826 & n10990 ) | ( n10826 & n10998 ) | ( n10990 & n10998 ) ;
  assign n11000 = n10998 ^ n10990 ^ n10826 ;
  assign n11001 = n11000 ^ n10877 ^ n10836 ;
  assign n11002 = ( n10836 & n10877 ) | ( n10836 & n11000 ) | ( n10877 & n11000 ) ;
  assign n11003 = ( n10846 & n10976 ) | ( n10846 & n11001 ) | ( n10976 & n11001 ) ;
  assign n11004 = n11001 ^ n10976 ^ n10846 ;
  assign n11005 = n11004 ^ n10855 ^ n10850 ;
  assign n11006 = ( n10850 & n10855 ) | ( n10850 & n11004 ) | ( n10855 & n11004 ) ;
  assign n11007 = x86 & n208 ;
  assign n11008 = n197 & n1569 ;
  assign n11009 = ( x88 & n194 ) | ( x88 & n11007 ) | ( n194 & n11007 ) ;
  assign n11010 = n11007 | n11009 ;
  assign n11011 = x87 & ~n192 ;
  assign n11012 = ( x87 & n11010 ) | ( x87 & ~n11011 ) | ( n11010 & ~n11011 ) ;
  assign n11013 = x85 & ~n242 ;
  assign n11014 = n11008 | n11012 ;
  assign n11015 = n11014 ^ x62 ^ 1'b0 ;
  assign n11016 = x84 & n325 ;
  assign n11017 = ( x85 & ~n11013 ) | ( x85 & n11016 ) | ( ~n11013 & n11016 ) ;
  assign n11018 = ( ~x20 & n10887 ) | ( ~x20 & n11017 ) | ( n10887 & n11017 ) ;
  assign n11019 = n11017 ^ n10887 ^ x20 ;
  assign n11020 = ( n10888 & n11015 ) | ( n10888 & ~n11019 ) | ( n11015 & ~n11019 ) ;
  assign n11021 = n11019 ^ n11015 ^ n10888 ;
  assign n11022 = x89 & n133 ;
  assign n11023 = ( x91 & n142 ) | ( x91 & n11022 ) | ( n142 & n11022 ) ;
  assign n11024 = n11022 | n11023 ;
  assign n11025 = x90 & ~n134 ;
  assign n11026 = ( x90 & n11024 ) | ( x90 & ~n11025 ) | ( n11024 & ~n11025 ) ;
  assign n11027 = n140 & n2114 ;
  assign n11028 = n11026 | n11027 ;
  assign n11029 = n11028 ^ x59 ^ 1'b0 ;
  assign n11030 = ( n10891 & ~n11021 ) | ( n10891 & n11029 ) | ( ~n11021 & n11029 ) ;
  assign n11031 = n11029 ^ n11021 ^ n10891 ;
  assign n11032 = x92 & n263 ;
  assign n11033 = ( x94 & n264 ) | ( x94 & n11032 ) | ( n264 & n11032 ) ;
  assign n11034 = n11032 | n11033 ;
  assign n11035 = x93 & ~n260 ;
  assign n11036 = ( x93 & n11034 ) | ( x93 & ~n11035 ) | ( n11034 & ~n11035 ) ;
  assign n11037 = n197 & n2114 ;
  assign n11038 = n272 & n2518 ;
  assign n11039 = n11036 | n11038 ;
  assign n11040 = n11039 ^ x56 ^ 1'b0 ;
  assign n11041 = ( n10900 & ~n11031 ) | ( n10900 & n11040 ) | ( ~n11031 & n11040 ) ;
  assign n11042 = n11040 ^ n11031 ^ n10900 ;
  assign n11043 = x95 & n408 ;
  assign n11044 = ( x97 & n403 ) | ( x97 & n11043 ) | ( n403 & n11043 ) ;
  assign n11045 = n11043 | n11044 ;
  assign n11046 = x96 & ~n410 ;
  assign n11047 = ( x96 & n11045 ) | ( x96 & ~n11046 ) | ( n11045 & ~n11046 ) ;
  assign n11048 = n402 & n3668 ;
  assign n11049 = n11047 | n11048 ;
  assign n11050 = n11049 ^ x53 ^ 1'b0 ;
  assign n11051 = ( n10916 & ~n11042 ) | ( n10916 & n11050 ) | ( ~n11042 & n11050 ) ;
  assign n11052 = n11050 ^ n11042 ^ n10916 ;
  assign n11053 = x98 & n561 ;
  assign n11054 = ( x100 & n551 ) | ( x100 & n11053 ) | ( n551 & n11053 ) ;
  assign n11055 = n11053 | n11054 ;
  assign n11056 = x99 & ~n550 ;
  assign n11057 = ( x99 & n11055 ) | ( x99 & ~n11056 ) | ( n11055 & ~n11056 ) ;
  assign n11058 = n553 & n4334 ;
  assign n11059 = n11057 | n11058 ;
  assign n11060 = n11059 ^ x50 ^ 1'b0 ;
  assign n11061 = ( n10922 & ~n11052 ) | ( n10922 & n11060 ) | ( ~n11052 & n11060 ) ;
  assign n11062 = n11060 ^ n11052 ^ n10922 ;
  assign n11063 = x89 & n208 ;
  assign n11064 = ( x91 & n194 ) | ( x91 & n11063 ) | ( n194 & n11063 ) ;
  assign n11065 = n11063 | n11064 ;
  assign n11066 = x90 & ~n192 ;
  assign n11067 = ( x90 & n11065 ) | ( x90 & ~n11066 ) | ( n11065 & ~n11066 ) ;
  assign n11068 = x101 & n744 ;
  assign n11069 = n11037 | n11067 ;
  assign n11070 = ( x103 & n730 ) | ( x103 & n11068 ) | ( n730 & n11068 ) ;
  assign n11071 = n11068 | n11070 ;
  assign n11072 = x102 & ~n732 ;
  assign n11073 = ( x102 & n11071 ) | ( x102 & ~n11072 ) | ( n11071 & ~n11072 ) ;
  assign n11074 = n731 & n7860 ;
  assign n11075 = n11073 | n11074 ;
  assign n11076 = n11075 ^ x47 ^ 1'b0 ;
  assign n11077 = ( n10937 & ~n11062 ) | ( n10937 & n11076 ) | ( ~n11062 & n11076 ) ;
  assign n11078 = n11076 ^ n11062 ^ n10937 ;
  assign n11079 = x104 & n888 ;
  assign n11080 = ( x106 & n878 ) | ( x106 & n11079 ) | ( n878 & n11079 ) ;
  assign n11081 = n11079 | n11080 ;
  assign n11082 = x105 & ~n877 ;
  assign n11083 = ( x105 & n11081 ) | ( x105 & ~n11082 ) | ( n11081 & ~n11082 ) ;
  assign n11084 = n880 & n8287 ;
  assign n11085 = n11083 | n11084 ;
  assign n11086 = n11085 ^ x44 ^ 1'b0 ;
  assign n11087 = n11086 ^ n11078 ^ n10947 ;
  assign n11088 = ( n10947 & ~n11078 ) | ( n10947 & n11086 ) | ( ~n11078 & n11086 ) ;
  assign n11089 = x107 & n1058 ;
  assign n11090 = ( x109 & n1065 ) | ( x109 & n11089 ) | ( n1065 & n11089 ) ;
  assign n11091 = n11089 | n11090 ;
  assign n11092 = x108 & ~n1060 ;
  assign n11093 = ( x108 & n11091 ) | ( x108 & ~n11092 ) | ( n11091 & ~n11092 ) ;
  assign n11094 = n1063 & n8680 ;
  assign n11095 = n11093 | n11094 ;
  assign n11096 = n11095 ^ x41 ^ 1'b0 ;
  assign n11097 = n11096 ^ n11087 ^ n10948 ;
  assign n11098 = ( n10948 & ~n11087 ) | ( n10948 & n11096 ) | ( ~n11087 & n11096 ) ;
  assign n11099 = x110 & n2156 ;
  assign n11100 = ( x112 & n2163 ) | ( x112 & n11099 ) | ( n2163 & n11099 ) ;
  assign n11101 = n11099 | n11100 ;
  assign n11102 = x111 & ~n2158 ;
  assign n11103 = n10876 ^ x23 ^ 1'b0 ;
  assign n11104 = n11069 ^ x62 ^ 1'b0 ;
  assign n11105 = n10864 ^ x23 ^ 1'b0 ;
  assign n11106 = ( x111 & n11101 ) | ( x111 & ~n11102 ) | ( n11101 & ~n11102 ) ;
  assign n11107 = n2161 & n9080 ;
  assign n11108 = n11106 | n11107 ;
  assign n11109 = n11108 ^ x38 ^ 1'b0 ;
  assign n11110 = ( n10958 & n11097 ) | ( n10958 & ~n11109 ) | ( n11097 & ~n11109 ) ;
  assign n11111 = n11109 ^ n11097 ^ n10958 ;
  assign n11112 = x113 & n2560 ;
  assign n11113 = ( x115 & n2567 ) | ( x115 & n11112 ) | ( n2567 & n11112 ) ;
  assign n11114 = n11112 | n11113 ;
  assign n11115 = x114 & ~n2562 ;
  assign n11116 = ( x114 & n11114 ) | ( x114 & ~n11115 ) | ( n11114 & ~n11115 ) ;
  assign n11117 = n2565 & n9414 ;
  assign n11118 = n11116 | n11117 ;
  assign n11119 = n11118 ^ x35 ^ 1'b0 ;
  assign n11120 = ( n10968 & n11111 ) | ( n10968 & n11119 ) | ( n11111 & n11119 ) ;
  assign n11121 = n11119 ^ n11111 ^ n10968 ;
  assign n11122 = x116 & n3025 ;
  assign n11123 = ( x118 & n3015 ) | ( x118 & n11122 ) | ( n3015 & n11122 ) ;
  assign n11124 = n11122 | n11123 ;
  assign n11125 = x117 & ~n3014 ;
  assign n11126 = ( x117 & n11124 ) | ( x117 & ~n11125 ) | ( n11124 & ~n11125 ) ;
  assign n11127 = n3017 & n9671 ;
  assign n11128 = n11126 | n11127 ;
  assign n11129 = n11128 ^ x32 ^ 1'b0 ;
  assign n11130 = n11129 ^ n11121 ^ n10979 ;
  assign n11131 = ( n10979 & n11121 ) | ( n10979 & n11129 ) | ( n11121 & n11129 ) ;
  assign n11132 = x119 & n3344 ;
  assign n11133 = ( x121 & n3342 ) | ( x121 & n11132 ) | ( n3342 & n11132 ) ;
  assign n11134 = n11132 | n11133 ;
  assign n11135 = x120 & ~n3347 ;
  assign n11136 = ( x120 & n11134 ) | ( x120 & ~n11135 ) | ( n11134 & ~n11135 ) ;
  assign n11137 = n3346 & n9808 ;
  assign n11138 = n11136 | n11137 ;
  assign n11139 = n11138 ^ x29 ^ 1'b0 ;
  assign n11140 = ( n10989 & n11130 ) | ( n10989 & n11139 ) | ( n11130 & n11139 ) ;
  assign n11141 = n11139 ^ n11130 ^ n10989 ;
  assign n11142 = x122 & n3734 ;
  assign n11143 = ( x124 & n3732 ) | ( x124 & n11142 ) | ( n3732 & n11142 ) ;
  assign n11144 = n11142 | n11143 ;
  assign n11145 = x123 & ~n3737 ;
  assign n11146 = ( x123 & n11144 ) | ( x123 & ~n11145 ) | ( n11144 & ~n11145 ) ;
  assign n11147 = n3736 & n9858 ;
  assign n11148 = n11146 | n11147 ;
  assign n11149 = n11148 ^ x26 ^ 1'b0 ;
  assign n11150 = ( n10999 & n11141 ) | ( n10999 & n11149 ) | ( n11141 & n11149 ) ;
  assign n11151 = n11149 ^ n11141 ^ n10999 ;
  assign n11152 = x87 & n208 ;
  assign n11153 = ( x89 & n194 ) | ( x89 & n11152 ) | ( n194 & n11152 ) ;
  assign n11154 = n11152 | n11153 ;
  assign n11155 = x88 & ~n192 ;
  assign n11156 = ( x88 & n11154 ) | ( x88 & ~n11155 ) | ( n11154 & ~n11155 ) ;
  assign n11157 = ( n11002 & n11103 ) | ( n11002 & n11151 ) | ( n11103 & n11151 ) ;
  assign n11158 = n11151 ^ n11103 ^ n11002 ;
  assign n11159 = ( n197 & n1654 ) | ( n197 & n11156 ) | ( n1654 & n11156 ) ;
  assign n11160 = x88 & n208 ;
  assign n11161 = ( x90 & n194 ) | ( x90 & n11160 ) | ( n194 & n11160 ) ;
  assign n11162 = n11160 | n11161 ;
  assign n11163 = x89 & ~n192 ;
  assign n11164 = n11156 | n11159 ;
  assign n11165 = ( x89 & n11162 ) | ( x89 & ~n11163 ) | ( n11162 & ~n11163 ) ;
  assign n11166 = ( n197 & n1741 ) | ( n197 & n11165 ) | ( n1741 & n11165 ) ;
  assign n11167 = n11165 | n11166 ;
  assign n11168 = n11164 ^ x62 ^ 1'b0 ;
  assign n11169 = n11158 ^ n11006 ^ n11003 ;
  assign n11170 = ( n11003 & n11006 ) | ( n11003 & n11158 ) | ( n11006 & n11158 ) ;
  assign n11171 = x90 & n133 ;
  assign n11172 = x91 & ~n134 ;
  assign n11173 = ( x92 & n142 ) | ( x92 & n11171 ) | ( n142 & n11171 ) ;
  assign n11174 = n11171 | n11173 ;
  assign n11175 = ( x91 & ~n11172 ) | ( x91 & n11174 ) | ( ~n11172 & n11174 ) ;
  assign n11176 = n140 & n2420 ;
  assign n11177 = n11175 | n11176 ;
  assign n11178 = x85 & n325 ;
  assign n11179 = x86 & ~n242 ;
  assign n11180 = ( x86 & n11178 ) | ( x86 & ~n11179 ) | ( n11178 & ~n11179 ) ;
  assign n11181 = n11180 ^ n11168 ^ n11018 ;
  assign n11182 = ( n11018 & n11168 ) | ( n11018 & ~n11180 ) | ( n11168 & ~n11180 ) ;
  assign n11183 = n11177 ^ x59 ^ 1'b0 ;
  assign n11184 = ( n11020 & ~n11181 ) | ( n11020 & n11183 ) | ( ~n11181 & n11183 ) ;
  assign n11185 = n11183 ^ n11181 ^ n11020 ;
  assign n11186 = x93 & n263 ;
  assign n11187 = ( x95 & n264 ) | ( x95 & n11186 ) | ( n264 & n11186 ) ;
  assign n11188 = n11186 | n11187 ;
  assign n11189 = x94 & ~n260 ;
  assign n11190 = ( x94 & n11188 ) | ( x94 & ~n11189 ) | ( n11188 & ~n11189 ) ;
  assign n11191 = n272 & n2854 ;
  assign n11192 = n11190 | n11191 ;
  assign n11193 = n11192 ^ x56 ^ 1'b0 ;
  assign n11194 = n11193 ^ n11185 ^ n11030 ;
  assign n11195 = ( n11030 & ~n11185 ) | ( n11030 & n11193 ) | ( ~n11185 & n11193 ) ;
  assign n11196 = x96 & n408 ;
  assign n11197 = ( x98 & n403 ) | ( x98 & n11196 ) | ( n403 & n11196 ) ;
  assign n11198 = n11196 | n11197 ;
  assign n11199 = x97 & ~n410 ;
  assign n11200 = ( x97 & n11198 ) | ( x97 & ~n11199 ) | ( n11198 & ~n11199 ) ;
  assign n11201 = n402 & n4052 ;
  assign n11202 = n11200 | n11201 ;
  assign n11203 = n11202 ^ x53 ^ 1'b0 ;
  assign n11204 = ( n11041 & ~n11194 ) | ( n11041 & n11203 ) | ( ~n11194 & n11203 ) ;
  assign n11205 = n11203 ^ n11194 ^ n11041 ;
  assign n11206 = x99 & n561 ;
  assign n11207 = ( x101 & n551 ) | ( x101 & n11206 ) | ( n551 & n11206 ) ;
  assign n11208 = n11206 | n11207 ;
  assign n11209 = x100 & ~n550 ;
  assign n11210 = ( x100 & n11208 ) | ( x100 & ~n11209 ) | ( n11208 & ~n11209 ) ;
  assign n11211 = n553 & n5687 ;
  assign n11212 = n11210 | n11211 ;
  assign n11213 = n11212 ^ x50 ^ 1'b0 ;
  assign n11214 = n11213 ^ n11205 ^ n11051 ;
  assign n11215 = ( n11051 & ~n11205 ) | ( n11051 & n11213 ) | ( ~n11205 & n11213 ) ;
  assign n11216 = x102 & n744 ;
  assign n11217 = ( x104 & n730 ) | ( x104 & n11216 ) | ( n730 & n11216 ) ;
  assign n11218 = n11216 | n11217 ;
  assign n11219 = x103 & ~n732 ;
  assign n11220 = ( x103 & n11218 ) | ( x103 & ~n11219 ) | ( n11218 & ~n11219 ) ;
  assign n11221 = n731 & n8012 ;
  assign n11222 = n11220 | n11221 ;
  assign n11223 = n11222 ^ x47 ^ 1'b0 ;
  assign n11224 = n11223 ^ n11214 ^ n11061 ;
  assign n11225 = ( n11061 & ~n11214 ) | ( n11061 & n11223 ) | ( ~n11214 & n11223 ) ;
  assign n11226 = x105 & n888 ;
  assign n11227 = ( x107 & n878 ) | ( x107 & n11226 ) | ( n878 & n11226 ) ;
  assign n11228 = n11226 | n11227 ;
  assign n11229 = x106 & ~n877 ;
  assign n11230 = ( x106 & n11228 ) | ( x106 & ~n11229 ) | ( n11228 & ~n11229 ) ;
  assign n11231 = n880 & n8440 ;
  assign n11232 = n11230 | n11231 ;
  assign n11233 = n11232 ^ x44 ^ 1'b0 ;
  assign n11234 = ( n11077 & ~n11224 ) | ( n11077 & n11233 ) | ( ~n11224 & n11233 ) ;
  assign n11235 = n11233 ^ n11224 ^ n11077 ;
  assign n11236 = x108 & n1058 ;
  assign n11237 = ( x110 & n1065 ) | ( x110 & n11236 ) | ( n1065 & n11236 ) ;
  assign n11238 = n11236 | n11237 ;
  assign n11239 = x109 & ~n1060 ;
  assign n11240 = ( x109 & n11238 ) | ( x109 & ~n11239 ) | ( n11238 & ~n11239 ) ;
  assign n11241 = n1063 & n8820 ;
  assign n11242 = n11240 | n11241 ;
  assign n11243 = n11242 ^ x41 ^ 1'b0 ;
  assign n11244 = ( n11088 & ~n11235 ) | ( n11088 & n11243 ) | ( ~n11235 & n11243 ) ;
  assign n11245 = n11243 ^ n11235 ^ n11088 ;
  assign n11246 = x111 & n2156 ;
  assign n11247 = ( x113 & n2163 ) | ( x113 & n11246 ) | ( n2163 & n11246 ) ;
  assign n11248 = n11246 | n11247 ;
  assign n11249 = x112 & ~n2158 ;
  assign n11250 = ( x112 & n11248 ) | ( x112 & ~n11249 ) | ( n11248 & ~n11249 ) ;
  assign n11251 = n2161 & n9199 ;
  assign n11252 = n11250 | n11251 ;
  assign n11253 = n11252 ^ x38 ^ 1'b0 ;
  assign n11254 = ( n11098 & ~n11245 ) | ( n11098 & n11253 ) | ( ~n11245 & n11253 ) ;
  assign n11255 = n11253 ^ n11245 ^ n11098 ;
  assign n11256 = x114 & n2560 ;
  assign n11257 = ( x116 & n2567 ) | ( x116 & n11256 ) | ( n2567 & n11256 ) ;
  assign n11258 = n11256 | n11257 ;
  assign n11259 = x115 & ~n2562 ;
  assign n11260 = ( x115 & n11258 ) | ( x115 & ~n11259 ) | ( n11258 & ~n11259 ) ;
  assign n11261 = n2565 & n9513 ;
  assign n11262 = n11260 | n11261 ;
  assign n11263 = n11262 ^ x35 ^ 1'b0 ;
  assign n11264 = n11263 ^ n11255 ^ n11110 ;
  assign n11265 = ( n11110 & n11255 ) | ( n11110 & ~n11263 ) | ( n11255 & ~n11263 ) ;
  assign n11266 = x117 & n3025 ;
  assign n11267 = ( x119 & n3015 ) | ( x119 & n11266 ) | ( n3015 & n11266 ) ;
  assign n11268 = n11266 | n11267 ;
  assign n11269 = x118 & ~n3014 ;
  assign n11270 = ( x118 & n11268 ) | ( x118 & ~n11269 ) | ( n11268 & ~n11269 ) ;
  assign n11271 = n3017 & n9733 ;
  assign n11272 = n11270 | n11271 ;
  assign n11273 = n11272 ^ x32 ^ 1'b0 ;
  assign n11274 = n11273 ^ n11264 ^ n11120 ;
  assign n11275 = ( n11120 & n11264 ) | ( n11120 & n11273 ) | ( n11264 & n11273 ) ;
  assign n11276 = x120 & n3344 ;
  assign n11277 = ( x122 & n3342 ) | ( x122 & n11276 ) | ( n3342 & n11276 ) ;
  assign n11278 = n11276 | n11277 ;
  assign n11279 = x121 & ~n3347 ;
  assign n11280 = ( x121 & n11278 ) | ( x121 & ~n11279 ) | ( n11278 & ~n11279 ) ;
  assign n11281 = ( n3346 & n9806 ) | ( n3346 & n11280 ) | ( n9806 & n11280 ) ;
  assign n11282 = n11280 | n11281 ;
  assign n11283 = n11282 ^ x29 ^ 1'b0 ;
  assign n11284 = n11283 ^ n11274 ^ n11131 ;
  assign n11285 = ( n11131 & n11274 ) | ( n11131 & n11283 ) | ( n11274 & n11283 ) ;
  assign n11286 = x123 & n3734 ;
  assign n11287 = ( x125 & n3732 ) | ( x125 & n11286 ) | ( n3732 & n11286 ) ;
  assign n11288 = n11286 | n11287 ;
  assign n11289 = x124 & ~n3737 ;
  assign n11290 = n10862 ^ x23 ^ 1'b0 ;
  assign n11291 = ( x124 & n11288 ) | ( x124 & ~n11289 ) | ( n11288 & ~n11289 ) ;
  assign n11292 = n3736 & n9883 ;
  assign n11293 = n11291 | n11292 ;
  assign n11294 = n11293 ^ x26 ^ 1'b0 ;
  assign n11295 = n11294 ^ n11284 ^ n11140 ;
  assign n11296 = ( n11140 & n11284 ) | ( n11140 & n11294 ) | ( n11284 & n11294 ) ;
  assign n11297 = n11295 ^ n11290 ^ n11150 ;
  assign n11298 = ( n11150 & n11290 ) | ( n11150 & n11295 ) | ( n11290 & n11295 ) ;
  assign n11299 = x126 & n3734 ;
  assign n11300 = x127 & ~n3737 ;
  assign n11301 = n11297 ^ n11170 ^ n11157 ;
  assign n11302 = ( n11157 & n11170 ) | ( n11157 & n11297 ) | ( n11170 & n11297 ) ;
  assign n11303 = ( x127 & n11299 ) | ( x127 & ~n11300 ) | ( n11299 & ~n11300 ) ;
  assign n11304 = ( n3736 & n9958 ) | ( n3736 & n11299 ) | ( n9958 & n11299 ) ;
  assign n11305 = x124 & n3734 ;
  assign n11306 = ( x126 & n3732 ) | ( x126 & n11305 ) | ( n3732 & n11305 ) ;
  assign n11307 = n11305 | n11306 ;
  assign n11308 = x125 & ~n3737 ;
  assign n11309 = n11303 | n11304 ;
  assign n11310 = x127 & n3734 ;
  assign n11311 = ( x125 & n11307 ) | ( x125 & ~n11308 ) | ( n11307 & ~n11308 ) ;
  assign n11312 = ( n3736 & n9968 ) | ( n3736 & n11310 ) | ( n9968 & n11310 ) ;
  assign n11313 = n11310 | n11312 ;
  assign n11314 = n3736 & n9917 ;
  assign n11315 = x125 & n3734 ;
  assign n11316 = ( x127 & n3732 ) | ( x127 & n11315 ) | ( n3732 & n11315 ) ;
  assign n11317 = n3736 & n9949 ;
  assign n11318 = x126 & ~n3737 ;
  assign n11319 = n11315 | n11316 ;
  assign n11320 = n11311 | n11314 ;
  assign n11321 = ( x126 & ~n11318 ) | ( x126 & n11319 ) | ( ~n11318 & n11319 ) ;
  assign n11322 = n11317 | n11321 ;
  assign n11323 = n11320 ^ x26 ^ 1'b0 ;
  assign n11324 = n11167 ^ x62 ^ 1'b0 ;
  assign n11325 = x91 & n133 ;
  assign n11326 = x92 & ~n134 ;
  assign n11327 = ( x93 & n142 ) | ( x93 & n11325 ) | ( n142 & n11325 ) ;
  assign n11328 = n11325 | n11327 ;
  assign n11329 = x86 & n325 ;
  assign n11330 = ( x92 & ~n11326 ) | ( x92 & n11328 ) | ( ~n11326 & n11328 ) ;
  assign n11331 = x87 & ~n242 ;
  assign n11332 = ( x87 & n11329 ) | ( x87 & ~n11331 ) | ( n11329 & ~n11331 ) ;
  assign n11333 = n140 & n2476 ;
  assign n11334 = n11330 | n11333 ;
  assign n11335 = ( n11180 & n11324 ) | ( n11180 & ~n11332 ) | ( n11324 & ~n11332 ) ;
  assign n11336 = n11332 ^ n11324 ^ n11180 ;
  assign n11337 = n11334 ^ x59 ^ 1'b0 ;
  assign n11338 = ( n11182 & ~n11336 ) | ( n11182 & n11337 ) | ( ~n11336 & n11337 ) ;
  assign n11339 = n11337 ^ n11336 ^ n11182 ;
  assign n11340 = x88 & ~n242 ;
  assign n11341 = x87 & n325 ;
  assign n11342 = ( x88 & ~n11340 ) | ( x88 & n11341 ) | ( ~n11340 & n11341 ) ;
  assign n11343 = ( ~x23 & n11332 ) | ( ~x23 & n11342 ) | ( n11332 & n11342 ) ;
  assign n11344 = n11342 ^ n11332 ^ x23 ;
  assign n11345 = ( n11104 & n11335 ) | ( n11104 & ~n11344 ) | ( n11335 & ~n11344 ) ;
  assign n11346 = n11344 ^ n11335 ^ n11104 ;
  assign n11347 = x94 & n263 ;
  assign n11348 = ( x96 & n264 ) | ( x96 & n11347 ) | ( n264 & n11347 ) ;
  assign n11349 = n11347 | n11348 ;
  assign n11350 = x95 & ~n260 ;
  assign n11351 = ( x95 & n11349 ) | ( x95 & ~n11350 ) | ( n11349 & ~n11350 ) ;
  assign n11352 = n272 & n2907 ;
  assign n11353 = n11351 | n11352 ;
  assign n11354 = n11353 ^ x56 ^ 1'b0 ;
  assign n11355 = ( n11184 & ~n11339 ) | ( n11184 & n11354 ) | ( ~n11339 & n11354 ) ;
  assign n11356 = n11354 ^ n11339 ^ n11184 ;
  assign n11357 = x97 & n408 ;
  assign n11358 = ( x99 & n403 ) | ( x99 & n11357 ) | ( n403 & n11357 ) ;
  assign n11359 = n11357 | n11358 ;
  assign n11360 = x98 & ~n410 ;
  assign n11361 = ( x98 & n11359 ) | ( x98 & ~n11360 ) | ( n11359 & ~n11360 ) ;
  assign n11362 = n402 & n4270 ;
  assign n11363 = n11361 | n11362 ;
  assign n11364 = n11363 ^ x53 ^ 1'b0 ;
  assign n11365 = n11364 ^ n11356 ^ n11195 ;
  assign n11366 = ( n11195 & ~n11356 ) | ( n11195 & n11364 ) | ( ~n11356 & n11364 ) ;
  assign n11367 = x100 & n561 ;
  assign n11368 = ( x102 & n551 ) | ( x102 & n11367 ) | ( n551 & n11367 ) ;
  assign n11369 = n11367 | n11368 ;
  assign n11370 = x101 & ~n550 ;
  assign n11371 = ( x101 & n11369 ) | ( x101 & ~n11370 ) | ( n11369 & ~n11370 ) ;
  assign n11372 = n553 & n5947 ;
  assign n11373 = n11371 | n11372 ;
  assign n11374 = n11373 ^ x50 ^ 1'b0 ;
  assign n11375 = n11374 ^ n11365 ^ n11204 ;
  assign n11376 = ( n11204 & ~n11365 ) | ( n11204 & n11374 ) | ( ~n11365 & n11374 ) ;
  assign n11377 = x103 & n744 ;
  assign n11378 = ( x105 & n730 ) | ( x105 & n11377 ) | ( n730 & n11377 ) ;
  assign n11379 = n11377 | n11378 ;
  assign n11380 = x104 & ~n732 ;
  assign n11381 = ( x104 & n11379 ) | ( x104 & ~n11380 ) | ( n11379 & ~n11380 ) ;
  assign n11382 = n731 & n8105 ;
  assign n11383 = n11381 | n11382 ;
  assign n11384 = n11383 ^ x47 ^ 1'b0 ;
  assign n11385 = ( n11215 & ~n11375 ) | ( n11215 & n11384 ) | ( ~n11375 & n11384 ) ;
  assign n11386 = n11384 ^ n11375 ^ n11215 ;
  assign n11387 = x106 & n888 ;
  assign n11388 = ( x108 & n878 ) | ( x108 & n11387 ) | ( n878 & n11387 ) ;
  assign n11389 = n11387 | n11388 ;
  assign n11390 = x107 & ~n877 ;
  assign n11391 = ( x107 & n11389 ) | ( x107 & ~n11390 ) | ( n11389 & ~n11390 ) ;
  assign n11392 = n880 & n8557 ;
  assign n11393 = n11391 | n11392 ;
  assign n11394 = n11393 ^ x44 ^ 1'b0 ;
  assign n11395 = ( n11225 & ~n11386 ) | ( n11225 & n11394 ) | ( ~n11386 & n11394 ) ;
  assign n11396 = n11394 ^ n11386 ^ n11225 ;
  assign n11397 = x109 & n1058 ;
  assign n11398 = ( x111 & n1065 ) | ( x111 & n11397 ) | ( n1065 & n11397 ) ;
  assign n11399 = n11397 | n11398 ;
  assign n11400 = x110 & ~n1060 ;
  assign n11401 = ( x110 & n11399 ) | ( x110 & ~n11400 ) | ( n11399 & ~n11400 ) ;
  assign n11402 = n1063 & n8946 ;
  assign n11403 = n11401 | n11402 ;
  assign n11404 = n11403 ^ x41 ^ 1'b0 ;
  assign n11405 = n11404 ^ n11396 ^ n11234 ;
  assign n11406 = ( n11234 & ~n11396 ) | ( n11234 & n11404 ) | ( ~n11396 & n11404 ) ;
  assign n11407 = x112 & n2156 ;
  assign n11408 = ( x114 & n2163 ) | ( x114 & n11407 ) | ( n2163 & n11407 ) ;
  assign n11409 = n11407 | n11408 ;
  assign n11410 = x113 & ~n2158 ;
  assign n11411 = ( x113 & n11409 ) | ( x113 & ~n11410 ) | ( n11409 & ~n11410 ) ;
  assign n11412 = n2161 & n9279 ;
  assign n11413 = n11411 | n11412 ;
  assign n11414 = n11413 ^ x38 ^ 1'b0 ;
  assign n11415 = ( n11244 & ~n11405 ) | ( n11244 & n11414 ) | ( ~n11405 & n11414 ) ;
  assign n11416 = n11414 ^ n11405 ^ n11244 ;
  assign n11417 = x115 & n2560 ;
  assign n11418 = ( x117 & n2567 ) | ( x117 & n11417 ) | ( n2567 & n11417 ) ;
  assign n11419 = n11417 | n11418 ;
  assign n11420 = x116 & ~n2562 ;
  assign n11421 = ( x116 & n11419 ) | ( x116 & ~n11420 ) | ( n11419 & ~n11420 ) ;
  assign n11422 = n2565 & n9569 ;
  assign n11423 = n11421 | n11422 ;
  assign n11424 = n11423 ^ x35 ^ 1'b0 ;
  assign n11425 = n11424 ^ n11416 ^ n11254 ;
  assign n11426 = ( n11254 & ~n11416 ) | ( n11254 & n11424 ) | ( ~n11416 & n11424 ) ;
  assign n11427 = x118 & n3025 ;
  assign n11428 = ( x120 & n3015 ) | ( x120 & n11427 ) | ( n3015 & n11427 ) ;
  assign n11429 = n11427 | n11428 ;
  assign n11430 = x119 & ~n3014 ;
  assign n11431 = ( x119 & n11429 ) | ( x119 & ~n11430 ) | ( n11429 & ~n11430 ) ;
  assign n11432 = n3017 & n9756 ;
  assign n11433 = n11431 | n11432 ;
  assign n11434 = n11433 ^ x32 ^ 1'b0 ;
  assign n11435 = ( n11265 & n11425 ) | ( n11265 & ~n11434 ) | ( n11425 & ~n11434 ) ;
  assign n11436 = n11434 ^ n11425 ^ n11265 ;
  assign n11437 = x121 & n3344 ;
  assign n11438 = ( x123 & n3342 ) | ( x123 & n11437 ) | ( n3342 & n11437 ) ;
  assign n11439 = n11437 | n11438 ;
  assign n11440 = x122 & ~n3347 ;
  assign n11441 = ( x122 & n11439 ) | ( x122 & ~n11440 ) | ( n11439 & ~n11440 ) ;
  assign n11442 = n3346 & n9828 ;
  assign n11443 = n11441 | n11442 ;
  assign n11444 = n11443 ^ x29 ^ 1'b0 ;
  assign n11445 = n11444 ^ n11436 ^ n11275 ;
  assign n11446 = ( n11275 & n11436 ) | ( n11275 & n11444 ) | ( n11436 & n11444 ) ;
  assign n11447 = n11445 ^ n11323 ^ n11285 ;
  assign n11448 = ( n11285 & n11323 ) | ( n11285 & n11445 ) | ( n11323 & n11445 ) ;
  assign n11449 = n11447 ^ n11296 ^ n11105 ;
  assign n11450 = ( n11105 & n11296 ) | ( n11105 & n11447 ) | ( n11296 & n11447 ) ;
  assign n11451 = n11449 ^ n11302 ^ n11298 ;
  assign n11452 = ( n11298 & n11302 ) | ( n11298 & n11449 ) | ( n11302 & n11449 ) ;
  assign n11453 = x92 & n133 ;
  assign n11454 = ( x94 & n142 ) | ( x94 & n11453 ) | ( n142 & n11453 ) ;
  assign n11455 = n11453 | n11454 ;
  assign n11456 = x93 & ~n134 ;
  assign n11457 = ( x93 & n11455 ) | ( x93 & ~n11456 ) | ( n11455 & ~n11456 ) ;
  assign n11458 = n140 & n2518 ;
  assign n11459 = n11457 | n11458 ;
  assign n11460 = n11459 ^ x59 ^ 1'b0 ;
  assign n11461 = ( n11338 & ~n11346 ) | ( n11338 & n11460 ) | ( ~n11346 & n11460 ) ;
  assign n11462 = n11460 ^ n11346 ^ n11338 ;
  assign n11463 = x95 & n263 ;
  assign n11464 = ( x97 & n264 ) | ( x97 & n11463 ) | ( n264 & n11463 ) ;
  assign n11465 = n11463 | n11464 ;
  assign n11466 = x96 & ~n260 ;
  assign n11467 = ( x96 & n11465 ) | ( x96 & ~n11466 ) | ( n11465 & ~n11466 ) ;
  assign n11468 = n272 & n3668 ;
  assign n11469 = n11467 | n11468 ;
  assign n11470 = n11469 ^ x56 ^ 1'b0 ;
  assign n11471 = n11470 ^ n11462 ^ n11355 ;
  assign n11472 = ( n11355 & ~n11462 ) | ( n11355 & n11470 ) | ( ~n11462 & n11470 ) ;
  assign n11473 = x98 & n408 ;
  assign n11474 = ( x100 & n403 ) | ( x100 & n11473 ) | ( n403 & n11473 ) ;
  assign n11475 = n11473 | n11474 ;
  assign n11476 = x99 & ~n410 ;
  assign n11477 = ( x99 & n11475 ) | ( x99 & ~n11476 ) | ( n11475 & ~n11476 ) ;
  assign n11478 = n402 & n4334 ;
  assign n11479 = n11477 | n11478 ;
  assign n11480 = n11479 ^ x53 ^ 1'b0 ;
  assign n11481 = n11480 ^ n11471 ^ n11366 ;
  assign n11482 = ( n11366 & ~n11471 ) | ( n11366 & n11480 ) | ( ~n11471 & n11480 ) ;
  assign n11483 = x90 & n208 ;
  assign n11484 = ( x92 & n194 ) | ( x92 & n11483 ) | ( n194 & n11483 ) ;
  assign n11485 = n11483 | n11484 ;
  assign n11486 = x91 & ~n192 ;
  assign n11487 = ( x91 & n11485 ) | ( x91 & ~n11486 ) | ( n11485 & ~n11486 ) ;
  assign n11488 = ( n197 & n2420 ) | ( n197 & n11487 ) | ( n2420 & n11487 ) ;
  assign n11489 = n11487 | n11488 ;
  assign n11490 = x101 & n561 ;
  assign n11491 = ( x103 & n551 ) | ( x103 & n11490 ) | ( n551 & n11490 ) ;
  assign n11492 = n11490 | n11491 ;
  assign n11493 = x102 & ~n550 ;
  assign n11494 = ( x102 & n11492 ) | ( x102 & ~n11493 ) | ( n11492 & ~n11493 ) ;
  assign n11495 = n553 & n7860 ;
  assign n11496 = n11494 | n11495 ;
  assign n11497 = n11496 ^ x50 ^ 1'b0 ;
  assign n11498 = n11497 ^ n11481 ^ n11376 ;
  assign n11499 = ( n11376 & ~n11481 ) | ( n11376 & n11497 ) | ( ~n11481 & n11497 ) ;
  assign n11500 = x104 & n744 ;
  assign n11501 = ( x106 & n730 ) | ( x106 & n11500 ) | ( n730 & n11500 ) ;
  assign n11502 = n11500 | n11501 ;
  assign n11503 = x105 & ~n732 ;
  assign n11504 = ( x105 & n11502 ) | ( x105 & ~n11503 ) | ( n11502 & ~n11503 ) ;
  assign n11505 = n731 & n8287 ;
  assign n11506 = n11504 | n11505 ;
  assign n11507 = n11506 ^ x47 ^ 1'b0 ;
  assign n11508 = ( n11385 & ~n11498 ) | ( n11385 & n11507 ) | ( ~n11498 & n11507 ) ;
  assign n11509 = n11507 ^ n11498 ^ n11385 ;
  assign n11510 = x107 & n888 ;
  assign n11511 = ( x109 & n878 ) | ( x109 & n11510 ) | ( n878 & n11510 ) ;
  assign n11512 = n11510 | n11511 ;
  assign n11513 = x108 & ~n877 ;
  assign n11514 = ( x108 & n11512 ) | ( x108 & ~n11513 ) | ( n11512 & ~n11513 ) ;
  assign n11515 = n880 & n8680 ;
  assign n11516 = n11514 | n11515 ;
  assign n11517 = n11516 ^ x44 ^ 1'b0 ;
  assign n11518 = n11517 ^ n11509 ^ n11395 ;
  assign n11519 = ( n11395 & ~n11509 ) | ( n11395 & n11517 ) | ( ~n11509 & n11517 ) ;
  assign n11520 = n11489 ^ x62 ^ 1'b0 ;
  assign n11521 = x110 & n1058 ;
  assign n11522 = ( x112 & n1065 ) | ( x112 & n11521 ) | ( n1065 & n11521 ) ;
  assign n11523 = n11521 | n11522 ;
  assign n11524 = x111 & ~n1060 ;
  assign n11525 = ( x111 & n11523 ) | ( x111 & ~n11524 ) | ( n11523 & ~n11524 ) ;
  assign n11526 = n1063 & n9080 ;
  assign n11527 = n11525 | n11526 ;
  assign n11528 = n11322 ^ x26 ^ 1'b0 ;
  assign n11529 = n11527 ^ x41 ^ 1'b0 ;
  assign n11530 = ( n11406 & ~n11518 ) | ( n11406 & n11529 ) | ( ~n11518 & n11529 ) ;
  assign n11531 = n11529 ^ n11518 ^ n11406 ;
  assign n11532 = x113 & n2156 ;
  assign n11533 = ( x115 & n2163 ) | ( x115 & n11532 ) | ( n2163 & n11532 ) ;
  assign n11534 = n11532 | n11533 ;
  assign n11535 = x114 & ~n2158 ;
  assign n11536 = ( x114 & n11534 ) | ( x114 & ~n11535 ) | ( n11534 & ~n11535 ) ;
  assign n11537 = n2161 & n9414 ;
  assign n11538 = n11536 | n11537 ;
  assign n11539 = n11538 ^ x38 ^ 1'b0 ;
  assign n11540 = n11539 ^ n11531 ^ n11415 ;
  assign n11541 = ( n11415 & ~n11531 ) | ( n11415 & n11539 ) | ( ~n11531 & n11539 ) ;
  assign n11542 = x116 & n2560 ;
  assign n11543 = ( x118 & n2567 ) | ( x118 & n11542 ) | ( n2567 & n11542 ) ;
  assign n11544 = n11542 | n11543 ;
  assign n11545 = x117 & ~n2562 ;
  assign n11546 = ( x117 & n11544 ) | ( x117 & ~n11545 ) | ( n11544 & ~n11545 ) ;
  assign n11547 = n2565 & n9671 ;
  assign n11548 = n11546 | n11547 ;
  assign n11549 = n11548 ^ x35 ^ 1'b0 ;
  assign n11550 = n11549 ^ n11540 ^ n11426 ;
  assign n11551 = ( n11426 & ~n11540 ) | ( n11426 & n11549 ) | ( ~n11540 & n11549 ) ;
  assign n11552 = x119 & n3025 ;
  assign n11553 = ( x121 & n3015 ) | ( x121 & n11552 ) | ( n3015 & n11552 ) ;
  assign n11554 = n11552 | n11553 ;
  assign n11555 = x120 & ~n3014 ;
  assign n11556 = ( x120 & n11554 ) | ( x120 & ~n11555 ) | ( n11554 & ~n11555 ) ;
  assign n11557 = n3017 & n9808 ;
  assign n11558 = n11556 | n11557 ;
  assign n11559 = n11558 ^ x32 ^ 1'b0 ;
  assign n11560 = ( n11435 & n11550 ) | ( n11435 & ~n11559 ) | ( n11550 & ~n11559 ) ;
  assign n11561 = n11559 ^ n11550 ^ n11435 ;
  assign n11562 = x122 & n3344 ;
  assign n11563 = ( x124 & n3342 ) | ( x124 & n11562 ) | ( n3342 & n11562 ) ;
  assign n11564 = n11562 | n11563 ;
  assign n11565 = x123 & ~n3347 ;
  assign n11566 = ( x123 & n11564 ) | ( x123 & ~n11565 ) | ( n11564 & ~n11565 ) ;
  assign n11567 = n3346 & n9858 ;
  assign n11568 = n11566 | n11567 ;
  assign n11569 = n11568 ^ x29 ^ 1'b0 ;
  assign n11570 = n11569 ^ n11561 ^ n11446 ;
  assign n11571 = ( n11446 & n11561 ) | ( n11446 & n11569 ) | ( n11561 & n11569 ) ;
  assign n11572 = ( n11448 & n11528 ) | ( n11448 & n11570 ) | ( n11528 & n11570 ) ;
  assign n11573 = n11570 ^ n11528 ^ n11448 ;
  assign n11574 = n11573 ^ n11452 ^ n11450 ;
  assign n11575 = ( n11450 & n11452 ) | ( n11450 & n11573 ) | ( n11452 & n11573 ) ;
  assign n11576 = x93 & n133 ;
  assign n11577 = x88 & n325 ;
  assign n11578 = x89 & ~n242 ;
  assign n11579 = ( x89 & n11577 ) | ( x89 & ~n11578 ) | ( n11577 & ~n11578 ) ;
  assign n11580 = ( x95 & n142 ) | ( x95 & n11576 ) | ( n142 & n11576 ) ;
  assign n11581 = n11576 | n11580 ;
  assign n11582 = x94 & ~n134 ;
  assign n11583 = ( x94 & n11581 ) | ( x94 & ~n11582 ) | ( n11581 & ~n11582 ) ;
  assign n11584 = ( n11343 & n11520 ) | ( n11343 & ~n11579 ) | ( n11520 & ~n11579 ) ;
  assign n11585 = n11579 ^ n11520 ^ n11343 ;
  assign n11586 = n140 & n2854 ;
  assign n11587 = n11583 | n11586 ;
  assign n11588 = n11587 ^ x59 ^ 1'b0 ;
  assign n11589 = n11588 ^ n11585 ^ n11345 ;
  assign n11590 = ( n11345 & ~n11585 ) | ( n11345 & n11588 ) | ( ~n11585 & n11588 ) ;
  assign n11591 = x96 & n263 ;
  assign n11592 = ( x98 & n264 ) | ( x98 & n11591 ) | ( n264 & n11591 ) ;
  assign n11593 = n11591 | n11592 ;
  assign n11594 = x97 & ~n260 ;
  assign n11595 = ( x97 & n11593 ) | ( x97 & ~n11594 ) | ( n11593 & ~n11594 ) ;
  assign n11596 = n272 & n4052 ;
  assign n11597 = n11595 | n11596 ;
  assign n11598 = n11597 ^ x56 ^ 1'b0 ;
  assign n11599 = ( n11461 & ~n11589 ) | ( n11461 & n11598 ) | ( ~n11589 & n11598 ) ;
  assign n11600 = n11598 ^ n11589 ^ n11461 ;
  assign n11601 = x99 & n408 ;
  assign n11602 = ( x101 & n403 ) | ( x101 & n11601 ) | ( n403 & n11601 ) ;
  assign n11603 = n11601 | n11602 ;
  assign n11604 = x100 & ~n410 ;
  assign n11605 = ( x100 & n11603 ) | ( x100 & ~n11604 ) | ( n11603 & ~n11604 ) ;
  assign n11606 = n402 & n5687 ;
  assign n11607 = n11605 | n11606 ;
  assign n11608 = n11607 ^ x53 ^ 1'b0 ;
  assign n11609 = ( n11472 & ~n11600 ) | ( n11472 & n11608 ) | ( ~n11600 & n11608 ) ;
  assign n11610 = n11608 ^ n11600 ^ n11472 ;
  assign n11611 = x102 & n561 ;
  assign n11612 = ( x104 & n551 ) | ( x104 & n11611 ) | ( n551 & n11611 ) ;
  assign n11613 = n11611 | n11612 ;
  assign n11614 = x103 & ~n550 ;
  assign n11615 = ( x103 & n11613 ) | ( x103 & ~n11614 ) | ( n11613 & ~n11614 ) ;
  assign n11616 = n553 & n8012 ;
  assign n11617 = n11615 | n11616 ;
  assign n11618 = n11617 ^ x50 ^ 1'b0 ;
  assign n11619 = ( n11482 & ~n11610 ) | ( n11482 & n11618 ) | ( ~n11610 & n11618 ) ;
  assign n11620 = n11618 ^ n11610 ^ n11482 ;
  assign n11621 = x105 & n744 ;
  assign n11622 = ( x107 & n730 ) | ( x107 & n11621 ) | ( n730 & n11621 ) ;
  assign n11623 = n11621 | n11622 ;
  assign n11624 = x106 & ~n732 ;
  assign n11625 = ( x106 & n11623 ) | ( x106 & ~n11624 ) | ( n11623 & ~n11624 ) ;
  assign n11626 = n731 & n8440 ;
  assign n11627 = n11625 | n11626 ;
  assign n11628 = n11627 ^ x47 ^ 1'b0 ;
  assign n11629 = n11628 ^ n11620 ^ n11499 ;
  assign n11630 = n11309 ^ x26 ^ 1'b0 ;
  assign n11631 = ( n11499 & ~n11620 ) | ( n11499 & n11628 ) | ( ~n11620 & n11628 ) ;
  assign n11632 = x108 & n888 ;
  assign n11633 = ( x110 & n878 ) | ( x110 & n11632 ) | ( n878 & n11632 ) ;
  assign n11634 = n11632 | n11633 ;
  assign n11635 = x109 & ~n877 ;
  assign n11636 = ( x109 & n11634 ) | ( x109 & ~n11635 ) | ( n11634 & ~n11635 ) ;
  assign n11637 = n880 & n8820 ;
  assign n11638 = n11636 | n11637 ;
  assign n11639 = n11638 ^ x44 ^ 1'b0 ;
  assign n11640 = ( n11508 & ~n11629 ) | ( n11508 & n11639 ) | ( ~n11629 & n11639 ) ;
  assign n11641 = n11639 ^ n11629 ^ n11508 ;
  assign n11642 = x111 & n1058 ;
  assign n11643 = ( x113 & n1065 ) | ( x113 & n11642 ) | ( n1065 & n11642 ) ;
  assign n11644 = n11642 | n11643 ;
  assign n11645 = x112 & ~n1060 ;
  assign n11646 = ( x112 & n11644 ) | ( x112 & ~n11645 ) | ( n11644 & ~n11645 ) ;
  assign n11647 = n1063 & n9199 ;
  assign n11648 = n11646 | n11647 ;
  assign n11649 = n11648 ^ x41 ^ 1'b0 ;
  assign n11650 = n11649 ^ n11641 ^ n11519 ;
  assign n11651 = ( n11519 & ~n11641 ) | ( n11519 & n11649 ) | ( ~n11641 & n11649 ) ;
  assign n11652 = x114 & n2156 ;
  assign n11653 = ( x116 & n2163 ) | ( x116 & n11652 ) | ( n2163 & n11652 ) ;
  assign n11654 = n11652 | n11653 ;
  assign n11655 = x115 & ~n2158 ;
  assign n11656 = ( x115 & n11654 ) | ( x115 & ~n11655 ) | ( n11654 & ~n11655 ) ;
  assign n11657 = n2161 & n9513 ;
  assign n11658 = n11656 | n11657 ;
  assign n11659 = n11658 ^ x38 ^ 1'b0 ;
  assign n11660 = ( n11530 & ~n11650 ) | ( n11530 & n11659 ) | ( ~n11650 & n11659 ) ;
  assign n11661 = n11659 ^ n11650 ^ n11530 ;
  assign n11662 = x117 & n2560 ;
  assign n11663 = ( x119 & n2567 ) | ( x119 & n11662 ) | ( n2567 & n11662 ) ;
  assign n11664 = n11662 | n11663 ;
  assign n11665 = x118 & ~n2562 ;
  assign n11666 = ( x118 & n11664 ) | ( x118 & ~n11665 ) | ( n11664 & ~n11665 ) ;
  assign n11667 = n2565 & n9733 ;
  assign n11668 = n11666 | n11667 ;
  assign n11669 = n11668 ^ x35 ^ 1'b0 ;
  assign n11670 = ( n11541 & ~n11661 ) | ( n11541 & n11669 ) | ( ~n11661 & n11669 ) ;
  assign n11671 = n11669 ^ n11661 ^ n11541 ;
  assign n11672 = x120 & n3025 ;
  assign n11673 = ( x122 & n3015 ) | ( x122 & n11672 ) | ( n3015 & n11672 ) ;
  assign n11674 = n11672 | n11673 ;
  assign n11675 = x121 & ~n3014 ;
  assign n11676 = ( x121 & n11674 ) | ( x121 & ~n11675 ) | ( n11674 & ~n11675 ) ;
  assign n11677 = ( n3017 & n9806 ) | ( n3017 & n11676 ) | ( n9806 & n11676 ) ;
  assign n11678 = n11676 | n11677 ;
  assign n11679 = n11678 ^ x32 ^ 1'b0 ;
  assign n11680 = ( n11551 & ~n11671 ) | ( n11551 & n11679 ) | ( ~n11671 & n11679 ) ;
  assign n11681 = n11679 ^ n11671 ^ n11551 ;
  assign n11682 = x123 & n3344 ;
  assign n11683 = ( x125 & n3342 ) | ( x125 & n11682 ) | ( n3342 & n11682 ) ;
  assign n11684 = n11682 | n11683 ;
  assign n11685 = x124 & ~n3347 ;
  assign n11686 = ( x124 & n11684 ) | ( x124 & ~n11685 ) | ( n11684 & ~n11685 ) ;
  assign n11687 = n3346 & n9883 ;
  assign n11688 = n11686 | n11687 ;
  assign n11689 = n11688 ^ x29 ^ 1'b0 ;
  assign n11690 = n11689 ^ n11681 ^ n11560 ;
  assign n11691 = ( n11560 & n11681 ) | ( n11560 & ~n11689 ) | ( n11681 & ~n11689 ) ;
  assign n11692 = ( n11571 & n11630 ) | ( n11571 & n11690 ) | ( n11630 & n11690 ) ;
  assign n11693 = n11690 ^ n11630 ^ n11571 ;
  assign n11694 = n11693 ^ n11575 ^ n11572 ;
  assign n11695 = ( n11572 & n11575 ) | ( n11572 & n11693 ) | ( n11575 & n11693 ) ;
  assign n11696 = x125 & n3344 ;
  assign n11697 = x124 & n3344 ;
  assign n11698 = ( x127 & n3342 ) | ( x127 & n11696 ) | ( n3342 & n11696 ) ;
  assign n11699 = n11696 | n11698 ;
  assign n11700 = x126 & ~n3347 ;
  assign n11701 = ( x126 & n11699 ) | ( x126 & ~n11700 ) | ( n11699 & ~n11700 ) ;
  assign n11702 = n3346 & n9949 ;
  assign n11703 = n11701 | n11702 ;
  assign n11704 = x93 & n208 ;
  assign n11705 = ( x126 & n3342 ) | ( x126 & n11697 ) | ( n3342 & n11697 ) ;
  assign n11706 = n197 & n2518 ;
  assign n11707 = n197 & n2854 ;
  assign n11708 = n11697 | n11705 ;
  assign n11709 = ( x95 & n194 ) | ( x95 & n11704 ) | ( n194 & n11704 ) ;
  assign n11710 = n11704 | n11709 ;
  assign n11711 = n11313 ^ x26 ^ 1'b0 ;
  assign n11712 = x125 & ~n3347 ;
  assign n11713 = ( x125 & n11708 ) | ( x125 & ~n11712 ) | ( n11708 & ~n11712 ) ;
  assign n11714 = x94 & ~n192 ;
  assign n11715 = x127 & ~n3347 ;
  assign n11716 = ( x94 & n11710 ) | ( x94 & ~n11714 ) | ( n11710 & ~n11714 ) ;
  assign n11717 = n3346 & n9917 ;
  assign n11718 = n11713 | n11717 ;
  assign n11719 = x91 & n208 ;
  assign n11720 = n11707 | n11716 ;
  assign n11721 = ( x93 & n194 ) | ( x93 & n11719 ) | ( n194 & n11719 ) ;
  assign n11722 = n11719 | n11721 ;
  assign n11723 = x92 & ~n192 ;
  assign n11724 = ( x92 & n11722 ) | ( x92 & ~n11723 ) | ( n11722 & ~n11723 ) ;
  assign n11725 = x126 & n3344 ;
  assign n11726 = ( x127 & ~n11715 ) | ( x127 & n11725 ) | ( ~n11715 & n11725 ) ;
  assign n11727 = ( n3346 & n9958 ) | ( n3346 & n11725 ) | ( n9958 & n11725 ) ;
  assign n11728 = x127 & n3344 ;
  assign n11729 = ( n3346 & n9968 ) | ( n3346 & n11728 ) | ( n9968 & n11728 ) ;
  assign n11730 = n11728 | n11729 ;
  assign n11731 = n11726 | n11727 ;
  assign n11732 = ( n197 & n2476 ) | ( n197 & n11724 ) | ( n2476 & n11724 ) ;
  assign n11733 = x90 & ~n242 ;
  assign n11734 = x89 & n325 ;
  assign n11735 = ( x90 & ~n11733 ) | ( x90 & n11734 ) | ( ~n11733 & n11734 ) ;
  assign n11736 = n11724 | n11732 ;
  assign n11737 = n11736 ^ x62 ^ 1'b0 ;
  assign n11738 = x94 & n133 ;
  assign n11739 = ( n11579 & ~n11735 ) | ( n11579 & n11737 ) | ( ~n11735 & n11737 ) ;
  assign n11740 = n11737 ^ n11735 ^ n11579 ;
  assign n11741 = ( x96 & n142 ) | ( x96 & n11738 ) | ( n142 & n11738 ) ;
  assign n11742 = n11738 | n11741 ;
  assign n11743 = x95 & ~n134 ;
  assign n11744 = ( x95 & n11742 ) | ( x95 & ~n11743 ) | ( n11742 & ~n11743 ) ;
  assign n11745 = n140 & n2907 ;
  assign n11746 = n11744 | n11745 ;
  assign n11747 = n11746 ^ x59 ^ 1'b0 ;
  assign n11748 = n11747 ^ n11740 ^ n11584 ;
  assign n11749 = ( n11584 & ~n11740 ) | ( n11584 & n11747 ) | ( ~n11740 & n11747 ) ;
  assign n11750 = x97 & n263 ;
  assign n11751 = ( x99 & n264 ) | ( x99 & n11750 ) | ( n264 & n11750 ) ;
  assign n11752 = n11750 | n11751 ;
  assign n11753 = x98 & ~n260 ;
  assign n11754 = ( x98 & n11752 ) | ( x98 & ~n11753 ) | ( n11752 & ~n11753 ) ;
  assign n11755 = n272 & n4270 ;
  assign n11756 = n11754 | n11755 ;
  assign n11757 = n11756 ^ x56 ^ 1'b0 ;
  assign n11758 = ( n11590 & ~n11748 ) | ( n11590 & n11757 ) | ( ~n11748 & n11757 ) ;
  assign n11759 = n11757 ^ n11748 ^ n11590 ;
  assign n11760 = x100 & n408 ;
  assign n11761 = ( x102 & n403 ) | ( x102 & n11760 ) | ( n403 & n11760 ) ;
  assign n11762 = n11760 | n11761 ;
  assign n11763 = x101 & ~n410 ;
  assign n11764 = ( x101 & n11762 ) | ( x101 & ~n11763 ) | ( n11762 & ~n11763 ) ;
  assign n11765 = n402 & n5947 ;
  assign n11766 = n11764 | n11765 ;
  assign n11767 = n11766 ^ x53 ^ 1'b0 ;
  assign n11768 = ( n11599 & ~n11759 ) | ( n11599 & n11767 ) | ( ~n11759 & n11767 ) ;
  assign n11769 = n11767 ^ n11759 ^ n11599 ;
  assign n11770 = x103 & n561 ;
  assign n11771 = ( x105 & n551 ) | ( x105 & n11770 ) | ( n551 & n11770 ) ;
  assign n11772 = n11770 | n11771 ;
  assign n11773 = x104 & ~n550 ;
  assign n11774 = ( x104 & n11772 ) | ( x104 & ~n11773 ) | ( n11772 & ~n11773 ) ;
  assign n11775 = n553 & n8105 ;
  assign n11776 = n11774 | n11775 ;
  assign n11777 = n11776 ^ x50 ^ 1'b0 ;
  assign n11778 = ( n11609 & ~n11769 ) | ( n11609 & n11777 ) | ( ~n11769 & n11777 ) ;
  assign n11779 = n11777 ^ n11769 ^ n11609 ;
  assign n11780 = x106 & n744 ;
  assign n11781 = ( x108 & n730 ) | ( x108 & n11780 ) | ( n730 & n11780 ) ;
  assign n11782 = n11780 | n11781 ;
  assign n11783 = x107 & ~n732 ;
  assign n11784 = ( x107 & n11782 ) | ( x107 & ~n11783 ) | ( n11782 & ~n11783 ) ;
  assign n11785 = n731 & n8557 ;
  assign n11786 = n11784 | n11785 ;
  assign n11787 = n11786 ^ x47 ^ 1'b0 ;
  assign n11788 = ( n11619 & ~n11779 ) | ( n11619 & n11787 ) | ( ~n11779 & n11787 ) ;
  assign n11789 = n11718 ^ x29 ^ 1'b0 ;
  assign n11790 = n11787 ^ n11779 ^ n11619 ;
  assign n11791 = x109 & n888 ;
  assign n11792 = ( x111 & n878 ) | ( x111 & n11791 ) | ( n878 & n11791 ) ;
  assign n11793 = n11791 | n11792 ;
  assign n11794 = x110 & ~n877 ;
  assign n11795 = ( x110 & n11793 ) | ( x110 & ~n11794 ) | ( n11793 & ~n11794 ) ;
  assign n11796 = n880 & n8946 ;
  assign n11797 = n11795 | n11796 ;
  assign n11798 = n11797 ^ x44 ^ 1'b0 ;
  assign n11799 = n11798 ^ n11790 ^ n11631 ;
  assign n11800 = ( n11631 & ~n11790 ) | ( n11631 & n11798 ) | ( ~n11790 & n11798 ) ;
  assign n11801 = x112 & n1058 ;
  assign n11802 = ( x114 & n1065 ) | ( x114 & n11801 ) | ( n1065 & n11801 ) ;
  assign n11803 = n11801 | n11802 ;
  assign n11804 = x113 & ~n1060 ;
  assign n11805 = ( x113 & n11803 ) | ( x113 & ~n11804 ) | ( n11803 & ~n11804 ) ;
  assign n11806 = n1063 & n9279 ;
  assign n11807 = n11805 | n11806 ;
  assign n11808 = n11807 ^ x41 ^ 1'b0 ;
  assign n11809 = ( n11640 & ~n11799 ) | ( n11640 & n11808 ) | ( ~n11799 & n11808 ) ;
  assign n11810 = n11808 ^ n11799 ^ n11640 ;
  assign n11811 = x115 & n2156 ;
  assign n11812 = ( x117 & n2163 ) | ( x117 & n11811 ) | ( n2163 & n11811 ) ;
  assign n11813 = n11811 | n11812 ;
  assign n11814 = x116 & ~n2158 ;
  assign n11815 = ( x116 & n11813 ) | ( x116 & ~n11814 ) | ( n11813 & ~n11814 ) ;
  assign n11816 = n2161 & n9569 ;
  assign n11817 = n11815 | n11816 ;
  assign n11818 = n11817 ^ x38 ^ 1'b0 ;
  assign n11819 = ( n11651 & ~n11810 ) | ( n11651 & n11818 ) | ( ~n11810 & n11818 ) ;
  assign n11820 = n11818 ^ n11810 ^ n11651 ;
  assign n11821 = x118 & n2560 ;
  assign n11822 = ( x120 & n2567 ) | ( x120 & n11821 ) | ( n2567 & n11821 ) ;
  assign n11823 = n11821 | n11822 ;
  assign n11824 = x119 & ~n2562 ;
  assign n11825 = ( x119 & n11823 ) | ( x119 & ~n11824 ) | ( n11823 & ~n11824 ) ;
  assign n11826 = n2565 & n9756 ;
  assign n11827 = n11825 | n11826 ;
  assign n11828 = n11827 ^ x35 ^ 1'b0 ;
  assign n11829 = ( n11660 & ~n11820 ) | ( n11660 & n11828 ) | ( ~n11820 & n11828 ) ;
  assign n11830 = n11828 ^ n11820 ^ n11660 ;
  assign n11831 = x121 & n3025 ;
  assign n11832 = ( x123 & n3015 ) | ( x123 & n11831 ) | ( n3015 & n11831 ) ;
  assign n11833 = n11831 | n11832 ;
  assign n11834 = x122 & ~n3014 ;
  assign n11835 = ( x122 & n11833 ) | ( x122 & ~n11834 ) | ( n11833 & ~n11834 ) ;
  assign n11836 = n3017 & n9828 ;
  assign n11837 = n11835 | n11836 ;
  assign n11838 = n11837 ^ x32 ^ 1'b0 ;
  assign n11839 = ( n11670 & ~n11830 ) | ( n11670 & n11838 ) | ( ~n11830 & n11838 ) ;
  assign n11840 = n11838 ^ n11830 ^ n11670 ;
  assign n11841 = ( n11680 & n11789 ) | ( n11680 & ~n11840 ) | ( n11789 & ~n11840 ) ;
  assign n11842 = n11840 ^ n11789 ^ n11680 ;
  assign n11843 = ( n11691 & ~n11711 ) | ( n11691 & n11842 ) | ( ~n11711 & n11842 ) ;
  assign n11844 = n11842 ^ n11711 ^ n11691 ;
  assign n11845 = ( n11692 & n11695 ) | ( n11692 & n11844 ) | ( n11695 & n11844 ) ;
  assign n11846 = n11844 ^ n11695 ^ n11692 ;
  assign n11847 = x92 & n208 ;
  assign n11848 = ( x94 & n194 ) | ( x94 & n11847 ) | ( n194 & n11847 ) ;
  assign n11849 = n11847 | n11848 ;
  assign n11850 = x93 & ~n192 ;
  assign n11851 = ( x93 & n11849 ) | ( x93 & ~n11850 ) | ( n11849 & ~n11850 ) ;
  assign n11852 = n11706 | n11851 ;
  assign n11853 = n197 & n2907 ;
  assign n11854 = x91 & ~n242 ;
  assign n11855 = x90 & n325 ;
  assign n11856 = ( x91 & ~n11854 ) | ( x91 & n11855 ) | ( ~n11854 & n11855 ) ;
  assign n11857 = n11852 ^ x62 ^ 1'b0 ;
  assign n11858 = n11856 ^ n11735 ^ x26 ;
  assign n11859 = ( ~x26 & n11735 ) | ( ~x26 & n11856 ) | ( n11735 & n11856 ) ;
  assign n11860 = ( n11739 & n11857 ) | ( n11739 & ~n11858 ) | ( n11857 & ~n11858 ) ;
  assign n11861 = n11858 ^ n11857 ^ n11739 ;
  assign n11862 = x95 & n133 ;
  assign n11863 = ( x97 & n142 ) | ( x97 & n11862 ) | ( n142 & n11862 ) ;
  assign n11864 = n11862 | n11863 ;
  assign n11865 = x96 & ~n134 ;
  assign n11866 = ( x96 & n11864 ) | ( x96 & ~n11865 ) | ( n11864 & ~n11865 ) ;
  assign n11867 = n140 & n3668 ;
  assign n11868 = n11866 | n11867 ;
  assign n11869 = n11868 ^ x59 ^ 1'b0 ;
  assign n11870 = n11869 ^ n11861 ^ n11749 ;
  assign n11871 = ( n11749 & ~n11861 ) | ( n11749 & n11869 ) | ( ~n11861 & n11869 ) ;
  assign n11872 = x94 & n208 ;
  assign n11873 = ( x96 & n194 ) | ( x96 & n11872 ) | ( n194 & n11872 ) ;
  assign n11874 = n11872 | n11873 ;
  assign n11875 = x95 & ~n192 ;
  assign n11876 = ( x95 & n11874 ) | ( x95 & ~n11875 ) | ( n11874 & ~n11875 ) ;
  assign n11877 = x98 & n263 ;
  assign n11878 = n11853 | n11876 ;
  assign n11879 = ( x100 & n264 ) | ( x100 & n11877 ) | ( n264 & n11877 ) ;
  assign n11880 = n11877 | n11879 ;
  assign n11881 = x99 & ~n260 ;
  assign n11882 = ( x99 & n11880 ) | ( x99 & ~n11881 ) | ( n11880 & ~n11881 ) ;
  assign n11883 = n272 & n4334 ;
  assign n11884 = n11882 | n11883 ;
  assign n11885 = n11884 ^ x56 ^ 1'b0 ;
  assign n11886 = n11885 ^ n11870 ^ n11758 ;
  assign n11887 = ( n11758 & ~n11870 ) | ( n11758 & n11885 ) | ( ~n11870 & n11885 ) ;
  assign n11888 = x101 & n408 ;
  assign n11889 = ( x103 & n403 ) | ( x103 & n11888 ) | ( n403 & n11888 ) ;
  assign n11890 = n11888 | n11889 ;
  assign n11891 = x102 & ~n410 ;
  assign n11892 = ( x102 & n11890 ) | ( x102 & ~n11891 ) | ( n11890 & ~n11891 ) ;
  assign n11893 = n402 & n7860 ;
  assign n11894 = n11892 | n11893 ;
  assign n11895 = n11894 ^ x53 ^ 1'b0 ;
  assign n11896 = ( n11768 & ~n11886 ) | ( n11768 & n11895 ) | ( ~n11886 & n11895 ) ;
  assign n11897 = n11895 ^ n11886 ^ n11768 ;
  assign n11898 = x104 & n561 ;
  assign n11899 = ( x106 & n551 ) | ( x106 & n11898 ) | ( n551 & n11898 ) ;
  assign n11900 = n11898 | n11899 ;
  assign n11901 = x105 & ~n550 ;
  assign n11902 = ( x105 & n11900 ) | ( x105 & ~n11901 ) | ( n11900 & ~n11901 ) ;
  assign n11903 = n553 & n8287 ;
  assign n11904 = n11902 | n11903 ;
  assign n11905 = n11904 ^ x50 ^ 1'b0 ;
  assign n11906 = n11905 ^ n11897 ^ n11778 ;
  assign n11907 = ( n11778 & ~n11897 ) | ( n11778 & n11905 ) | ( ~n11897 & n11905 ) ;
  assign n11908 = x107 & n744 ;
  assign n11909 = ( x109 & n730 ) | ( x109 & n11908 ) | ( n730 & n11908 ) ;
  assign n11910 = n11908 | n11909 ;
  assign n11911 = x108 & ~n732 ;
  assign n11912 = ( x108 & n11910 ) | ( x108 & ~n11911 ) | ( n11910 & ~n11911 ) ;
  assign n11913 = n731 & n8680 ;
  assign n11914 = n11912 | n11913 ;
  assign n11915 = n11914 ^ x47 ^ 1'b0 ;
  assign n11916 = n11915 ^ n11906 ^ n11788 ;
  assign n11917 = ( n11788 & ~n11906 ) | ( n11788 & n11915 ) | ( ~n11906 & n11915 ) ;
  assign n11918 = x110 & n888 ;
  assign n11919 = ( x112 & n878 ) | ( x112 & n11918 ) | ( n878 & n11918 ) ;
  assign n11920 = n11918 | n11919 ;
  assign n11921 = x111 & ~n877 ;
  assign n11922 = ( x111 & n11920 ) | ( x111 & ~n11921 ) | ( n11920 & ~n11921 ) ;
  assign n11923 = n880 & n9080 ;
  assign n11924 = n11922 | n11923 ;
  assign n11925 = n11924 ^ x44 ^ 1'b0 ;
  assign n11926 = ( n11800 & ~n11916 ) | ( n11800 & n11925 ) | ( ~n11916 & n11925 ) ;
  assign n11927 = n11925 ^ n11916 ^ n11800 ;
  assign n11928 = x113 & n1058 ;
  assign n11929 = ( x115 & n1065 ) | ( x115 & n11928 ) | ( n1065 & n11928 ) ;
  assign n11930 = n11928 | n11929 ;
  assign n11931 = x114 & ~n1060 ;
  assign n11932 = ( x114 & n11930 ) | ( x114 & ~n11931 ) | ( n11930 & ~n11931 ) ;
  assign n11933 = n1063 & n9414 ;
  assign n11934 = n11932 | n11933 ;
  assign n11935 = n11934 ^ x41 ^ 1'b0 ;
  assign n11936 = ( n11809 & ~n11927 ) | ( n11809 & n11935 ) | ( ~n11927 & n11935 ) ;
  assign n11937 = n11935 ^ n11927 ^ n11809 ;
  assign n11938 = x116 & n2156 ;
  assign n11939 = ( x118 & n2163 ) | ( x118 & n11938 ) | ( n2163 & n11938 ) ;
  assign n11940 = n11938 | n11939 ;
  assign n11941 = x117 & ~n2158 ;
  assign n11942 = ( x117 & n11940 ) | ( x117 & ~n11941 ) | ( n11940 & ~n11941 ) ;
  assign n11943 = n2161 & n9671 ;
  assign n11944 = n11942 | n11943 ;
  assign n11945 = n11944 ^ x38 ^ 1'b0 ;
  assign n11946 = ( n11819 & ~n11937 ) | ( n11819 & n11945 ) | ( ~n11937 & n11945 ) ;
  assign n11947 = n11945 ^ n11937 ^ n11819 ;
  assign n11948 = x119 & n2560 ;
  assign n11949 = ( x121 & n2567 ) | ( x121 & n11948 ) | ( n2567 & n11948 ) ;
  assign n11950 = n11948 | n11949 ;
  assign n11951 = x120 & ~n2562 ;
  assign n11952 = ( x120 & n11950 ) | ( x120 & ~n11951 ) | ( n11950 & ~n11951 ) ;
  assign n11953 = n2565 & n9808 ;
  assign n11954 = n11952 | n11953 ;
  assign n11955 = n11954 ^ x35 ^ 1'b0 ;
  assign n11956 = n11955 ^ n11947 ^ n11829 ;
  assign n11957 = ( n11829 & ~n11947 ) | ( n11829 & n11955 ) | ( ~n11947 & n11955 ) ;
  assign n11958 = x122 & n3025 ;
  assign n11959 = ( x124 & n3015 ) | ( x124 & n11958 ) | ( n3015 & n11958 ) ;
  assign n11960 = n11958 | n11959 ;
  assign n11961 = x123 & ~n3014 ;
  assign n11962 = ( x123 & n11960 ) | ( x123 & ~n11961 ) | ( n11960 & ~n11961 ) ;
  assign n11963 = n3017 & n9858 ;
  assign n11964 = n11703 ^ x29 ^ 1'b0 ;
  assign n11965 = n11962 | n11963 ;
  assign n11966 = n11965 ^ x32 ^ 1'b0 ;
  assign n11967 = n11966 ^ n11956 ^ n11839 ;
  assign n11968 = ( n11839 & ~n11956 ) | ( n11839 & n11966 ) | ( ~n11956 & n11966 ) ;
  assign n11969 = ( n11841 & n11964 ) | ( n11841 & ~n11967 ) | ( n11964 & ~n11967 ) ;
  assign n11970 = n11731 ^ x29 ^ 1'b0 ;
  assign n11971 = n11878 ^ x62 ^ 1'b0 ;
  assign n11972 = n11730 ^ x29 ^ 1'b0 ;
  assign n11973 = n11720 ^ x62 ^ 1'b0 ;
  assign n11974 = n11967 ^ n11964 ^ n11841 ;
  assign n11975 = n11974 ^ n11845 ^ n11843 ;
  assign n11976 = ( n11843 & ~n11845 ) | ( n11843 & n11974 ) | ( ~n11845 & n11974 ) ;
  assign n11977 = x96 & n133 ;
  assign n11978 = ( x98 & n142 ) | ( x98 & n11977 ) | ( n142 & n11977 ) ;
  assign n11979 = n11977 | n11978 ;
  assign n11980 = x97 & ~n134 ;
  assign n11981 = ( x97 & n11979 ) | ( x97 & ~n11980 ) | ( n11979 & ~n11980 ) ;
  assign n11982 = x92 & ~n242 ;
  assign n11983 = x91 & n325 ;
  assign n11984 = ( x92 & ~n11982 ) | ( x92 & n11983 ) | ( ~n11982 & n11983 ) ;
  assign n11985 = n140 & n4052 ;
  assign n11986 = n11981 | n11985 ;
  assign n11987 = n11986 ^ x59 ^ 1'b0 ;
  assign n11988 = ( n11859 & n11973 ) | ( n11859 & ~n11984 ) | ( n11973 & ~n11984 ) ;
  assign n11989 = n11984 ^ n11973 ^ n11859 ;
  assign n11990 = n11989 ^ n11987 ^ n11860 ;
  assign n11991 = ( n11860 & n11987 ) | ( n11860 & ~n11989 ) | ( n11987 & ~n11989 ) ;
  assign n11992 = x99 & n263 ;
  assign n11993 = ( x101 & n264 ) | ( x101 & n11992 ) | ( n264 & n11992 ) ;
  assign n11994 = n11992 | n11993 ;
  assign n11995 = x100 & ~n260 ;
  assign n11996 = ( x100 & n11994 ) | ( x100 & ~n11995 ) | ( n11994 & ~n11995 ) ;
  assign n11997 = n272 & n5687 ;
  assign n11998 = n11996 | n11997 ;
  assign n11999 = n11998 ^ x56 ^ 1'b0 ;
  assign n12000 = n11999 ^ n11990 ^ n11871 ;
  assign n12001 = ( n11871 & ~n11990 ) | ( n11871 & n11999 ) | ( ~n11990 & n11999 ) ;
  assign n12002 = x102 & n408 ;
  assign n12003 = ( x104 & n403 ) | ( x104 & n12002 ) | ( n403 & n12002 ) ;
  assign n12004 = n12002 | n12003 ;
  assign n12005 = x103 & ~n410 ;
  assign n12006 = ( x103 & n12004 ) | ( x103 & ~n12005 ) | ( n12004 & ~n12005 ) ;
  assign n12007 = n402 & n8012 ;
  assign n12008 = n12006 | n12007 ;
  assign n12009 = n12008 ^ x53 ^ 1'b0 ;
  assign n12010 = ( n11887 & ~n12000 ) | ( n11887 & n12009 ) | ( ~n12000 & n12009 ) ;
  assign n12011 = n12009 ^ n12000 ^ n11887 ;
  assign n12012 = x105 & n561 ;
  assign n12013 = ( x107 & n551 ) | ( x107 & n12012 ) | ( n551 & n12012 ) ;
  assign n12014 = n12012 | n12013 ;
  assign n12015 = x106 & ~n550 ;
  assign n12016 = ( x106 & n12014 ) | ( x106 & ~n12015 ) | ( n12014 & ~n12015 ) ;
  assign n12017 = n553 & n8440 ;
  assign n12018 = n12016 | n12017 ;
  assign n12019 = n12018 ^ x50 ^ 1'b0 ;
  assign n12020 = ( n11896 & ~n12011 ) | ( n11896 & n12019 ) | ( ~n12011 & n12019 ) ;
  assign n12021 = n12019 ^ n12011 ^ n11896 ;
  assign n12022 = x108 & n744 ;
  assign n12023 = ( x110 & n730 ) | ( x110 & n12022 ) | ( n730 & n12022 ) ;
  assign n12024 = n12022 | n12023 ;
  assign n12025 = x109 & ~n732 ;
  assign n12026 = ( x109 & n12024 ) | ( x109 & ~n12025 ) | ( n12024 & ~n12025 ) ;
  assign n12027 = n731 & n8820 ;
  assign n12028 = n12026 | n12027 ;
  assign n12029 = n12028 ^ x47 ^ 1'b0 ;
  assign n12030 = n12029 ^ n12021 ^ n11907 ;
  assign n12031 = ( n11907 & ~n12021 ) | ( n11907 & n12029 ) | ( ~n12021 & n12029 ) ;
  assign n12032 = x111 & n888 ;
  assign n12033 = ( x113 & n878 ) | ( x113 & n12032 ) | ( n878 & n12032 ) ;
  assign n12034 = n12032 | n12033 ;
  assign n12035 = x112 & ~n877 ;
  assign n12036 = ( x112 & n12034 ) | ( x112 & ~n12035 ) | ( n12034 & ~n12035 ) ;
  assign n12037 = n880 & n9199 ;
  assign n12038 = n12036 | n12037 ;
  assign n12039 = n12038 ^ x44 ^ 1'b0 ;
  assign n12040 = n12039 ^ n12030 ^ n11917 ;
  assign n12041 = ( n11917 & ~n12030 ) | ( n11917 & n12039 ) | ( ~n12030 & n12039 ) ;
  assign n12042 = x114 & n1058 ;
  assign n12043 = ( x116 & n1065 ) | ( x116 & n12042 ) | ( n1065 & n12042 ) ;
  assign n12044 = n12042 | n12043 ;
  assign n12045 = x115 & ~n1060 ;
  assign n12046 = ( x115 & n12044 ) | ( x115 & ~n12045 ) | ( n12044 & ~n12045 ) ;
  assign n12047 = n1063 & n9513 ;
  assign n12048 = n12046 | n12047 ;
  assign n12049 = n12048 ^ x41 ^ 1'b0 ;
  assign n12050 = ( n11926 & ~n12040 ) | ( n11926 & n12049 ) | ( ~n12040 & n12049 ) ;
  assign n12051 = n12049 ^ n12040 ^ n11926 ;
  assign n12052 = x117 & n2156 ;
  assign n12053 = ( x119 & n2163 ) | ( x119 & n12052 ) | ( n2163 & n12052 ) ;
  assign n12054 = n12052 | n12053 ;
  assign n12055 = x118 & ~n2158 ;
  assign n12056 = ( x118 & n12054 ) | ( x118 & ~n12055 ) | ( n12054 & ~n12055 ) ;
  assign n12057 = n2161 & n9733 ;
  assign n12058 = n12056 | n12057 ;
  assign n12059 = n12058 ^ x38 ^ 1'b0 ;
  assign n12060 = n12059 ^ n12051 ^ n11936 ;
  assign n12061 = ( n11936 & ~n12051 ) | ( n11936 & n12059 ) | ( ~n12051 & n12059 ) ;
  assign n12062 = x120 & n2560 ;
  assign n12063 = ( x122 & n2567 ) | ( x122 & n12062 ) | ( n2567 & n12062 ) ;
  assign n12064 = n12062 | n12063 ;
  assign n12065 = x121 & ~n2562 ;
  assign n12066 = ( x121 & n12064 ) | ( x121 & ~n12065 ) | ( n12064 & ~n12065 ) ;
  assign n12067 = n2565 & n9806 ;
  assign n12068 = n12066 | n12067 ;
  assign n12069 = n12068 ^ x35 ^ 1'b0 ;
  assign n12070 = ( n11946 & ~n12060 ) | ( n11946 & n12069 ) | ( ~n12060 & n12069 ) ;
  assign n12071 = n12069 ^ n12060 ^ n11946 ;
  assign n12072 = x123 & n3025 ;
  assign n12073 = ( x125 & n3015 ) | ( x125 & n12072 ) | ( n3015 & n12072 ) ;
  assign n12074 = n12072 | n12073 ;
  assign n12075 = x124 & ~n3014 ;
  assign n12076 = ( x124 & n12074 ) | ( x124 & ~n12075 ) | ( n12074 & ~n12075 ) ;
  assign n12077 = n3017 & n9883 ;
  assign n12078 = n12076 | n12077 ;
  assign n12079 = n12078 ^ x32 ^ 1'b0 ;
  assign n12080 = ( n11957 & ~n12071 ) | ( n11957 & n12079 ) | ( ~n12071 & n12079 ) ;
  assign n12081 = n12079 ^ n12071 ^ n11957 ;
  assign n12082 = n12081 ^ n11970 ^ n11968 ;
  assign n12083 = n12082 ^ n11976 ^ n11969 ;
  assign n12084 = ( n11968 & n11970 ) | ( n11968 & ~n12081 ) | ( n11970 & ~n12081 ) ;
  assign n12085 = ( ~n11969 & n11976 ) | ( ~n11969 & n12082 ) | ( n11976 & n12082 ) ;
  assign n12086 = x97 & n133 ;
  assign n12087 = x92 & n325 ;
  assign n12088 = x93 & ~n242 ;
  assign n12089 = ( x93 & n12087 ) | ( x93 & ~n12088 ) | ( n12087 & ~n12088 ) ;
  assign n12090 = ( x99 & n142 ) | ( x99 & n12086 ) | ( n142 & n12086 ) ;
  assign n12091 = n12086 | n12090 ;
  assign n12092 = x98 & ~n134 ;
  assign n12093 = ( x98 & n12091 ) | ( x98 & ~n12092 ) | ( n12091 & ~n12092 ) ;
  assign n12094 = ( n11984 & n11988 ) | ( n11984 & ~n12089 ) | ( n11988 & ~n12089 ) ;
  assign n12095 = n12089 ^ n11988 ^ n11984 ;
  assign n12096 = n140 & n4270 ;
  assign n12097 = n12093 | n12096 ;
  assign n12098 = n12097 ^ x59 ^ 1'b0 ;
  assign n12099 = n12098 ^ n12095 ^ n11971 ;
  assign n12100 = ( n11971 & ~n12095 ) | ( n11971 & n12098 ) | ( ~n12095 & n12098 ) ;
  assign n12101 = x100 & n263 ;
  assign n12102 = ( x102 & n264 ) | ( x102 & n12101 ) | ( n264 & n12101 ) ;
  assign n12103 = n12101 | n12102 ;
  assign n12104 = x101 & ~n260 ;
  assign n12105 = ( x101 & n12103 ) | ( x101 & ~n12104 ) | ( n12103 & ~n12104 ) ;
  assign n12106 = n272 & n5947 ;
  assign n12107 = n12105 | n12106 ;
  assign n12108 = n12107 ^ x56 ^ 1'b0 ;
  assign n12109 = ( n11991 & ~n12099 ) | ( n11991 & n12108 ) | ( ~n12099 & n12108 ) ;
  assign n12110 = n12108 ^ n12099 ^ n11991 ;
  assign n12111 = x103 & n408 ;
  assign n12112 = ( x105 & n403 ) | ( x105 & n12111 ) | ( n403 & n12111 ) ;
  assign n12113 = n12111 | n12112 ;
  assign n12114 = x104 & ~n410 ;
  assign n12115 = ( x104 & n12113 ) | ( x104 & ~n12114 ) | ( n12113 & ~n12114 ) ;
  assign n12116 = n402 & n8105 ;
  assign n12117 = n12115 | n12116 ;
  assign n12118 = n12117 ^ x53 ^ 1'b0 ;
  assign n12119 = n12118 ^ n12110 ^ n12001 ;
  assign n12120 = ( n12001 & ~n12110 ) | ( n12001 & n12118 ) | ( ~n12110 & n12118 ) ;
  assign n12121 = x106 & n561 ;
  assign n12122 = ( x108 & n551 ) | ( x108 & n12121 ) | ( n551 & n12121 ) ;
  assign n12123 = n12121 | n12122 ;
  assign n12124 = x107 & ~n550 ;
  assign n12125 = ( x107 & n12123 ) | ( x107 & ~n12124 ) | ( n12123 & ~n12124 ) ;
  assign n12126 = n553 & n8557 ;
  assign n12127 = n12125 | n12126 ;
  assign n12128 = n12127 ^ x50 ^ 1'b0 ;
  assign n12129 = ( n12010 & ~n12119 ) | ( n12010 & n12128 ) | ( ~n12119 & n12128 ) ;
  assign n12130 = n12128 ^ n12119 ^ n12010 ;
  assign n12131 = x109 & n744 ;
  assign n12132 = ( x111 & n730 ) | ( x111 & n12131 ) | ( n730 & n12131 ) ;
  assign n12133 = n12131 | n12132 ;
  assign n12134 = x110 & ~n732 ;
  assign n12135 = ( x110 & n12133 ) | ( x110 & ~n12134 ) | ( n12133 & ~n12134 ) ;
  assign n12136 = n731 & n8946 ;
  assign n12137 = n12135 | n12136 ;
  assign n12138 = n12137 ^ x47 ^ 1'b0 ;
  assign n12139 = ( n12020 & ~n12130 ) | ( n12020 & n12138 ) | ( ~n12130 & n12138 ) ;
  assign n12140 = n12138 ^ n12130 ^ n12020 ;
  assign n12141 = x112 & n888 ;
  assign n12142 = ( x114 & n878 ) | ( x114 & n12141 ) | ( n878 & n12141 ) ;
  assign n12143 = n12141 | n12142 ;
  assign n12144 = x113 & ~n877 ;
  assign n12145 = ( x113 & n12143 ) | ( x113 & ~n12144 ) | ( n12143 & ~n12144 ) ;
  assign n12146 = n880 & n9279 ;
  assign n12147 = n12145 | n12146 ;
  assign n12148 = n12147 ^ x44 ^ 1'b0 ;
  assign n12149 = n12148 ^ n12140 ^ n12031 ;
  assign n12150 = ( n12031 & ~n12140 ) | ( n12031 & n12148 ) | ( ~n12140 & n12148 ) ;
  assign n12151 = x115 & n1058 ;
  assign n12152 = ( x117 & n1065 ) | ( x117 & n12151 ) | ( n1065 & n12151 ) ;
  assign n12153 = n12151 | n12152 ;
  assign n12154 = x116 & ~n1060 ;
  assign n12155 = ( x116 & n12153 ) | ( x116 & ~n12154 ) | ( n12153 & ~n12154 ) ;
  assign n12156 = n1063 & n9569 ;
  assign n12157 = n12155 | n12156 ;
  assign n12158 = n12157 ^ x41 ^ 1'b0 ;
  assign n12159 = ( n12041 & ~n12149 ) | ( n12041 & n12158 ) | ( ~n12149 & n12158 ) ;
  assign n12160 = n12158 ^ n12149 ^ n12041 ;
  assign n12161 = x118 & n2156 ;
  assign n12162 = ( x120 & n2163 ) | ( x120 & n12161 ) | ( n2163 & n12161 ) ;
  assign n12163 = n12161 | n12162 ;
  assign n12164 = x119 & ~n2158 ;
  assign n12165 = ( x119 & n12163 ) | ( x119 & ~n12164 ) | ( n12163 & ~n12164 ) ;
  assign n12166 = n2161 & n9756 ;
  assign n12167 = n12165 | n12166 ;
  assign n12168 = n12167 ^ x38 ^ 1'b0 ;
  assign n12169 = n12168 ^ n12160 ^ n12050 ;
  assign n12170 = ( n12050 & ~n12160 ) | ( n12050 & n12168 ) | ( ~n12160 & n12168 ) ;
  assign n12171 = x125 & n3025 ;
  assign n12172 = ( x127 & n3015 ) | ( x127 & n12171 ) | ( n3015 & n12171 ) ;
  assign n12173 = n12171 | n12172 ;
  assign n12174 = x126 & ~n3014 ;
  assign n12175 = ( x126 & n12173 ) | ( x126 & ~n12174 ) | ( n12173 & ~n12174 ) ;
  assign n12176 = x124 & n3025 ;
  assign n12177 = ( x126 & n3015 ) | ( x126 & n12176 ) | ( n3015 & n12176 ) ;
  assign n12178 = n12176 | n12177 ;
  assign n12179 = n3017 & n9949 ;
  assign n12180 = n12175 | n12179 ;
  assign n12181 = x125 & ~n3014 ;
  assign n12182 = ( x125 & n12178 ) | ( x125 & ~n12181 ) | ( n12178 & ~n12181 ) ;
  assign n12183 = x127 & ~n3014 ;
  assign n12184 = x126 & n3025 ;
  assign n12185 = ( x127 & ~n12183 ) | ( x127 & n12184 ) | ( ~n12183 & n12184 ) ;
  assign n12186 = ( n3017 & n9958 ) | ( n3017 & n12184 ) | ( n9958 & n12184 ) ;
  assign n12187 = n12185 | n12186 ;
  assign n12188 = n3017 & n9917 ;
  assign n12189 = n12182 | n12188 ;
  assign n12190 = x121 & n2560 ;
  assign n12191 = x127 & n3025 ;
  assign n12192 = n12189 ^ x32 ^ 1'b0 ;
  assign n12193 = ( n3017 & n9968 ) | ( n3017 & n12191 ) | ( n9968 & n12191 ) ;
  assign n12194 = n12191 | n12193 ;
  assign n12195 = ( x123 & n2567 ) | ( x123 & n12190 ) | ( n2567 & n12190 ) ;
  assign n12196 = n12190 | n12195 ;
  assign n12197 = x122 & ~n2562 ;
  assign n12198 = ( x122 & n12196 ) | ( x122 & ~n12197 ) | ( n12196 & ~n12197 ) ;
  assign n12199 = n2565 & n9828 ;
  assign n12200 = n12198 | n12199 ;
  assign n12201 = n12200 ^ x35 ^ 1'b0 ;
  assign n12202 = n12201 ^ n12169 ^ n12061 ;
  assign n12203 = ( n12061 & ~n12169 ) | ( n12061 & n12201 ) | ( ~n12169 & n12201 ) ;
  assign n12204 = ( n12070 & n12192 ) | ( n12070 & ~n12202 ) | ( n12192 & ~n12202 ) ;
  assign n12205 = n12202 ^ n12192 ^ n12070 ;
  assign n12206 = ( n11972 & n12080 ) | ( n11972 & ~n12205 ) | ( n12080 & ~n12205 ) ;
  assign n12207 = n12205 ^ n12080 ^ n11972 ;
  assign n12208 = n12207 ^ n12085 ^ n12084 ;
  assign n12209 = ( ~n12084 & n12085 ) | ( ~n12084 & n12207 ) | ( n12085 & n12207 ) ;
  assign n12210 = x95 & n208 ;
  assign n12211 = ( x97 & n194 ) | ( x97 & n12210 ) | ( n194 & n12210 ) ;
  assign n12212 = n12210 | n12211 ;
  assign n12213 = x96 & ~n192 ;
  assign n12214 = ( x96 & n12212 ) | ( x96 & ~n12213 ) | ( n12212 & ~n12213 ) ;
  assign n12215 = n197 & n3668 ;
  assign n12216 = x93 & n325 ;
  assign n12217 = n12214 | n12215 ;
  assign n12218 = x94 & ~n242 ;
  assign n12219 = ( x94 & n12216 ) | ( x94 & ~n12218 ) | ( n12216 & ~n12218 ) ;
  assign n12220 = n12219 ^ n12089 ^ x29 ;
  assign n12221 = ( ~x29 & n12089 ) | ( ~x29 & n12219 ) | ( n12089 & n12219 ) ;
  assign n12222 = n12217 ^ x62 ^ 1'b0 ;
  assign n12223 = ( n12094 & ~n12220 ) | ( n12094 & n12222 ) | ( ~n12220 & n12222 ) ;
  assign n12224 = n12222 ^ n12220 ^ n12094 ;
  assign n12225 = x98 & n133 ;
  assign n12226 = ( x100 & n142 ) | ( x100 & n12225 ) | ( n142 & n12225 ) ;
  assign n12227 = n12225 | n12226 ;
  assign n12228 = x99 & ~n134 ;
  assign n12229 = ( x99 & n12227 ) | ( x99 & ~n12228 ) | ( n12227 & ~n12228 ) ;
  assign n12230 = n140 & n4334 ;
  assign n12231 = n12229 | n12230 ;
  assign n12232 = n12231 ^ x59 ^ 1'b0 ;
  assign n12233 = n12232 ^ n12224 ^ n12100 ;
  assign n12234 = n12180 ^ x32 ^ 1'b0 ;
  assign n12235 = ( n12100 & ~n12224 ) | ( n12100 & n12232 ) | ( ~n12224 & n12232 ) ;
  assign n12236 = x101 & n263 ;
  assign n12237 = ( x103 & n264 ) | ( x103 & n12236 ) | ( n264 & n12236 ) ;
  assign n12238 = n12236 | n12237 ;
  assign n12239 = n197 & n4334 ;
  assign n12240 = x102 & ~n260 ;
  assign n12241 = n12187 ^ x32 ^ 1'b0 ;
  assign n12242 = ( x102 & n12238 ) | ( x102 & ~n12240 ) | ( n12238 & ~n12240 ) ;
  assign n12243 = n272 & n7860 ;
  assign n12244 = n12242 | n12243 ;
  assign n12245 = n12244 ^ x56 ^ 1'b0 ;
  assign n12246 = ( n12109 & ~n12233 ) | ( n12109 & n12245 ) | ( ~n12233 & n12245 ) ;
  assign n12247 = n197 & n4270 ;
  assign n12248 = n12245 ^ n12233 ^ n12109 ;
  assign n12249 = x104 & n408 ;
  assign n12250 = ( x106 & n403 ) | ( x106 & n12249 ) | ( n403 & n12249 ) ;
  assign n12251 = n12249 | n12250 ;
  assign n12252 = x105 & ~n410 ;
  assign n12253 = ( x105 & n12251 ) | ( x105 & ~n12252 ) | ( n12251 & ~n12252 ) ;
  assign n12254 = n402 & n8287 ;
  assign n12255 = n12253 | n12254 ;
  assign n12256 = n12255 ^ x53 ^ 1'b0 ;
  assign n12257 = ( n12120 & ~n12248 ) | ( n12120 & n12256 ) | ( ~n12248 & n12256 ) ;
  assign n12258 = n12256 ^ n12248 ^ n12120 ;
  assign n12259 = x107 & n561 ;
  assign n12260 = ( x109 & n551 ) | ( x109 & n12259 ) | ( n551 & n12259 ) ;
  assign n12261 = n12259 | n12260 ;
  assign n12262 = x108 & ~n550 ;
  assign n12263 = ( x108 & n12261 ) | ( x108 & ~n12262 ) | ( n12261 & ~n12262 ) ;
  assign n12264 = n553 & n8680 ;
  assign n12265 = n12263 | n12264 ;
  assign n12266 = n12265 ^ x50 ^ 1'b0 ;
  assign n12267 = n12266 ^ n12258 ^ n12129 ;
  assign n12268 = ( n12129 & ~n12258 ) | ( n12129 & n12266 ) | ( ~n12258 & n12266 ) ;
  assign n12269 = x110 & n744 ;
  assign n12270 = ( x112 & n730 ) | ( x112 & n12269 ) | ( n730 & n12269 ) ;
  assign n12271 = n12269 | n12270 ;
  assign n12272 = x111 & ~n732 ;
  assign n12273 = ( x111 & n12271 ) | ( x111 & ~n12272 ) | ( n12271 & ~n12272 ) ;
  assign n12274 = n731 & n9080 ;
  assign n12275 = n12273 | n12274 ;
  assign n12276 = n12275 ^ x47 ^ 1'b0 ;
  assign n12277 = n12276 ^ n12267 ^ n12139 ;
  assign n12278 = ( n12139 & ~n12267 ) | ( n12139 & n12276 ) | ( ~n12267 & n12276 ) ;
  assign n12279 = x113 & n888 ;
  assign n12280 = ( x115 & n878 ) | ( x115 & n12279 ) | ( n878 & n12279 ) ;
  assign n12281 = n12279 | n12280 ;
  assign n12282 = x114 & ~n877 ;
  assign n12283 = ( x114 & n12281 ) | ( x114 & ~n12282 ) | ( n12281 & ~n12282 ) ;
  assign n12284 = n880 & n9414 ;
  assign n12285 = n12283 | n12284 ;
  assign n12286 = n12285 ^ x44 ^ 1'b0 ;
  assign n12287 = n12286 ^ n12277 ^ n12150 ;
  assign n12288 = ( n12150 & ~n12277 ) | ( n12150 & n12286 ) | ( ~n12277 & n12286 ) ;
  assign n12289 = x116 & n1058 ;
  assign n12290 = ( x118 & n1065 ) | ( x118 & n12289 ) | ( n1065 & n12289 ) ;
  assign n12291 = n12289 | n12290 ;
  assign n12292 = x117 & ~n1060 ;
  assign n12293 = ( x117 & n12291 ) | ( x117 & ~n12292 ) | ( n12291 & ~n12292 ) ;
  assign n12294 = n1063 & n9671 ;
  assign n12295 = n12293 | n12294 ;
  assign n12296 = n12295 ^ x41 ^ 1'b0 ;
  assign n12297 = ( n12159 & ~n12287 ) | ( n12159 & n12296 ) | ( ~n12287 & n12296 ) ;
  assign n12298 = n12296 ^ n12287 ^ n12159 ;
  assign n12299 = x119 & n2156 ;
  assign n12300 = ( x121 & n2163 ) | ( x121 & n12299 ) | ( n2163 & n12299 ) ;
  assign n12301 = n12299 | n12300 ;
  assign n12302 = x120 & ~n2158 ;
  assign n12303 = ( x120 & n12301 ) | ( x120 & ~n12302 ) | ( n12301 & ~n12302 ) ;
  assign n12304 = n2161 & n9808 ;
  assign n12305 = n12303 | n12304 ;
  assign n12306 = n12305 ^ x38 ^ 1'b0 ;
  assign n12307 = ( n12170 & ~n12298 ) | ( n12170 & n12306 ) | ( ~n12298 & n12306 ) ;
  assign n12308 = n12306 ^ n12298 ^ n12170 ;
  assign n12309 = n197 & n4052 ;
  assign n12310 = x98 & n208 ;
  assign n12311 = ( x100 & n194 ) | ( x100 & n12310 ) | ( n194 & n12310 ) ;
  assign n12312 = n12310 | n12311 ;
  assign n12313 = x99 & ~n192 ;
  assign n12314 = ( x99 & n12312 ) | ( x99 & ~n12313 ) | ( n12312 & ~n12313 ) ;
  assign n12315 = x122 & n2560 ;
  assign n12316 = n12239 | n12314 ;
  assign n12317 = ( x124 & n2567 ) | ( x124 & n12315 ) | ( n2567 & n12315 ) ;
  assign n12318 = n12315 | n12317 ;
  assign n12319 = x123 & ~n2562 ;
  assign n12320 = ( x123 & n12318 ) | ( x123 & ~n12319 ) | ( n12318 & ~n12319 ) ;
  assign n12321 = n2565 & n9858 ;
  assign n12322 = n12320 | n12321 ;
  assign n12323 = n12322 ^ x35 ^ 1'b0 ;
  assign n12324 = n12316 ^ x62 ^ 1'b0 ;
  assign n12325 = ( n12203 & ~n12308 ) | ( n12203 & n12323 ) | ( ~n12308 & n12323 ) ;
  assign n12326 = n12323 ^ n12308 ^ n12203 ;
  assign n12327 = x96 & n208 ;
  assign n12328 = ( x98 & n194 ) | ( x98 & n12327 ) | ( n194 & n12327 ) ;
  assign n12329 = n12327 | n12328 ;
  assign n12330 = x97 & ~n192 ;
  assign n12331 = ( x97 & n12329 ) | ( x97 & ~n12330 ) | ( n12329 & ~n12330 ) ;
  assign n12332 = n12326 ^ n12234 ^ n12204 ;
  assign n12333 = n12309 | n12331 ;
  assign n12334 = ( ~n12206 & n12209 ) | ( ~n12206 & n12332 ) | ( n12209 & n12332 ) ;
  assign n12335 = n12332 ^ n12209 ^ n12206 ;
  assign n12336 = n12333 ^ x62 ^ 1'b0 ;
  assign n12337 = ( n12204 & n12234 ) | ( n12204 & ~n12326 ) | ( n12234 & ~n12326 ) ;
  assign n12338 = x97 & n208 ;
  assign n12339 = x98 & ~n192 ;
  assign n12340 = ( x99 & n194 ) | ( x99 & n12338 ) | ( n194 & n12338 ) ;
  assign n12341 = n12338 | n12340 ;
  assign n12342 = ( x98 & ~n12339 ) | ( x98 & n12341 ) | ( ~n12339 & n12341 ) ;
  assign n12343 = x99 & n133 ;
  assign n12344 = ( x101 & n142 ) | ( x101 & n12343 ) | ( n142 & n12343 ) ;
  assign n12345 = n12343 | n12344 ;
  assign n12346 = n12247 | n12342 ;
  assign n12347 = n140 & n5687 ;
  assign n12348 = x100 & ~n134 ;
  assign n12349 = ( x100 & n12345 ) | ( x100 & ~n12348 ) | ( n12345 & ~n12348 ) ;
  assign n12350 = n12347 | n12349 ;
  assign n12351 = x94 & n325 ;
  assign n12352 = x95 & ~n242 ;
  assign n12353 = ( x95 & n12351 ) | ( x95 & ~n12352 ) | ( n12351 & ~n12352 ) ;
  assign n12354 = n12353 ^ n12336 ^ n12221 ;
  assign n12355 = n12350 ^ x59 ^ 1'b0 ;
  assign n12356 = ( n12221 & n12336 ) | ( n12221 & ~n12353 ) | ( n12336 & ~n12353 ) ;
  assign n12357 = n12355 ^ n12354 ^ n12223 ;
  assign n12358 = ( n12223 & ~n12354 ) | ( n12223 & n12355 ) | ( ~n12354 & n12355 ) ;
  assign n12359 = x102 & n263 ;
  assign n12360 = ( x104 & n264 ) | ( x104 & n12359 ) | ( n264 & n12359 ) ;
  assign n12361 = n12359 | n12360 ;
  assign n12362 = x103 & ~n260 ;
  assign n12363 = ( x103 & n12361 ) | ( x103 & ~n12362 ) | ( n12361 & ~n12362 ) ;
  assign n12364 = n272 & n8012 ;
  assign n12365 = n12363 | n12364 ;
  assign n12366 = n12365 ^ x56 ^ 1'b0 ;
  assign n12367 = n12366 ^ n12357 ^ n12235 ;
  assign n12368 = ( n12235 & ~n12357 ) | ( n12235 & n12366 ) | ( ~n12357 & n12366 ) ;
  assign n12369 = x105 & n408 ;
  assign n12370 = ( x107 & n403 ) | ( x107 & n12369 ) | ( n403 & n12369 ) ;
  assign n12371 = n12369 | n12370 ;
  assign n12372 = x106 & ~n410 ;
  assign n12373 = ( x106 & n12371 ) | ( x106 & ~n12372 ) | ( n12371 & ~n12372 ) ;
  assign n12374 = n402 & n8440 ;
  assign n12375 = n12373 | n12374 ;
  assign n12376 = n12375 ^ x53 ^ 1'b0 ;
  assign n12377 = n12376 ^ n12367 ^ n12246 ;
  assign n12378 = ( n12246 & ~n12367 ) | ( n12246 & n12376 ) | ( ~n12367 & n12376 ) ;
  assign n12379 = x108 & n561 ;
  assign n12380 = ( x110 & n551 ) | ( x110 & n12379 ) | ( n551 & n12379 ) ;
  assign n12381 = n12379 | n12380 ;
  assign n12382 = x109 & ~n550 ;
  assign n12383 = ( x109 & n12381 ) | ( x109 & ~n12382 ) | ( n12381 & ~n12382 ) ;
  assign n12384 = n553 & n8820 ;
  assign n12385 = n12383 | n12384 ;
  assign n12386 = n12385 ^ x50 ^ 1'b0 ;
  assign n12387 = n12386 ^ n12377 ^ n12257 ;
  assign n12388 = ( n12257 & ~n12377 ) | ( n12257 & n12386 ) | ( ~n12377 & n12386 ) ;
  assign n12389 = x111 & n744 ;
  assign n12390 = ( x113 & n730 ) | ( x113 & n12389 ) | ( n730 & n12389 ) ;
  assign n12391 = n12389 | n12390 ;
  assign n12392 = x112 & ~n732 ;
  assign n12393 = ( x112 & n12391 ) | ( x112 & ~n12392 ) | ( n12391 & ~n12392 ) ;
  assign n12394 = n731 & n9199 ;
  assign n12395 = n12393 | n12394 ;
  assign n12396 = n12395 ^ x47 ^ 1'b0 ;
  assign n12397 = n12396 ^ n12387 ^ n12268 ;
  assign n12398 = ( n12268 & ~n12387 ) | ( n12268 & n12396 ) | ( ~n12387 & n12396 ) ;
  assign n12399 = x114 & n888 ;
  assign n12400 = ( x116 & n878 ) | ( x116 & n12399 ) | ( n878 & n12399 ) ;
  assign n12401 = n12399 | n12400 ;
  assign n12402 = x115 & ~n877 ;
  assign n12403 = ( x115 & n12401 ) | ( x115 & ~n12402 ) | ( n12401 & ~n12402 ) ;
  assign n12404 = n880 & n9513 ;
  assign n12405 = n12403 | n12404 ;
  assign n12406 = n12405 ^ x44 ^ 1'b0 ;
  assign n12407 = ( n12278 & ~n12397 ) | ( n12278 & n12406 ) | ( ~n12397 & n12406 ) ;
  assign n12408 = n12406 ^ n12397 ^ n12278 ;
  assign n12409 = x117 & n1058 ;
  assign n12410 = ( x119 & n1065 ) | ( x119 & n12409 ) | ( n1065 & n12409 ) ;
  assign n12411 = n12409 | n12410 ;
  assign n12412 = x118 & ~n1060 ;
  assign n12413 = ( x118 & n12411 ) | ( x118 & ~n12412 ) | ( n12411 & ~n12412 ) ;
  assign n12414 = n1063 & n9733 ;
  assign n12415 = n12413 | n12414 ;
  assign n12416 = n12415 ^ x41 ^ 1'b0 ;
  assign n12417 = n12416 ^ n12408 ^ n12288 ;
  assign n12418 = ( n12288 & ~n12408 ) | ( n12288 & n12416 ) | ( ~n12408 & n12416 ) ;
  assign n12419 = x120 & n2156 ;
  assign n12420 = ( x122 & n2163 ) | ( x122 & n12419 ) | ( n2163 & n12419 ) ;
  assign n12421 = n12419 | n12420 ;
  assign n12422 = x121 & ~n2158 ;
  assign n12423 = ( x121 & n12421 ) | ( x121 & ~n12422 ) | ( n12421 & ~n12422 ) ;
  assign n12424 = n2161 & n9806 ;
  assign n12425 = n12423 | n12424 ;
  assign n12426 = n12425 ^ x38 ^ 1'b0 ;
  assign n12427 = ( n12297 & ~n12417 ) | ( n12297 & n12426 ) | ( ~n12417 & n12426 ) ;
  assign n12428 = n12426 ^ n12417 ^ n12297 ;
  assign n12429 = x123 & n2560 ;
  assign n12430 = ( x125 & n2567 ) | ( x125 & n12429 ) | ( n2567 & n12429 ) ;
  assign n12431 = n12429 | n12430 ;
  assign n12432 = x124 & ~n2562 ;
  assign n12433 = ( x124 & n12431 ) | ( x124 & ~n12432 ) | ( n12431 & ~n12432 ) ;
  assign n12434 = n2565 & n9883 ;
  assign n12435 = n12433 | n12434 ;
  assign n12436 = n12435 ^ x35 ^ 1'b0 ;
  assign n12437 = ( n12307 & ~n12428 ) | ( n12307 & n12436 ) | ( ~n12428 & n12436 ) ;
  assign n12438 = n12436 ^ n12428 ^ n12307 ;
  assign n12439 = n12438 ^ n12325 ^ n12241 ;
  assign n12440 = n12439 ^ n12337 ^ n12334 ;
  assign n12441 = ( n12241 & n12325 ) | ( n12241 & ~n12438 ) | ( n12325 & ~n12438 ) ;
  assign n12442 = ( n12334 & ~n12337 ) | ( n12334 & n12439 ) | ( ~n12337 & n12439 ) ;
  assign n12443 = x95 & n325 ;
  assign n12444 = x96 & ~n242 ;
  assign n12445 = ( x96 & n12443 ) | ( x96 & ~n12444 ) | ( n12443 & ~n12444 ) ;
  assign n12446 = x100 & n133 ;
  assign n12447 = ( x102 & n142 ) | ( x102 & n12446 ) | ( n142 & n12446 ) ;
  assign n12448 = n12446 | n12447 ;
  assign n12449 = x101 & ~n134 ;
  assign n12450 = ( x101 & n12448 ) | ( x101 & ~n12449 ) | ( n12448 & ~n12449 ) ;
  assign n12451 = n12346 ^ x62 ^ 1'b0 ;
  assign n12452 = n140 & n5947 ;
  assign n12453 = n12450 | n12452 ;
  assign n12454 = n12453 ^ x59 ^ 1'b0 ;
  assign n12455 = n12445 ^ n12356 ^ n12353 ;
  assign n12456 = ( n12353 & n12356 ) | ( n12353 & ~n12445 ) | ( n12356 & ~n12445 ) ;
  assign n12457 = n12455 ^ n12454 ^ n12451 ;
  assign n12458 = ( n12451 & n12454 ) | ( n12451 & ~n12455 ) | ( n12454 & ~n12455 ) ;
  assign n12459 = x103 & n263 ;
  assign n12460 = ( x105 & n264 ) | ( x105 & n12459 ) | ( n264 & n12459 ) ;
  assign n12461 = n12459 | n12460 ;
  assign n12462 = x104 & ~n260 ;
  assign n12463 = ( x104 & n12461 ) | ( x104 & ~n12462 ) | ( n12461 & ~n12462 ) ;
  assign n12464 = n272 & n8105 ;
  assign n12465 = n12463 | n12464 ;
  assign n12466 = n12465 ^ x56 ^ 1'b0 ;
  assign n12467 = ( n12358 & ~n12457 ) | ( n12358 & n12466 ) | ( ~n12457 & n12466 ) ;
  assign n12468 = n12466 ^ n12457 ^ n12358 ;
  assign n12469 = x106 & n408 ;
  assign n12470 = ( x108 & n403 ) | ( x108 & n12469 ) | ( n403 & n12469 ) ;
  assign n12471 = n12469 | n12470 ;
  assign n12472 = x107 & ~n410 ;
  assign n12473 = ( x107 & n12471 ) | ( x107 & ~n12472 ) | ( n12471 & ~n12472 ) ;
  assign n12474 = n402 & n8557 ;
  assign n12475 = n12473 | n12474 ;
  assign n12476 = n12475 ^ x53 ^ 1'b0 ;
  assign n12477 = n12476 ^ n12468 ^ n12368 ;
  assign n12478 = ( n12368 & ~n12468 ) | ( n12368 & n12476 ) | ( ~n12468 & n12476 ) ;
  assign n12479 = x109 & n561 ;
  assign n12480 = ( x111 & n551 ) | ( x111 & n12479 ) | ( n551 & n12479 ) ;
  assign n12481 = n12479 | n12480 ;
  assign n12482 = x110 & ~n550 ;
  assign n12483 = ( x110 & n12481 ) | ( x110 & ~n12482 ) | ( n12481 & ~n12482 ) ;
  assign n12484 = n553 & n8946 ;
  assign n12485 = n12483 | n12484 ;
  assign n12486 = n12485 ^ x50 ^ 1'b0 ;
  assign n12487 = n12486 ^ n12477 ^ n12378 ;
  assign n12488 = ( n12378 & ~n12477 ) | ( n12378 & n12486 ) | ( ~n12477 & n12486 ) ;
  assign n12489 = x112 & n744 ;
  assign n12490 = ( x114 & n730 ) | ( x114 & n12489 ) | ( n730 & n12489 ) ;
  assign n12491 = n12489 | n12490 ;
  assign n12492 = x113 & ~n732 ;
  assign n12493 = ( x113 & n12491 ) | ( x113 & ~n12492 ) | ( n12491 & ~n12492 ) ;
  assign n12494 = n731 & n9279 ;
  assign n12495 = n12493 | n12494 ;
  assign n12496 = n12495 ^ x47 ^ 1'b0 ;
  assign n12497 = ( n12388 & ~n12487 ) | ( n12388 & n12496 ) | ( ~n12487 & n12496 ) ;
  assign n12498 = n12496 ^ n12487 ^ n12388 ;
  assign n12499 = x115 & n888 ;
  assign n12500 = ( x117 & n878 ) | ( x117 & n12499 ) | ( n878 & n12499 ) ;
  assign n12501 = n12499 | n12500 ;
  assign n12502 = x116 & ~n877 ;
  assign n12503 = ( x116 & n12501 ) | ( x116 & ~n12502 ) | ( n12501 & ~n12502 ) ;
  assign n12504 = n880 & n9569 ;
  assign n12505 = n12503 | n12504 ;
  assign n12506 = n12505 ^ x44 ^ 1'b0 ;
  assign n12507 = n12506 ^ n12498 ^ n12398 ;
  assign n12508 = ( n12398 & ~n12498 ) | ( n12398 & n12506 ) | ( ~n12498 & n12506 ) ;
  assign n12509 = x118 & n1058 ;
  assign n12510 = ( x120 & n1065 ) | ( x120 & n12509 ) | ( n1065 & n12509 ) ;
  assign n12511 = n12509 | n12510 ;
  assign n12512 = x119 & ~n1060 ;
  assign n12513 = ( x119 & n12511 ) | ( x119 & ~n12512 ) | ( n12511 & ~n12512 ) ;
  assign n12514 = n1063 & n9756 ;
  assign n12515 = n12513 | n12514 ;
  assign n12516 = n12515 ^ x41 ^ 1'b0 ;
  assign n12517 = n12516 ^ n12507 ^ n12407 ;
  assign n12518 = ( n12407 & ~n12507 ) | ( n12407 & n12516 ) | ( ~n12507 & n12516 ) ;
  assign n12519 = x121 & n2156 ;
  assign n12520 = ( x123 & n2163 ) | ( x123 & n12519 ) | ( n2163 & n12519 ) ;
  assign n12521 = n12519 | n12520 ;
  assign n12522 = x122 & ~n2158 ;
  assign n12523 = ( x122 & n12521 ) | ( x122 & ~n12522 ) | ( n12521 & ~n12522 ) ;
  assign n12524 = n2161 & n9828 ;
  assign n12525 = n12523 | n12524 ;
  assign n12526 = n12525 ^ x38 ^ 1'b0 ;
  assign n12527 = n12526 ^ n12517 ^ n12418 ;
  assign n12528 = ( n12418 & ~n12517 ) | ( n12418 & n12526 ) | ( ~n12517 & n12526 ) ;
  assign n12529 = n12194 ^ x32 ^ 1'b0 ;
  assign n12530 = x125 & n2560 ;
  assign n12531 = ( x127 & n2567 ) | ( x127 & n12530 ) | ( n2567 & n12530 ) ;
  assign n12532 = n12530 | n12531 ;
  assign n12533 = x124 & n2560 ;
  assign n12534 = ( x126 & n2567 ) | ( x126 & n12533 ) | ( n2567 & n12533 ) ;
  assign n12535 = n12533 | n12534 ;
  assign n12536 = x126 & ~n2562 ;
  assign n12537 = ( x126 & n12532 ) | ( x126 & ~n12536 ) | ( n12532 & ~n12536 ) ;
  assign n12538 = n2565 & n9949 ;
  assign n12539 = n12537 | n12538 ;
  assign n12540 = x127 & ~n2562 ;
  assign n12541 = x125 & ~n2562 ;
  assign n12542 = ( x125 & n12535 ) | ( x125 & ~n12541 ) | ( n12535 & ~n12541 ) ;
  assign n12543 = x126 & n2560 ;
  assign n12544 = ( x127 & ~n12540 ) | ( x127 & n12543 ) | ( ~n12540 & n12543 ) ;
  assign n12545 = ( n2565 & n9958 ) | ( n2565 & n12543 ) | ( n9958 & n12543 ) ;
  assign n12546 = n12544 | n12545 ;
  assign n12547 = x127 & n2560 ;
  assign n12548 = n2565 & n9917 ;
  assign n12549 = n12542 | n12548 ;
  assign n12550 = n12549 ^ x35 ^ 1'b0 ;
  assign n12551 = n12550 ^ n12527 ^ n12427 ;
  assign n12552 = ( n12427 & ~n12527 ) | ( n12427 & n12550 ) | ( ~n12527 & n12550 ) ;
  assign n12553 = ( n12437 & n12529 ) | ( n12437 & ~n12551 ) | ( n12529 & ~n12551 ) ;
  assign n12554 = n12551 ^ n12529 ^ n12437 ;
  assign n12555 = ( ~n12441 & n12442 ) | ( ~n12441 & n12554 ) | ( n12442 & n12554 ) ;
  assign n12556 = n12554 ^ n12442 ^ n12441 ;
  assign n12557 = x97 & ~n242 ;
  assign n12558 = ( n2565 & n9968 ) | ( n2565 & n12547 ) | ( n9968 & n12547 ) ;
  assign n12559 = n12547 | n12558 ;
  assign n12560 = x96 & n325 ;
  assign n12561 = ( x97 & ~n12557 ) | ( x97 & n12560 ) | ( ~n12557 & n12560 ) ;
  assign n12562 = ( ~x32 & n12445 ) | ( ~x32 & n12561 ) | ( n12445 & n12561 ) ;
  assign n12563 = n12561 ^ n12445 ^ x32 ;
  assign n12564 = n12563 ^ n12456 ^ n12324 ;
  assign n12565 = ( n12324 & n12456 ) | ( n12324 & ~n12563 ) | ( n12456 & ~n12563 ) ;
  assign n12566 = x101 & n133 ;
  assign n12567 = ( x103 & n142 ) | ( x103 & n12566 ) | ( n142 & n12566 ) ;
  assign n12568 = n12566 | n12567 ;
  assign n12569 = x102 & ~n134 ;
  assign n12570 = ( x102 & n12568 ) | ( x102 & ~n12569 ) | ( n12568 & ~n12569 ) ;
  assign n12571 = n140 & n7860 ;
  assign n12572 = n12570 | n12571 ;
  assign n12573 = n12572 ^ x59 ^ 1'b0 ;
  assign n12574 = n12573 ^ n12564 ^ n12458 ;
  assign n12575 = ( n12458 & ~n12564 ) | ( n12458 & n12573 ) | ( ~n12564 & n12573 ) ;
  assign n12576 = x104 & n263 ;
  assign n12577 = ( x106 & n264 ) | ( x106 & n12576 ) | ( n264 & n12576 ) ;
  assign n12578 = n12576 | n12577 ;
  assign n12579 = x105 & ~n260 ;
  assign n12580 = ( x105 & n12578 ) | ( x105 & ~n12579 ) | ( n12578 & ~n12579 ) ;
  assign n12581 = n272 & n8287 ;
  assign n12582 = n12580 | n12581 ;
  assign n12583 = n12582 ^ x56 ^ 1'b0 ;
  assign n12584 = ( n12467 & ~n12574 ) | ( n12467 & n12583 ) | ( ~n12574 & n12583 ) ;
  assign n12585 = n12583 ^ n12574 ^ n12467 ;
  assign n12586 = x107 & n408 ;
  assign n12587 = ( x109 & n403 ) | ( x109 & n12586 ) | ( n403 & n12586 ) ;
  assign n12588 = n12586 | n12587 ;
  assign n12589 = x108 & ~n410 ;
  assign n12590 = ( x108 & n12588 ) | ( x108 & ~n12589 ) | ( n12588 & ~n12589 ) ;
  assign n12591 = n402 & n8680 ;
  assign n12592 = n12590 | n12591 ;
  assign n12593 = n12592 ^ x53 ^ 1'b0 ;
  assign n12594 = n12593 ^ n12585 ^ n12478 ;
  assign n12595 = ( n12478 & ~n12585 ) | ( n12478 & n12593 ) | ( ~n12585 & n12593 ) ;
  assign n12596 = x110 & n561 ;
  assign n12597 = ( x112 & n551 ) | ( x112 & n12596 ) | ( n551 & n12596 ) ;
  assign n12598 = n12596 | n12597 ;
  assign n12599 = x111 & ~n550 ;
  assign n12600 = ( x111 & n12598 ) | ( x111 & ~n12599 ) | ( n12598 & ~n12599 ) ;
  assign n12601 = n553 & n9080 ;
  assign n12602 = n12600 | n12601 ;
  assign n12603 = n12539 ^ x35 ^ 1'b0 ;
  assign n12604 = n12602 ^ x50 ^ 1'b0 ;
  assign n12605 = n12604 ^ n12594 ^ n12488 ;
  assign n12606 = ( n12488 & ~n12594 ) | ( n12488 & n12604 ) | ( ~n12594 & n12604 ) ;
  assign n12607 = x113 & n744 ;
  assign n12608 = ( x115 & n730 ) | ( x115 & n12607 ) | ( n730 & n12607 ) ;
  assign n12609 = n12607 | n12608 ;
  assign n12610 = x114 & ~n732 ;
  assign n12611 = ( x114 & n12609 ) | ( x114 & ~n12610 ) | ( n12609 & ~n12610 ) ;
  assign n12612 = n731 & n9414 ;
  assign n12613 = n12611 | n12612 ;
  assign n12614 = n12613 ^ x47 ^ 1'b0 ;
  assign n12615 = n12614 ^ n12605 ^ n12497 ;
  assign n12616 = ( n12497 & ~n12605 ) | ( n12497 & n12614 ) | ( ~n12605 & n12614 ) ;
  assign n12617 = x116 & n888 ;
  assign n12618 = ( x118 & n878 ) | ( x118 & n12617 ) | ( n878 & n12617 ) ;
  assign n12619 = n12617 | n12618 ;
  assign n12620 = x117 & ~n877 ;
  assign n12621 = ( x117 & n12619 ) | ( x117 & ~n12620 ) | ( n12619 & ~n12620 ) ;
  assign n12622 = n880 & n9671 ;
  assign n12623 = n12621 | n12622 ;
  assign n12624 = n12623 ^ x44 ^ 1'b0 ;
  assign n12625 = n12624 ^ n12615 ^ n12508 ;
  assign n12626 = ( n12508 & ~n12615 ) | ( n12508 & n12624 ) | ( ~n12615 & n12624 ) ;
  assign n12627 = x119 & n1058 ;
  assign n12628 = ( x121 & n1065 ) | ( x121 & n12627 ) | ( n1065 & n12627 ) ;
  assign n12629 = n12627 | n12628 ;
  assign n12630 = x120 & ~n1060 ;
  assign n12631 = ( x120 & n12629 ) | ( x120 & ~n12630 ) | ( n12629 & ~n12630 ) ;
  assign n12632 = n1063 & n9808 ;
  assign n12633 = n12631 | n12632 ;
  assign n12634 = n12633 ^ x41 ^ 1'b0 ;
  assign n12635 = n12634 ^ n12625 ^ n12518 ;
  assign n12636 = ( n12518 & ~n12625 ) | ( n12518 & n12634 ) | ( ~n12625 & n12634 ) ;
  assign n12637 = x122 & n2156 ;
  assign n12638 = ( x124 & n2163 ) | ( x124 & n12637 ) | ( n2163 & n12637 ) ;
  assign n12639 = n12637 | n12638 ;
  assign n12640 = x123 & ~n2158 ;
  assign n12641 = ( x123 & n12639 ) | ( x123 & ~n12640 ) | ( n12639 & ~n12640 ) ;
  assign n12642 = n2161 & n9858 ;
  assign n12643 = n12641 | n12642 ;
  assign n12644 = n12643 ^ x38 ^ 1'b0 ;
  assign n12645 = ( n12528 & ~n12635 ) | ( n12528 & n12644 ) | ( ~n12635 & n12644 ) ;
  assign n12646 = n12644 ^ n12635 ^ n12528 ;
  assign n12647 = n12646 ^ n12603 ^ n12552 ;
  assign n12648 = ( n12552 & n12603 ) | ( n12552 & ~n12646 ) | ( n12603 & ~n12646 ) ;
  assign n12649 = n12647 ^ n12555 ^ n12553 ;
  assign n12650 = ( ~n12553 & n12555 ) | ( ~n12553 & n12647 ) | ( n12555 & n12647 ) ;
  assign n12651 = x99 & n208 ;
  assign n12652 = ( x101 & n194 ) | ( x101 & n12651 ) | ( n194 & n12651 ) ;
  assign n12653 = n197 & n5687 ;
  assign n12654 = n12651 | n12652 ;
  assign n12655 = x100 & ~n192 ;
  assign n12656 = ( x100 & n12654 ) | ( x100 & ~n12655 ) | ( n12654 & ~n12655 ) ;
  assign n12657 = x102 & n133 ;
  assign n12658 = n12653 | n12656 ;
  assign n12659 = x97 & n325 ;
  assign n12660 = ( x104 & n142 ) | ( x104 & n12657 ) | ( n142 & n12657 ) ;
  assign n12661 = n12657 | n12660 ;
  assign n12662 = x98 & ~n242 ;
  assign n12663 = ( x98 & n12659 ) | ( x98 & ~n12662 ) | ( n12659 & ~n12662 ) ;
  assign n12664 = n12658 ^ x62 ^ 1'b0 ;
  assign n12665 = n12664 ^ n12663 ^ n12562 ;
  assign n12666 = ( n12562 & ~n12663 ) | ( n12562 & n12664 ) | ( ~n12663 & n12664 ) ;
  assign n12667 = x103 & ~n134 ;
  assign n12668 = ( x103 & n12661 ) | ( x103 & ~n12667 ) | ( n12661 & ~n12667 ) ;
  assign n12669 = n140 & n8012 ;
  assign n12670 = n12668 | n12669 ;
  assign n12671 = n12670 ^ x59 ^ 1'b0 ;
  assign n12672 = n12671 ^ n12665 ^ n12565 ;
  assign n12673 = n197 & n7860 ;
  assign n12674 = ( n12565 & ~n12665 ) | ( n12565 & n12671 ) | ( ~n12665 & n12671 ) ;
  assign n12675 = x105 & n263 ;
  assign n12676 = ( x107 & n264 ) | ( x107 & n12675 ) | ( n264 & n12675 ) ;
  assign n12677 = n12675 | n12676 ;
  assign n12678 = x106 & ~n260 ;
  assign n12679 = ( x106 & n12677 ) | ( x106 & ~n12678 ) | ( n12677 & ~n12678 ) ;
  assign n12680 = n272 & n8440 ;
  assign n12681 = n12679 | n12680 ;
  assign n12682 = n12681 ^ x56 ^ 1'b0 ;
  assign n12683 = ( n12575 & ~n12672 ) | ( n12575 & n12682 ) | ( ~n12672 & n12682 ) ;
  assign n12684 = n12682 ^ n12672 ^ n12575 ;
  assign n12685 = x108 & n408 ;
  assign n12686 = ( x110 & n403 ) | ( x110 & n12685 ) | ( n403 & n12685 ) ;
  assign n12687 = n12685 | n12686 ;
  assign n12688 = x109 & ~n410 ;
  assign n12689 = ( x109 & n12687 ) | ( x109 & ~n12688 ) | ( n12687 & ~n12688 ) ;
  assign n12690 = n402 & n8820 ;
  assign n12691 = n12689 | n12690 ;
  assign n12692 = n12691 ^ x53 ^ 1'b0 ;
  assign n12693 = n12692 ^ n12684 ^ n12584 ;
  assign n12694 = ( n12584 & ~n12684 ) | ( n12584 & n12692 ) | ( ~n12684 & n12692 ) ;
  assign n12695 = x111 & n561 ;
  assign n12696 = ( x113 & n551 ) | ( x113 & n12695 ) | ( n551 & n12695 ) ;
  assign n12697 = n12695 | n12696 ;
  assign n12698 = x112 & ~n550 ;
  assign n12699 = ( x112 & n12697 ) | ( x112 & ~n12698 ) | ( n12697 & ~n12698 ) ;
  assign n12700 = n553 & n9199 ;
  assign n12701 = n12699 | n12700 ;
  assign n12702 = n12701 ^ x50 ^ 1'b0 ;
  assign n12703 = n12702 ^ n12693 ^ n12595 ;
  assign n12704 = ( n12595 & ~n12693 ) | ( n12595 & n12702 ) | ( ~n12693 & n12702 ) ;
  assign n12705 = x114 & n744 ;
  assign n12706 = ( x116 & n730 ) | ( x116 & n12705 ) | ( n730 & n12705 ) ;
  assign n12707 = n12705 | n12706 ;
  assign n12708 = x115 & ~n732 ;
  assign n12709 = ( x115 & n12707 ) | ( x115 & ~n12708 ) | ( n12707 & ~n12708 ) ;
  assign n12710 = n731 & n9513 ;
  assign n12711 = n12709 | n12710 ;
  assign n12712 = n12711 ^ x47 ^ 1'b0 ;
  assign n12713 = ( n12606 & ~n12703 ) | ( n12606 & n12712 ) | ( ~n12703 & n12712 ) ;
  assign n12714 = n12712 ^ n12703 ^ n12606 ;
  assign n12715 = x117 & n888 ;
  assign n12716 = ( x119 & n878 ) | ( x119 & n12715 ) | ( n878 & n12715 ) ;
  assign n12717 = n12715 | n12716 ;
  assign n12718 = x118 & ~n877 ;
  assign n12719 = ( x118 & n12717 ) | ( x118 & ~n12718 ) | ( n12717 & ~n12718 ) ;
  assign n12720 = n880 & n9733 ;
  assign n12721 = n12719 | n12720 ;
  assign n12722 = n12721 ^ x44 ^ 1'b0 ;
  assign n12723 = n12722 ^ n12714 ^ n12616 ;
  assign n12724 = ( n12616 & ~n12714 ) | ( n12616 & n12722 ) | ( ~n12714 & n12722 ) ;
  assign n12725 = x101 & n208 ;
  assign n12726 = ( x103 & n194 ) | ( x103 & n12725 ) | ( n194 & n12725 ) ;
  assign n12727 = n12725 | n12726 ;
  assign n12728 = x102 & ~n192 ;
  assign n12729 = ( x102 & n12727 ) | ( x102 & ~n12728 ) | ( n12727 & ~n12728 ) ;
  assign n12730 = x120 & n1058 ;
  assign n12731 = n12673 | n12729 ;
  assign n12732 = ( x122 & n1065 ) | ( x122 & n12730 ) | ( n1065 & n12730 ) ;
  assign n12733 = n12730 | n12732 ;
  assign n12734 = x121 & ~n1060 ;
  assign n12735 = ( x121 & n12733 ) | ( x121 & ~n12734 ) | ( n12733 & ~n12734 ) ;
  assign n12736 = n1063 & n9806 ;
  assign n12737 = n12735 | n12736 ;
  assign n12738 = n12737 ^ x41 ^ 1'b0 ;
  assign n12739 = n12738 ^ n12723 ^ n12626 ;
  assign n12740 = ( n12626 & ~n12723 ) | ( n12626 & n12738 ) | ( ~n12723 & n12738 ) ;
  assign n12741 = x123 & n2156 ;
  assign n12742 = ( x125 & n2163 ) | ( x125 & n12741 ) | ( n2163 & n12741 ) ;
  assign n12743 = n12741 | n12742 ;
  assign n12744 = x124 & ~n2158 ;
  assign n12745 = ( x124 & n12743 ) | ( x124 & ~n12744 ) | ( n12743 & ~n12744 ) ;
  assign n12746 = n2161 & n9883 ;
  assign n12747 = n12745 | n12746 ;
  assign n12748 = n12747 ^ x38 ^ 1'b0 ;
  assign n12749 = n12748 ^ n12739 ^ n12636 ;
  assign n12750 = ( n12636 & ~n12739 ) | ( n12636 & n12748 ) | ( ~n12739 & n12748 ) ;
  assign n12751 = x124 & n2156 ;
  assign n12752 = ( x126 & n2163 ) | ( x126 & n12751 ) | ( n2163 & n12751 ) ;
  assign n12753 = n12751 | n12752 ;
  assign n12754 = n12546 ^ x35 ^ 1'b0 ;
  assign n12755 = x125 & n2156 ;
  assign n12756 = ( x127 & n2163 ) | ( x127 & n12755 ) | ( n2163 & n12755 ) ;
  assign n12757 = n12755 | n12756 ;
  assign n12758 = x126 & ~n2158 ;
  assign n12759 = ( x126 & n12757 ) | ( x126 & ~n12758 ) | ( n12757 & ~n12758 ) ;
  assign n12760 = x125 & ~n2158 ;
  assign n12761 = ( x125 & n12753 ) | ( x125 & ~n12760 ) | ( n12753 & ~n12760 ) ;
  assign n12762 = n12754 ^ n12749 ^ n12645 ;
  assign n12763 = ( n12645 & ~n12749 ) | ( n12645 & n12754 ) | ( ~n12749 & n12754 ) ;
  assign n12764 = n2161 & n9949 ;
  assign n12765 = n12759 | n12764 ;
  assign n12766 = x100 & n208 ;
  assign n12767 = ( x102 & n194 ) | ( x102 & n12766 ) | ( n194 & n12766 ) ;
  assign n12768 = n12559 ^ x35 ^ 1'b0 ;
  assign n12769 = n12766 | n12767 ;
  assign n12770 = x127 & ~n2158 ;
  assign n12771 = x101 & ~n192 ;
  assign n12772 = ( x101 & n12769 ) | ( x101 & ~n12771 ) | ( n12769 & ~n12771 ) ;
  assign n12773 = x126 & n2156 ;
  assign n12774 = ( x127 & ~n12770 ) | ( x127 & n12773 ) | ( ~n12770 & n12773 ) ;
  assign n12775 = ( n2161 & n9958 ) | ( n2161 & n12773 ) | ( n9958 & n12773 ) ;
  assign n12776 = n12774 | n12775 ;
  assign n12777 = n197 & n5947 ;
  assign n12778 = x127 & n2156 ;
  assign n12779 = ( n2161 & n9968 ) | ( n2161 & n12778 ) | ( n9968 & n12778 ) ;
  assign n12780 = n2161 & n9917 ;
  assign n12781 = n12772 | n12777 ;
  assign n12782 = n12761 | n12780 ;
  assign n12783 = n12781 ^ x62 ^ 1'b0 ;
  assign n12784 = n12762 ^ n12650 ^ n12648 ;
  assign n12785 = n12778 | n12779 ;
  assign n12786 = ( ~n12648 & n12650 ) | ( ~n12648 & n12762 ) | ( n12650 & n12762 ) ;
  assign n12787 = x103 & n133 ;
  assign n12788 = x98 & n325 ;
  assign n12789 = x99 & ~n242 ;
  assign n12790 = ( x99 & n12788 ) | ( x99 & ~n12789 ) | ( n12788 & ~n12789 ) ;
  assign n12791 = ( x105 & n142 ) | ( x105 & n12787 ) | ( n142 & n12787 ) ;
  assign n12792 = n12787 | n12791 ;
  assign n12793 = x104 & ~n134 ;
  assign n12794 = ( x104 & n12792 ) | ( x104 & ~n12793 ) | ( n12792 & ~n12793 ) ;
  assign n12795 = ( n12663 & n12666 ) | ( n12663 & ~n12790 ) | ( n12666 & ~n12790 ) ;
  assign n12796 = n12790 ^ n12666 ^ n12663 ;
  assign n12797 = n140 & n8105 ;
  assign n12798 = n12794 | n12797 ;
  assign n12799 = n12798 ^ x59 ^ 1'b0 ;
  assign n12800 = n12799 ^ n12796 ^ n12783 ;
  assign n12801 = ( n12783 & ~n12796 ) | ( n12783 & n12799 ) | ( ~n12796 & n12799 ) ;
  assign n12802 = x106 & n263 ;
  assign n12803 = ( x108 & n264 ) | ( x108 & n12802 ) | ( n264 & n12802 ) ;
  assign n12804 = n12802 | n12803 ;
  assign n12805 = x107 & ~n260 ;
  assign n12806 = ( x107 & n12804 ) | ( x107 & ~n12805 ) | ( n12804 & ~n12805 ) ;
  assign n12807 = n272 & n8557 ;
  assign n12808 = n12806 | n12807 ;
  assign n12809 = n12808 ^ x56 ^ 1'b0 ;
  assign n12810 = ( n12674 & ~n12800 ) | ( n12674 & n12809 ) | ( ~n12800 & n12809 ) ;
  assign n12811 = n12809 ^ n12800 ^ n12674 ;
  assign n12812 = x109 & n408 ;
  assign n12813 = ( x111 & n403 ) | ( x111 & n12812 ) | ( n403 & n12812 ) ;
  assign n12814 = n12812 | n12813 ;
  assign n12815 = x110 & ~n410 ;
  assign n12816 = ( x110 & n12814 ) | ( x110 & ~n12815 ) | ( n12814 & ~n12815 ) ;
  assign n12817 = n402 & n8946 ;
  assign n12818 = n12816 | n12817 ;
  assign n12819 = n12818 ^ x53 ^ 1'b0 ;
  assign n12820 = n12819 ^ n12811 ^ n12683 ;
  assign n12821 = ( n12683 & ~n12811 ) | ( n12683 & n12819 ) | ( ~n12811 & n12819 ) ;
  assign n12822 = x112 & n561 ;
  assign n12823 = ( x114 & n551 ) | ( x114 & n12822 ) | ( n551 & n12822 ) ;
  assign n12824 = n12822 | n12823 ;
  assign n12825 = x113 & ~n550 ;
  assign n12826 = ( x113 & n12824 ) | ( x113 & ~n12825 ) | ( n12824 & ~n12825 ) ;
  assign n12827 = n553 & n9279 ;
  assign n12828 = n12826 | n12827 ;
  assign n12829 = n12828 ^ x50 ^ 1'b0 ;
  assign n12830 = ( n12694 & ~n12820 ) | ( n12694 & n12829 ) | ( ~n12820 & n12829 ) ;
  assign n12831 = n12829 ^ n12820 ^ n12694 ;
  assign n12832 = x115 & n744 ;
  assign n12833 = ( x117 & n730 ) | ( x117 & n12832 ) | ( n730 & n12832 ) ;
  assign n12834 = n12832 | n12833 ;
  assign n12835 = x116 & ~n732 ;
  assign n12836 = ( x116 & n12834 ) | ( x116 & ~n12835 ) | ( n12834 & ~n12835 ) ;
  assign n12837 = n731 & n9569 ;
  assign n12838 = n12836 | n12837 ;
  assign n12839 = n12838 ^ x47 ^ 1'b0 ;
  assign n12840 = ( n12704 & ~n12831 ) | ( n12704 & n12839 ) | ( ~n12831 & n12839 ) ;
  assign n12841 = n12839 ^ n12831 ^ n12704 ;
  assign n12842 = x118 & n888 ;
  assign n12843 = ( x120 & n878 ) | ( x120 & n12842 ) | ( n878 & n12842 ) ;
  assign n12844 = n12842 | n12843 ;
  assign n12845 = x119 & ~n877 ;
  assign n12846 = ( x119 & n12844 ) | ( x119 & ~n12845 ) | ( n12844 & ~n12845 ) ;
  assign n12847 = n880 & n9756 ;
  assign n12848 = n12846 | n12847 ;
  assign n12849 = n12848 ^ x44 ^ 1'b0 ;
  assign n12850 = n12849 ^ n12841 ^ n12713 ;
  assign n12851 = ( n12713 & ~n12841 ) | ( n12713 & n12849 ) | ( ~n12841 & n12849 ) ;
  assign n12852 = x121 & n1058 ;
  assign n12853 = ( x123 & n1065 ) | ( x123 & n12852 ) | ( n1065 & n12852 ) ;
  assign n12854 = n12852 | n12853 ;
  assign n12855 = x122 & ~n1060 ;
  assign n12856 = ( x122 & n12854 ) | ( x122 & ~n12855 ) | ( n12854 & ~n12855 ) ;
  assign n12857 = n1063 & n9828 ;
  assign n12858 = n12856 | n12857 ;
  assign n12859 = n12731 ^ x62 ^ 1'b0 ;
  assign n12860 = n12782 ^ x38 ^ 1'b0 ;
  assign n12861 = n12858 ^ x41 ^ 1'b0 ;
  assign n12862 = ( n12724 & ~n12850 ) | ( n12724 & n12861 ) | ( ~n12850 & n12861 ) ;
  assign n12863 = n12861 ^ n12850 ^ n12724 ;
  assign n12864 = x104 & n133 ;
  assign n12865 = n12863 ^ n12860 ^ n12740 ;
  assign n12866 = ( n12740 & n12860 ) | ( n12740 & ~n12863 ) | ( n12860 & ~n12863 ) ;
  assign n12867 = ( n12750 & n12768 ) | ( n12750 & ~n12865 ) | ( n12768 & ~n12865 ) ;
  assign n12868 = x105 & ~n134 ;
  assign n12869 = n12865 ^ n12768 ^ n12750 ;
  assign n12870 = x113 & n561 ;
  assign n12871 = ( x106 & n142 ) | ( x106 & n12864 ) | ( n142 & n12864 ) ;
  assign n12872 = n12864 | n12871 ;
  assign n12873 = ( x115 & n551 ) | ( x115 & n12870 ) | ( n551 & n12870 ) ;
  assign n12874 = ( x105 & ~n12868 ) | ( x105 & n12872 ) | ( ~n12868 & n12872 ) ;
  assign n12875 = x110 & n408 ;
  assign n12876 = n12870 | n12873 ;
  assign n12877 = x114 & ~n550 ;
  assign n12878 = ( x114 & n12876 ) | ( x114 & ~n12877 ) | ( n12876 & ~n12877 ) ;
  assign n12879 = ( x112 & n403 ) | ( x112 & n12875 ) | ( n403 & n12875 ) ;
  assign n12880 = n12875 | n12879 ;
  assign n12881 = n140 & n8287 ;
  assign n12882 = n12874 | n12881 ;
  assign n12883 = x111 & ~n410 ;
  assign n12884 = ( x111 & n12880 ) | ( x111 & ~n12883 ) | ( n12880 & ~n12883 ) ;
  assign n12885 = ( ~n12763 & n12786 ) | ( ~n12763 & n12869 ) | ( n12786 & n12869 ) ;
  assign n12886 = n12869 ^ n12786 ^ n12763 ;
  assign n12887 = x99 & n325 ;
  assign n12888 = x100 & ~n242 ;
  assign n12889 = ( x100 & n12887 ) | ( x100 & ~n12888 ) | ( n12887 & ~n12888 ) ;
  assign n12890 = n12889 ^ n12790 ^ x35 ;
  assign n12891 = ( ~x35 & n12790 ) | ( ~x35 & n12889 ) | ( n12790 & n12889 ) ;
  assign n12892 = n402 & n9080 ;
  assign n12893 = n12884 | n12892 ;
  assign n12894 = n553 & n9414 ;
  assign n12895 = n12882 ^ x59 ^ 1'b0 ;
  assign n12896 = n12878 | n12894 ;
  assign n12897 = n12890 ^ n12859 ^ n12795 ;
  assign n12898 = n12896 ^ x50 ^ 1'b0 ;
  assign n12899 = n12893 ^ x53 ^ 1'b0 ;
  assign n12900 = ( n12795 & n12859 ) | ( n12795 & ~n12890 ) | ( n12859 & ~n12890 ) ;
  assign n12901 = x107 & n263 ;
  assign n12902 = n12897 ^ n12895 ^ n12801 ;
  assign n12903 = ( n12801 & n12895 ) | ( n12801 & ~n12897 ) | ( n12895 & ~n12897 ) ;
  assign n12904 = x108 & ~n260 ;
  assign n12905 = ( x109 & n264 ) | ( x109 & n12901 ) | ( n264 & n12901 ) ;
  assign n12906 = n12901 | n12905 ;
  assign n12907 = ( x108 & ~n12904 ) | ( x108 & n12906 ) | ( ~n12904 & n12906 ) ;
  assign n12908 = n272 & n8680 ;
  assign n12909 = n12907 | n12908 ;
  assign n12910 = n12909 ^ x56 ^ 1'b0 ;
  assign n12911 = n12910 ^ n12902 ^ n12810 ;
  assign n12912 = n12911 ^ n12899 ^ n12821 ;
  assign n12913 = ( n12810 & ~n12902 ) | ( n12810 & n12910 ) | ( ~n12902 & n12910 ) ;
  assign n12914 = ( n12821 & n12899 ) | ( n12821 & ~n12911 ) | ( n12899 & ~n12911 ) ;
  assign n12915 = n12912 ^ n12898 ^ n12830 ;
  assign n12916 = ( n12830 & n12898 ) | ( n12830 & ~n12912 ) | ( n12898 & ~n12912 ) ;
  assign n12917 = n12765 ^ x38 ^ 1'b0 ;
  assign n12918 = x116 & n744 ;
  assign n12919 = n12776 ^ x38 ^ 1'b0 ;
  assign n12920 = ( x118 & n730 ) | ( x118 & n12918 ) | ( n730 & n12918 ) ;
  assign n12921 = n12918 | n12920 ;
  assign n12922 = x117 & ~n732 ;
  assign n12923 = ( x117 & n12921 ) | ( x117 & ~n12922 ) | ( n12921 & ~n12922 ) ;
  assign n12924 = n731 & n9671 ;
  assign n12925 = n12923 | n12924 ;
  assign n12926 = n12925 ^ x47 ^ 1'b0 ;
  assign n12927 = n12926 ^ n12915 ^ n12840 ;
  assign n12928 = ( n12840 & ~n12915 ) | ( n12840 & n12926 ) | ( ~n12915 & n12926 ) ;
  assign n12929 = x119 & n888 ;
  assign n12930 = ( x121 & n878 ) | ( x121 & n12929 ) | ( n878 & n12929 ) ;
  assign n12931 = n12929 | n12930 ;
  assign n12932 = x120 & ~n877 ;
  assign n12933 = ( x120 & n12931 ) | ( x120 & ~n12932 ) | ( n12931 & ~n12932 ) ;
  assign n12934 = n197 & n8012 ;
  assign n12935 = n880 & n9808 ;
  assign n12936 = n12933 | n12935 ;
  assign n12937 = n12936 ^ x44 ^ 1'b0 ;
  assign n12938 = n12937 ^ n12927 ^ n12851 ;
  assign n12939 = ( n12851 & ~n12927 ) | ( n12851 & n12937 ) | ( ~n12927 & n12937 ) ;
  assign n12940 = x122 & n1058 ;
  assign n12941 = ( x124 & n1065 ) | ( x124 & n12940 ) | ( n1065 & n12940 ) ;
  assign n12942 = n12940 | n12941 ;
  assign n12943 = x123 & ~n1060 ;
  assign n12944 = ( x123 & n12942 ) | ( x123 & ~n12943 ) | ( n12942 & ~n12943 ) ;
  assign n12945 = n1063 & n9858 ;
  assign n12946 = n12944 | n12945 ;
  assign n12947 = n12946 ^ x41 ^ 1'b0 ;
  assign n12948 = ( n12862 & ~n12938 ) | ( n12862 & n12947 ) | ( ~n12938 & n12947 ) ;
  assign n12949 = n12947 ^ n12938 ^ n12862 ;
  assign n12950 = n12949 ^ n12917 ^ n12866 ;
  assign n12951 = ( ~n12867 & n12885 ) | ( ~n12867 & n12950 ) | ( n12885 & n12950 ) ;
  assign n12952 = n12950 ^ n12885 ^ n12867 ;
  assign n12953 = x105 & n133 ;
  assign n12954 = ( x107 & n142 ) | ( x107 & n12953 ) | ( n142 & n12953 ) ;
  assign n12955 = n12953 | n12954 ;
  assign n12956 = x106 & ~n134 ;
  assign n12957 = ( x106 & n12955 ) | ( x106 & ~n12956 ) | ( n12955 & ~n12956 ) ;
  assign n12958 = n140 & n8440 ;
  assign n12959 = n12957 | n12958 ;
  assign n12960 = x102 & n208 ;
  assign n12961 = n12959 ^ x59 ^ 1'b0 ;
  assign n12962 = ( n12866 & n12917 ) | ( n12866 & ~n12949 ) | ( n12917 & ~n12949 ) ;
  assign n12963 = x101 & ~n242 ;
  assign n12964 = x100 & n325 ;
  assign n12965 = n197 & n8105 ;
  assign n12966 = ( x101 & ~n12963 ) | ( x101 & n12964 ) | ( ~n12963 & n12964 ) ;
  assign n12967 = ( x104 & n194 ) | ( x104 & n12960 ) | ( n194 & n12960 ) ;
  assign n12968 = n12960 | n12967 ;
  assign n12969 = x103 & ~n192 ;
  assign n12970 = ( x103 & n12968 ) | ( x103 & ~n12969 ) | ( n12968 & ~n12969 ) ;
  assign n12971 = n12934 | n12970 ;
  assign n12972 = n12971 ^ x62 ^ 1'b0 ;
  assign n12973 = ( n12891 & ~n12966 ) | ( n12891 & n12972 ) | ( ~n12966 & n12972 ) ;
  assign n12974 = n12972 ^ n12966 ^ n12891 ;
  assign n12975 = ( n12900 & n12961 ) | ( n12900 & ~n12974 ) | ( n12961 & ~n12974 ) ;
  assign n12976 = n12974 ^ n12961 ^ n12900 ;
  assign n12977 = x108 & n263 ;
  assign n12978 = ( x110 & n264 ) | ( x110 & n12977 ) | ( n264 & n12977 ) ;
  assign n12979 = n12977 | n12978 ;
  assign n12980 = x109 & ~n260 ;
  assign n12981 = ( x109 & n12979 ) | ( x109 & ~n12980 ) | ( n12979 & ~n12980 ) ;
  assign n12982 = n272 & n8820 ;
  assign n12983 = n12981 | n12982 ;
  assign n12984 = n12983 ^ x56 ^ 1'b0 ;
  assign n12985 = ( n12903 & ~n12976 ) | ( n12903 & n12984 ) | ( ~n12976 & n12984 ) ;
  assign n12986 = n12984 ^ n12976 ^ n12903 ;
  assign n12987 = x111 & n408 ;
  assign n12988 = ( x113 & n403 ) | ( x113 & n12987 ) | ( n403 & n12987 ) ;
  assign n12989 = n12987 | n12988 ;
  assign n12990 = x112 & ~n410 ;
  assign n12991 = ( x112 & n12989 ) | ( x112 & ~n12990 ) | ( n12989 & ~n12990 ) ;
  assign n12992 = n402 & n9199 ;
  assign n12993 = n12991 | n12992 ;
  assign n12994 = n12993 ^ x53 ^ 1'b0 ;
  assign n12995 = ( n12913 & ~n12986 ) | ( n12913 & n12994 ) | ( ~n12986 & n12994 ) ;
  assign n12996 = n12994 ^ n12986 ^ n12913 ;
  assign n12997 = x114 & n561 ;
  assign n12998 = ( x116 & n551 ) | ( x116 & n12997 ) | ( n551 & n12997 ) ;
  assign n12999 = n12997 | n12998 ;
  assign n13000 = x115 & ~n550 ;
  assign n13001 = ( x115 & n12999 ) | ( x115 & ~n13000 ) | ( n12999 & ~n13000 ) ;
  assign n13002 = n553 & n9513 ;
  assign n13003 = n13001 | n13002 ;
  assign n13004 = n13003 ^ x50 ^ 1'b0 ;
  assign n13005 = n13004 ^ n12996 ^ n12914 ;
  assign n13006 = ( n12914 & ~n12996 ) | ( n12914 & n13004 ) | ( ~n12996 & n13004 ) ;
  assign n13007 = x117 & n744 ;
  assign n13008 = ( x119 & n730 ) | ( x119 & n13007 ) | ( n730 & n13007 ) ;
  assign n13009 = n13007 | n13008 ;
  assign n13010 = x118 & ~n732 ;
  assign n13011 = ( x118 & n13009 ) | ( x118 & ~n13010 ) | ( n13009 & ~n13010 ) ;
  assign n13012 = n731 & n9733 ;
  assign n13013 = n13011 | n13012 ;
  assign n13014 = n13013 ^ x47 ^ 1'b0 ;
  assign n13015 = ( n12916 & ~n13005 ) | ( n12916 & n13014 ) | ( ~n13005 & n13014 ) ;
  assign n13016 = n13014 ^ n13005 ^ n12916 ;
  assign n13017 = x120 & n888 ;
  assign n13018 = ( x122 & n878 ) | ( x122 & n13017 ) | ( n878 & n13017 ) ;
  assign n13019 = n13017 | n13018 ;
  assign n13020 = x121 & ~n877 ;
  assign n13021 = ( x121 & n13019 ) | ( x121 & ~n13020 ) | ( n13019 & ~n13020 ) ;
  assign n13022 = n880 & n9806 ;
  assign n13023 = n13021 | n13022 ;
  assign n13024 = n13023 ^ x44 ^ 1'b0 ;
  assign n13025 = ( n12928 & ~n13016 ) | ( n12928 & n13024 ) | ( ~n13016 & n13024 ) ;
  assign n13026 = n13024 ^ n13016 ^ n12928 ;
  assign n13027 = x123 & n1058 ;
  assign n13028 = ( x125 & n1065 ) | ( x125 & n13027 ) | ( n1065 & n13027 ) ;
  assign n13029 = n13027 | n13028 ;
  assign n13030 = x124 & ~n1060 ;
  assign n13031 = ( x124 & n13029 ) | ( x124 & ~n13030 ) | ( n13029 & ~n13030 ) ;
  assign n13032 = n1063 & n9883 ;
  assign n13033 = n13031 | n13032 ;
  assign n13034 = n13033 ^ x41 ^ 1'b0 ;
  assign n13035 = ( n12939 & ~n13026 ) | ( n12939 & n13034 ) | ( ~n13026 & n13034 ) ;
  assign n13036 = n13034 ^ n13026 ^ n12939 ;
  assign n13037 = ( n12919 & n12948 ) | ( n12919 & ~n13036 ) | ( n12948 & ~n13036 ) ;
  assign n13038 = n13036 ^ n12948 ^ n12919 ;
  assign n13039 = n13038 ^ n12962 ^ n12951 ;
  assign n13040 = ( n12951 & ~n12962 ) | ( n12951 & n13038 ) | ( ~n12962 & n13038 ) ;
  assign n13041 = x104 & ~n192 ;
  assign n13042 = x103 & n208 ;
  assign n13043 = ( x105 & n194 ) | ( x105 & n13042 ) | ( n194 & n13042 ) ;
  assign n13044 = n13042 | n13043 ;
  assign n13045 = ( x104 & ~n13041 ) | ( x104 & n13044 ) | ( ~n13041 & n13044 ) ;
  assign n13046 = n12785 ^ x38 ^ 1'b0 ;
  assign n13047 = x125 & n1058 ;
  assign n13048 = x124 & n1058 ;
  assign n13049 = n12965 | n13045 ;
  assign n13050 = ( x127 & n1065 ) | ( x127 & n13047 ) | ( n1065 & n13047 ) ;
  assign n13051 = ( x126 & n1065 ) | ( x126 & n13048 ) | ( n1065 & n13048 ) ;
  assign n13052 = n13048 | n13051 ;
  assign n13053 = n1063 & n9917 ;
  assign n13054 = n13047 | n13050 ;
  assign n13055 = x125 & ~n1060 ;
  assign n13056 = ( x125 & n13052 ) | ( x125 & ~n13055 ) | ( n13052 & ~n13055 ) ;
  assign n13057 = x106 & n133 ;
  assign n13058 = n13053 | n13056 ;
  assign n13059 = ( x108 & n142 ) | ( x108 & n13057 ) | ( n142 & n13057 ) ;
  assign n13060 = n13057 | n13059 ;
  assign n13061 = x107 & ~n134 ;
  assign n13062 = ( x107 & n13060 ) | ( x107 & ~n13061 ) | ( n13060 & ~n13061 ) ;
  assign n13063 = x126 & ~n1060 ;
  assign n13064 = ( x126 & n13054 ) | ( x126 & ~n13063 ) | ( n13054 & ~n13063 ) ;
  assign n13065 = n1063 & n9949 ;
  assign n13066 = n13064 | n13065 ;
  assign n13067 = n140 & n8557 ;
  assign n13068 = n13062 | n13067 ;
  assign n13069 = n13058 ^ x41 ^ 1'b0 ;
  assign n13070 = n13049 ^ x62 ^ 1'b0 ;
  assign n13071 = x127 & n1058 ;
  assign n13072 = n13068 ^ x59 ^ 1'b0 ;
  assign n13073 = x127 & ~n1060 ;
  assign n13074 = x126 & n1058 ;
  assign n13075 = ( x127 & ~n13073 ) | ( x127 & n13074 ) | ( ~n13073 & n13074 ) ;
  assign n13076 = ( n1063 & n9958 ) | ( n1063 & n13074 ) | ( n9958 & n13074 ) ;
  assign n13077 = ( n1063 & n9968 ) | ( n1063 & n13071 ) | ( n9968 & n13071 ) ;
  assign n13078 = n13071 | n13077 ;
  assign n13079 = x101 & n325 ;
  assign n13080 = n13075 | n13076 ;
  assign n13081 = x102 & ~n242 ;
  assign n13082 = ( x102 & n13079 ) | ( x102 & ~n13081 ) | ( n13079 & ~n13081 ) ;
  assign n13083 = n13082 ^ n12973 ^ n12966 ;
  assign n13084 = ( ~n12966 & n12973 ) | ( ~n12966 & n13082 ) | ( n12973 & n13082 ) ;
  assign n13085 = ( n13070 & n13072 ) | ( n13070 & ~n13083 ) | ( n13072 & ~n13083 ) ;
  assign n13086 = n13083 ^ n13072 ^ n13070 ;
  assign n13087 = x109 & n263 ;
  assign n13088 = ( x111 & n264 ) | ( x111 & n13087 ) | ( n264 & n13087 ) ;
  assign n13089 = n13087 | n13088 ;
  assign n13090 = x110 & ~n260 ;
  assign n13091 = ( x110 & n13089 ) | ( x110 & ~n13090 ) | ( n13089 & ~n13090 ) ;
  assign n13092 = n272 & n8946 ;
  assign n13093 = n13091 | n13092 ;
  assign n13094 = n13093 ^ x56 ^ 1'b0 ;
  assign n13095 = ( n12975 & ~n13086 ) | ( n12975 & n13094 ) | ( ~n13086 & n13094 ) ;
  assign n13096 = n13094 ^ n13086 ^ n12975 ;
  assign n13097 = x112 & n408 ;
  assign n13098 = ( x114 & n403 ) | ( x114 & n13097 ) | ( n403 & n13097 ) ;
  assign n13099 = n13097 | n13098 ;
  assign n13100 = x113 & ~n410 ;
  assign n13101 = ( x113 & n13099 ) | ( x113 & ~n13100 ) | ( n13099 & ~n13100 ) ;
  assign n13102 = n402 & n9279 ;
  assign n13103 = n13101 | n13102 ;
  assign n13104 = n13103 ^ x53 ^ 1'b0 ;
  assign n13105 = ( n12985 & ~n13096 ) | ( n12985 & n13104 ) | ( ~n13096 & n13104 ) ;
  assign n13106 = n13104 ^ n13096 ^ n12985 ;
  assign n13107 = x115 & n561 ;
  assign n13108 = ( x117 & n551 ) | ( x117 & n13107 ) | ( n551 & n13107 ) ;
  assign n13109 = n13107 | n13108 ;
  assign n13110 = x116 & ~n550 ;
  assign n13111 = ( x116 & n13109 ) | ( x116 & ~n13110 ) | ( n13109 & ~n13110 ) ;
  assign n13112 = n553 & n9569 ;
  assign n13113 = n13111 | n13112 ;
  assign n13114 = n13113 ^ x50 ^ 1'b0 ;
  assign n13115 = ( n12995 & ~n13106 ) | ( n12995 & n13114 ) | ( ~n13106 & n13114 ) ;
  assign n13116 = n13114 ^ n13106 ^ n12995 ;
  assign n13117 = x118 & n744 ;
  assign n13118 = ( x120 & n730 ) | ( x120 & n13117 ) | ( n730 & n13117 ) ;
  assign n13119 = n13117 | n13118 ;
  assign n13120 = x119 & ~n732 ;
  assign n13121 = ( x119 & n13119 ) | ( x119 & ~n13120 ) | ( n13119 & ~n13120 ) ;
  assign n13122 = n731 & n9756 ;
  assign n13123 = n13121 | n13122 ;
  assign n13124 = n13123 ^ x47 ^ 1'b0 ;
  assign n13125 = ( n13006 & ~n13116 ) | ( n13006 & n13124 ) | ( ~n13116 & n13124 ) ;
  assign n13126 = n13124 ^ n13116 ^ n13006 ;
  assign n13127 = x121 & n888 ;
  assign n13128 = ( x123 & n878 ) | ( x123 & n13127 ) | ( n878 & n13127 ) ;
  assign n13129 = n13127 | n13128 ;
  assign n13130 = x122 & ~n877 ;
  assign n13131 = ( x122 & n13129 ) | ( x122 & ~n13130 ) | ( n13129 & ~n13130 ) ;
  assign n13132 = n880 & n9828 ;
  assign n13133 = n13131 | n13132 ;
  assign n13134 = n13133 ^ x44 ^ 1'b0 ;
  assign n13135 = ( n13015 & ~n13126 ) | ( n13015 & n13134 ) | ( ~n13126 & n13134 ) ;
  assign n13136 = n13134 ^ n13126 ^ n13015 ;
  assign n13137 = ( n13025 & n13069 ) | ( n13025 & ~n13136 ) | ( n13069 & ~n13136 ) ;
  assign n13138 = n13136 ^ n13069 ^ n13025 ;
  assign n13139 = n13138 ^ n13046 ^ n13035 ;
  assign n13140 = n13139 ^ n13040 ^ n13037 ;
  assign n13141 = ( n13035 & n13046 ) | ( n13035 & ~n13138 ) | ( n13046 & ~n13138 ) ;
  assign n13142 = ( ~n13037 & n13040 ) | ( ~n13037 & n13139 ) | ( n13040 & n13139 ) ;
  assign n13143 = x104 & n208 ;
  assign n13144 = ( x106 & n194 ) | ( x106 & n13143 ) | ( n194 & n13143 ) ;
  assign n13145 = n13143 | n13144 ;
  assign n13146 = x105 & ~n192 ;
  assign n13147 = ( x105 & n13145 ) | ( x105 & ~n13146 ) | ( n13145 & ~n13146 ) ;
  assign n13148 = n197 & n8287 ;
  assign n13149 = n13147 | n13148 ;
  assign n13150 = x103 & ~n242 ;
  assign n13151 = x102 & n325 ;
  assign n13152 = ( x103 & ~n13150 ) | ( x103 & n13151 ) | ( ~n13150 & n13151 ) ;
  assign n13153 = ( ~x38 & n12966 ) | ( ~x38 & n13152 ) | ( n12966 & n13152 ) ;
  assign n13154 = n13152 ^ n12966 ^ x38 ;
  assign n13155 = n13149 ^ x62 ^ 1'b0 ;
  assign n13156 = n13155 ^ n13154 ^ n13084 ;
  assign n13157 = ( n13084 & ~n13154 ) | ( n13084 & n13155 ) | ( ~n13154 & n13155 ) ;
  assign n13158 = x105 & n208 ;
  assign n13159 = ( x107 & n194 ) | ( x107 & n13158 ) | ( n194 & n13158 ) ;
  assign n13160 = n13158 | n13159 ;
  assign n13161 = x106 & ~n192 ;
  assign n13162 = ( x106 & n13160 ) | ( x106 & ~n13161 ) | ( n13160 & ~n13161 ) ;
  assign n13163 = ( n197 & n8440 ) | ( n197 & n13162 ) | ( n8440 & n13162 ) ;
  assign n13164 = n13162 | n13163 ;
  assign n13165 = x107 & n133 ;
  assign n13166 = ( x109 & n142 ) | ( x109 & n13165 ) | ( n142 & n13165 ) ;
  assign n13167 = n13165 | n13166 ;
  assign n13168 = x108 & ~n134 ;
  assign n13169 = ( x108 & n13167 ) | ( x108 & ~n13168 ) | ( n13167 & ~n13168 ) ;
  assign n13170 = n140 & n8680 ;
  assign n13171 = n13169 | n13170 ;
  assign n13172 = n13164 ^ x62 ^ 1'b0 ;
  assign n13173 = n13171 ^ x59 ^ 1'b0 ;
  assign n13174 = ( n13085 & ~n13156 ) | ( n13085 & n13173 ) | ( ~n13156 & n13173 ) ;
  assign n13175 = n13173 ^ n13156 ^ n13085 ;
  assign n13176 = x110 & n263 ;
  assign n13177 = n13080 ^ x41 ^ 1'b0 ;
  assign n13178 = n13066 ^ x41 ^ 1'b0 ;
  assign n13179 = ( x112 & n264 ) | ( x112 & n13176 ) | ( n264 & n13176 ) ;
  assign n13180 = n13176 | n13179 ;
  assign n13181 = x111 & ~n260 ;
  assign n13182 = ( x111 & n13180 ) | ( x111 & ~n13181 ) | ( n13180 & ~n13181 ) ;
  assign n13183 = n272 & n9080 ;
  assign n13184 = n13182 | n13183 ;
  assign n13185 = n13184 ^ x56 ^ 1'b0 ;
  assign n13186 = n13185 ^ n13175 ^ n13095 ;
  assign n13187 = ( n13095 & ~n13175 ) | ( n13095 & n13185 ) | ( ~n13175 & n13185 ) ;
  assign n13188 = x113 & n408 ;
  assign n13189 = ( x115 & n403 ) | ( x115 & n13188 ) | ( n403 & n13188 ) ;
  assign n13190 = n13188 | n13189 ;
  assign n13191 = x114 & ~n410 ;
  assign n13192 = ( x114 & n13190 ) | ( x114 & ~n13191 ) | ( n13190 & ~n13191 ) ;
  assign n13193 = n402 & n9414 ;
  assign n13194 = n13192 | n13193 ;
  assign n13195 = n13194 ^ x53 ^ 1'b0 ;
  assign n13196 = n13195 ^ n13186 ^ n13105 ;
  assign n13197 = ( n13105 & ~n13186 ) | ( n13105 & n13195 ) | ( ~n13186 & n13195 ) ;
  assign n13198 = x107 & n208 ;
  assign n13199 = n197 & n8680 ;
  assign n13200 = ( x109 & n194 ) | ( x109 & n13198 ) | ( n194 & n13198 ) ;
  assign n13201 = n13198 | n13200 ;
  assign n13202 = x108 & ~n192 ;
  assign n13203 = ( x108 & n13201 ) | ( x108 & ~n13202 ) | ( n13201 & ~n13202 ) ;
  assign n13204 = x116 & n561 ;
  assign n13205 = n13199 | n13203 ;
  assign n13206 = ( x118 & n551 ) | ( x118 & n13204 ) | ( n551 & n13204 ) ;
  assign n13207 = n13204 | n13206 ;
  assign n13208 = x117 & ~n550 ;
  assign n13209 = ( x117 & n13207 ) | ( x117 & ~n13208 ) | ( n13207 & ~n13208 ) ;
  assign n13210 = n553 & n9671 ;
  assign n13211 = n13209 | n13210 ;
  assign n13212 = n13211 ^ x50 ^ 1'b0 ;
  assign n13213 = n197 & n8557 ;
  assign n13214 = n13212 ^ n13196 ^ n13115 ;
  assign n13215 = ( n13115 & ~n13196 ) | ( n13115 & n13212 ) | ( ~n13196 & n13212 ) ;
  assign n13216 = x106 & n208 ;
  assign n13217 = ( x108 & n194 ) | ( x108 & n13216 ) | ( n194 & n13216 ) ;
  assign n13218 = n13216 | n13217 ;
  assign n13219 = x107 & ~n192 ;
  assign n13220 = ( x107 & n13218 ) | ( x107 & ~n13219 ) | ( n13218 & ~n13219 ) ;
  assign n13221 = x119 & n744 ;
  assign n13222 = n13213 | n13220 ;
  assign n13223 = ( x121 & n730 ) | ( x121 & n13221 ) | ( n730 & n13221 ) ;
  assign n13224 = n13221 | n13223 ;
  assign n13225 = x120 & ~n732 ;
  assign n13226 = ( x120 & n13224 ) | ( x120 & ~n13225 ) | ( n13224 & ~n13225 ) ;
  assign n13227 = n731 & n9808 ;
  assign n13228 = n13226 | n13227 ;
  assign n13229 = n13228 ^ x47 ^ 1'b0 ;
  assign n13230 = n13229 ^ n13214 ^ n13125 ;
  assign n13231 = ( n13125 & ~n13214 ) | ( n13125 & n13229 ) | ( ~n13214 & n13229 ) ;
  assign n13232 = x122 & n888 ;
  assign n13233 = ( x124 & n878 ) | ( x124 & n13232 ) | ( n878 & n13232 ) ;
  assign n13234 = n13232 | n13233 ;
  assign n13235 = x123 & ~n877 ;
  assign n13236 = ( x123 & n13234 ) | ( x123 & ~n13235 ) | ( n13234 & ~n13235 ) ;
  assign n13237 = n880 & n9858 ;
  assign n13238 = n13236 | n13237 ;
  assign n13239 = n13238 ^ x44 ^ 1'b0 ;
  assign n13240 = n13239 ^ n13230 ^ n13135 ;
  assign n13241 = ( n13135 & ~n13230 ) | ( n13135 & n13239 ) | ( ~n13230 & n13239 ) ;
  assign n13242 = n13240 ^ n13178 ^ n13137 ;
  assign n13243 = n13242 ^ n13142 ^ n13141 ;
  assign n13244 = ( ~n13141 & n13142 ) | ( ~n13141 & n13242 ) | ( n13142 & n13242 ) ;
  assign n13245 = ( n13137 & n13178 ) | ( n13137 & ~n13240 ) | ( n13178 & ~n13240 ) ;
  assign n13246 = x108 & n133 ;
  assign n13247 = ( x110 & n142 ) | ( x110 & n13246 ) | ( n142 & n13246 ) ;
  assign n13248 = n13246 | n13247 ;
  assign n13249 = x109 & ~n134 ;
  assign n13250 = ( x109 & n13248 ) | ( x109 & ~n13249 ) | ( n13248 & ~n13249 ) ;
  assign n13251 = n140 & n8820 ;
  assign n13252 = n13250 | n13251 ;
  assign n13253 = x104 & ~n242 ;
  assign n13254 = x103 & n325 ;
  assign n13255 = ( x104 & ~n13253 ) | ( x104 & n13254 ) | ( ~n13253 & n13254 ) ;
  assign n13256 = ( n13153 & n13172 ) | ( n13153 & ~n13255 ) | ( n13172 & ~n13255 ) ;
  assign n13257 = n13255 ^ n13172 ^ n13153 ;
  assign n13258 = n13252 ^ x59 ^ 1'b0 ;
  assign n13259 = n13258 ^ n13257 ^ n13157 ;
  assign n13260 = ( n13157 & ~n13257 ) | ( n13157 & n13258 ) | ( ~n13257 & n13258 ) ;
  assign n13261 = x111 & n263 ;
  assign n13262 = ( x113 & n264 ) | ( x113 & n13261 ) | ( n264 & n13261 ) ;
  assign n13263 = n13261 | n13262 ;
  assign n13264 = x112 & ~n260 ;
  assign n13265 = ( x112 & n13263 ) | ( x112 & ~n13264 ) | ( n13263 & ~n13264 ) ;
  assign n13266 = n272 & n9199 ;
  assign n13267 = n13265 | n13266 ;
  assign n13268 = n13267 ^ x56 ^ 1'b0 ;
  assign n13269 = n13268 ^ n13259 ^ n13174 ;
  assign n13270 = ( n13174 & ~n13259 ) | ( n13174 & n13268 ) | ( ~n13259 & n13268 ) ;
  assign n13271 = x114 & n408 ;
  assign n13272 = ( x116 & n403 ) | ( x116 & n13271 ) | ( n403 & n13271 ) ;
  assign n13273 = n13271 | n13272 ;
  assign n13274 = x115 & ~n410 ;
  assign n13275 = ( x115 & n13273 ) | ( x115 & ~n13274 ) | ( n13273 & ~n13274 ) ;
  assign n13276 = n402 & n9513 ;
  assign n13277 = n13275 | n13276 ;
  assign n13278 = n13277 ^ x53 ^ 1'b0 ;
  assign n13279 = ( n13187 & ~n13269 ) | ( n13187 & n13278 ) | ( ~n13269 & n13278 ) ;
  assign n13280 = n13278 ^ n13269 ^ n13187 ;
  assign n13281 = x117 & n561 ;
  assign n13282 = ( x119 & n551 ) | ( x119 & n13281 ) | ( n551 & n13281 ) ;
  assign n13283 = n13281 | n13282 ;
  assign n13284 = x118 & ~n550 ;
  assign n13285 = ( x118 & n13283 ) | ( x118 & ~n13284 ) | ( n13283 & ~n13284 ) ;
  assign n13286 = n553 & n9733 ;
  assign n13287 = n13285 | n13286 ;
  assign n13288 = n13287 ^ x50 ^ 1'b0 ;
  assign n13289 = ( n13197 & ~n13280 ) | ( n13197 & n13288 ) | ( ~n13280 & n13288 ) ;
  assign n13290 = n13288 ^ n13280 ^ n13197 ;
  assign n13291 = x120 & n744 ;
  assign n13292 = ( x122 & n730 ) | ( x122 & n13291 ) | ( n730 & n13291 ) ;
  assign n13293 = n13291 | n13292 ;
  assign n13294 = x121 & ~n732 ;
  assign n13295 = ( x121 & n13293 ) | ( x121 & ~n13294 ) | ( n13293 & ~n13294 ) ;
  assign n13296 = n731 & n9806 ;
  assign n13297 = n13295 | n13296 ;
  assign n13298 = n13297 ^ x47 ^ 1'b0 ;
  assign n13299 = n13298 ^ n13290 ^ n13215 ;
  assign n13300 = ( n13215 & ~n13290 ) | ( n13215 & n13298 ) | ( ~n13290 & n13298 ) ;
  assign n13301 = x123 & n888 ;
  assign n13302 = ( x125 & n878 ) | ( x125 & n13301 ) | ( n878 & n13301 ) ;
  assign n13303 = n13301 | n13302 ;
  assign n13304 = x124 & ~n877 ;
  assign n13305 = ( x124 & n13303 ) | ( x124 & ~n13304 ) | ( n13303 & ~n13304 ) ;
  assign n13306 = n880 & n9883 ;
  assign n13307 = n13305 | n13306 ;
  assign n13308 = n13307 ^ x44 ^ 1'b0 ;
  assign n13309 = ( n13231 & ~n13299 ) | ( n13231 & n13308 ) | ( ~n13299 & n13308 ) ;
  assign n13310 = n13308 ^ n13299 ^ n13231 ;
  assign n13311 = x124 & n888 ;
  assign n13312 = ( x126 & n878 ) | ( x126 & n13311 ) | ( n878 & n13311 ) ;
  assign n13313 = n13311 | n13312 ;
  assign n13314 = x125 & n888 ;
  assign n13315 = ( x127 & n878 ) | ( x127 & n13314 ) | ( n878 & n13314 ) ;
  assign n13316 = n13314 | n13315 ;
  assign n13317 = x125 & ~n877 ;
  assign n13318 = ( x125 & n13313 ) | ( x125 & ~n13317 ) | ( n13313 & ~n13317 ) ;
  assign n13319 = x126 & ~n877 ;
  assign n13320 = ( x126 & n13316 ) | ( x126 & ~n13319 ) | ( n13316 & ~n13319 ) ;
  assign n13321 = n880 & n9949 ;
  assign n13322 = n13320 | n13321 ;
  assign n13323 = x127 & ~n877 ;
  assign n13324 = n880 & n9917 ;
  assign n13325 = n13318 | n13324 ;
  assign n13326 = ( n13177 & n13241 ) | ( n13177 & ~n13310 ) | ( n13241 & ~n13310 ) ;
  assign n13327 = n13310 ^ n13241 ^ n13177 ;
  assign n13328 = x126 & n888 ;
  assign n13329 = ( x127 & ~n13323 ) | ( x127 & n13328 ) | ( ~n13323 & n13328 ) ;
  assign n13330 = x127 & n888 ;
  assign n13331 = ( n880 & n9968 ) | ( n880 & n13330 ) | ( n9968 & n13330 ) ;
  assign n13332 = ( n880 & n9958 ) | ( n880 & n13328 ) | ( n9958 & n13328 ) ;
  assign n13333 = n13330 | n13331 ;
  assign n13334 = n13329 | n13332 ;
  assign n13335 = n13327 ^ n13245 ^ n13244 ;
  assign n13336 = ( n13244 & ~n13245 ) | ( n13244 & n13327 ) | ( ~n13245 & n13327 ) ;
  assign n13337 = x109 & n133 ;
  assign n13338 = ( x111 & n142 ) | ( x111 & n13337 ) | ( n142 & n13337 ) ;
  assign n13339 = n13337 | n13338 ;
  assign n13340 = n13078 ^ x41 ^ 1'b0 ;
  assign n13341 = x110 & ~n134 ;
  assign n13342 = ( x110 & n13339 ) | ( x110 & ~n13341 ) | ( n13339 & ~n13341 ) ;
  assign n13343 = n140 & n8946 ;
  assign n13344 = x105 & ~n242 ;
  assign n13345 = n13342 | n13343 ;
  assign n13346 = x104 & n325 ;
  assign n13347 = ( x105 & ~n13344 ) | ( x105 & n13346 ) | ( ~n13344 & n13346 ) ;
  assign n13348 = n13345 ^ x59 ^ 1'b0 ;
  assign n13349 = n13347 ^ n13256 ^ n13255 ;
  assign n13350 = ( ~n13255 & n13256 ) | ( ~n13255 & n13347 ) | ( n13256 & n13347 ) ;
  assign n13351 = n13222 ^ x62 ^ 1'b0 ;
  assign n13352 = ( n13348 & ~n13349 ) | ( n13348 & n13351 ) | ( ~n13349 & n13351 ) ;
  assign n13353 = n13351 ^ n13349 ^ n13348 ;
  assign n13354 = n13325 ^ x44 ^ 1'b0 ;
  assign n13355 = x112 & n263 ;
  assign n13356 = ( x114 & n264 ) | ( x114 & n13355 ) | ( n264 & n13355 ) ;
  assign n13357 = n13205 ^ x62 ^ 1'b0 ;
  assign n13358 = n13355 | n13356 ;
  assign n13359 = x113 & ~n260 ;
  assign n13360 = ( x113 & n13358 ) | ( x113 & ~n13359 ) | ( n13358 & ~n13359 ) ;
  assign n13361 = n272 & n9279 ;
  assign n13362 = n13360 | n13361 ;
  assign n13363 = n13362 ^ x56 ^ 1'b0 ;
  assign n13364 = n13363 ^ n13353 ^ n13260 ;
  assign n13365 = ( n13260 & ~n13353 ) | ( n13260 & n13363 ) | ( ~n13353 & n13363 ) ;
  assign n13366 = x115 & n408 ;
  assign n13367 = ( x117 & n403 ) | ( x117 & n13366 ) | ( n403 & n13366 ) ;
  assign n13368 = n13366 | n13367 ;
  assign n13369 = x116 & ~n410 ;
  assign n13370 = ( x116 & n13368 ) | ( x116 & ~n13369 ) | ( n13368 & ~n13369 ) ;
  assign n13371 = n402 & n9569 ;
  assign n13372 = n13370 | n13371 ;
  assign n13373 = n13372 ^ x53 ^ 1'b0 ;
  assign n13374 = ( n13270 & ~n13364 ) | ( n13270 & n13373 ) | ( ~n13364 & n13373 ) ;
  assign n13375 = n13373 ^ n13364 ^ n13270 ;
  assign n13376 = x118 & n561 ;
  assign n13377 = ( x120 & n551 ) | ( x120 & n13376 ) | ( n551 & n13376 ) ;
  assign n13378 = n13376 | n13377 ;
  assign n13379 = x119 & ~n550 ;
  assign n13380 = ( x119 & n13378 ) | ( x119 & ~n13379 ) | ( n13378 & ~n13379 ) ;
  assign n13381 = n553 & n9756 ;
  assign n13382 = n13380 | n13381 ;
  assign n13383 = n13382 ^ x50 ^ 1'b0 ;
  assign n13384 = n13383 ^ n13375 ^ n13279 ;
  assign n13385 = ( n13279 & ~n13375 ) | ( n13279 & n13383 ) | ( ~n13375 & n13383 ) ;
  assign n13386 = x121 & n744 ;
  assign n13387 = ( x123 & n730 ) | ( x123 & n13386 ) | ( n730 & n13386 ) ;
  assign n13388 = n13386 | n13387 ;
  assign n13389 = x122 & ~n732 ;
  assign n13390 = ( x122 & n13388 ) | ( x122 & ~n13389 ) | ( n13388 & ~n13389 ) ;
  assign n13391 = n731 & n9828 ;
  assign n13392 = n13390 | n13391 ;
  assign n13393 = n13392 ^ x47 ^ 1'b0 ;
  assign n13394 = ( n13289 & ~n13384 ) | ( n13289 & n13393 ) | ( ~n13384 & n13393 ) ;
  assign n13395 = n13393 ^ n13384 ^ n13289 ;
  assign n13396 = n13395 ^ n13354 ^ n13300 ;
  assign n13397 = ( n13309 & n13340 ) | ( n13309 & ~n13396 ) | ( n13340 & ~n13396 ) ;
  assign n13398 = ( n13300 & n13354 ) | ( n13300 & ~n13395 ) | ( n13354 & ~n13395 ) ;
  assign n13399 = n13396 ^ n13340 ^ n13309 ;
  assign n13400 = ( ~n13326 & n13336 ) | ( ~n13326 & n13399 ) | ( n13336 & n13399 ) ;
  assign n13401 = n13399 ^ n13336 ^ n13326 ;
  assign n13402 = x105 & n325 ;
  assign n13403 = x106 & ~n242 ;
  assign n13404 = ( x106 & n13402 ) | ( x106 & ~n13403 ) | ( n13402 & ~n13403 ) ;
  assign n13405 = n13404 ^ n13255 ^ x41 ;
  assign n13406 = ( ~x41 & n13255 ) | ( ~x41 & n13404 ) | ( n13255 & n13404 ) ;
  assign n13407 = ( n13350 & n13357 ) | ( n13350 & ~n13405 ) | ( n13357 & ~n13405 ) ;
  assign n13408 = n13405 ^ n13357 ^ n13350 ;
  assign n13409 = x110 & n133 ;
  assign n13410 = ( x112 & n142 ) | ( x112 & n13409 ) | ( n142 & n13409 ) ;
  assign n13411 = n13409 | n13410 ;
  assign n13412 = x111 & ~n134 ;
  assign n13413 = ( x111 & n13411 ) | ( x111 & ~n13412 ) | ( n13411 & ~n13412 ) ;
  assign n13414 = n140 & n9080 ;
  assign n13415 = n13413 | n13414 ;
  assign n13416 = n13415 ^ x59 ^ 1'b0 ;
  assign n13417 = ( n13352 & ~n13408 ) | ( n13352 & n13416 ) | ( ~n13408 & n13416 ) ;
  assign n13418 = n13416 ^ n13408 ^ n13352 ;
  assign n13419 = x113 & n263 ;
  assign n13420 = ( x115 & n264 ) | ( x115 & n13419 ) | ( n264 & n13419 ) ;
  assign n13421 = n13419 | n13420 ;
  assign n13422 = x114 & ~n260 ;
  assign n13423 = ( x114 & n13421 ) | ( x114 & ~n13422 ) | ( n13421 & ~n13422 ) ;
  assign n13424 = n272 & n9414 ;
  assign n13425 = n13423 | n13424 ;
  assign n13426 = n13425 ^ x56 ^ 1'b0 ;
  assign n13427 = n13426 ^ n13418 ^ n13365 ;
  assign n13428 = ( n13365 & ~n13418 ) | ( n13365 & n13426 ) | ( ~n13418 & n13426 ) ;
  assign n13429 = x116 & n408 ;
  assign n13430 = ( x118 & n403 ) | ( x118 & n13429 ) | ( n403 & n13429 ) ;
  assign n13431 = n13429 | n13430 ;
  assign n13432 = x117 & ~n410 ;
  assign n13433 = ( x117 & n13431 ) | ( x117 & ~n13432 ) | ( n13431 & ~n13432 ) ;
  assign n13434 = n402 & n9671 ;
  assign n13435 = n13433 | n13434 ;
  assign n13436 = n13435 ^ x53 ^ 1'b0 ;
  assign n13437 = n13436 ^ n13427 ^ n13374 ;
  assign n13438 = ( n13374 & ~n13427 ) | ( n13374 & n13436 ) | ( ~n13427 & n13436 ) ;
  assign n13439 = x119 & n561 ;
  assign n13440 = ( x121 & n551 ) | ( x121 & n13439 ) | ( n551 & n13439 ) ;
  assign n13441 = n13439 | n13440 ;
  assign n13442 = x120 & ~n550 ;
  assign n13443 = ( x120 & n13441 ) | ( x120 & ~n13442 ) | ( n13441 & ~n13442 ) ;
  assign n13444 = n553 & n9808 ;
  assign n13445 = n13443 | n13444 ;
  assign n13446 = n13445 ^ x50 ^ 1'b0 ;
  assign n13447 = ( n13385 & ~n13437 ) | ( n13385 & n13446 ) | ( ~n13437 & n13446 ) ;
  assign n13448 = n13446 ^ n13437 ^ n13385 ;
  assign n13449 = x108 & n208 ;
  assign n13450 = ( x110 & n194 ) | ( x110 & n13449 ) | ( n194 & n13449 ) ;
  assign n13451 = n13449 | n13450 ;
  assign n13452 = x109 & ~n192 ;
  assign n13453 = ( x109 & n13451 ) | ( x109 & ~n13452 ) | ( n13451 & ~n13452 ) ;
  assign n13454 = ( n197 & n8820 ) | ( n197 & n13453 ) | ( n8820 & n13453 ) ;
  assign n13455 = n13453 | n13454 ;
  assign n13456 = n13322 ^ x44 ^ 1'b0 ;
  assign n13457 = x122 & n744 ;
  assign n13458 = ( x124 & n730 ) | ( x124 & n13457 ) | ( n730 & n13457 ) ;
  assign n13459 = n13457 | n13458 ;
  assign n13460 = x123 & ~n732 ;
  assign n13461 = ( x123 & n13459 ) | ( x123 & ~n13460 ) | ( n13459 & ~n13460 ) ;
  assign n13462 = n731 & n9858 ;
  assign n13463 = n13461 | n13462 ;
  assign n13464 = n13463 ^ x47 ^ 1'b0 ;
  assign n13465 = n13464 ^ n13448 ^ n13394 ;
  assign n13466 = ( n13394 & ~n13448 ) | ( n13394 & n13464 ) | ( ~n13448 & n13464 ) ;
  assign n13467 = n13465 ^ n13456 ^ n13398 ;
  assign n13468 = ( ~n13397 & n13400 ) | ( ~n13397 & n13467 ) | ( n13400 & n13467 ) ;
  assign n13469 = ( n13398 & n13456 ) | ( n13398 & ~n13465 ) | ( n13456 & ~n13465 ) ;
  assign n13470 = x123 & n744 ;
  assign n13471 = ( x125 & n730 ) | ( x125 & n13470 ) | ( n730 & n13470 ) ;
  assign n13472 = n13470 | n13471 ;
  assign n13473 = x124 & ~n732 ;
  assign n13474 = n13467 ^ n13400 ^ n13397 ;
  assign n13475 = x124 & n744 ;
  assign n13476 = ( x124 & n13472 ) | ( x124 & ~n13473 ) | ( n13472 & ~n13473 ) ;
  assign n13477 = x125 & n744 ;
  assign n13478 = ( x127 & n730 ) | ( x127 & n13477 ) | ( n730 & n13477 ) ;
  assign n13479 = ( x126 & n730 ) | ( x126 & n13475 ) | ( n730 & n13475 ) ;
  assign n13480 = n13477 | n13478 ;
  assign n13481 = n13475 | n13479 ;
  assign n13482 = n13334 ^ x44 ^ 1'b0 ;
  assign n13483 = x127 & n744 ;
  assign n13484 = ( n731 & n9968 ) | ( n731 & n13483 ) | ( n9968 & n13483 ) ;
  assign n13485 = n13483 | n13484 ;
  assign n13486 = x125 & ~n732 ;
  assign n13487 = ( x125 & n13481 ) | ( x125 & ~n13486 ) | ( n13481 & ~n13486 ) ;
  assign n13488 = n731 & n9917 ;
  assign n13489 = n13487 | n13488 ;
  assign n13490 = n731 & n9883 ;
  assign n13491 = n13476 | n13490 ;
  assign n13492 = x127 & ~n732 ;
  assign n13493 = x126 & n744 ;
  assign n13494 = ( x127 & ~n13492 ) | ( x127 & n13493 ) | ( ~n13492 & n13493 ) ;
  assign n13495 = ( n731 & n9958 ) | ( n731 & n13493 ) | ( n9958 & n13493 ) ;
  assign n13496 = n731 & n9949 ;
  assign n13497 = x126 & ~n732 ;
  assign n13498 = ( x126 & n13480 ) | ( x126 & ~n13497 ) | ( n13480 & ~n13497 ) ;
  assign n13499 = n13496 | n13498 ;
  assign n13500 = n13489 ^ x47 ^ 1'b0 ;
  assign n13501 = n13485 ^ x47 ^ 1'b0 ;
  assign n13502 = n13491 ^ x47 ^ 1'b0 ;
  assign n13503 = n13494 | n13495 ;
  assign n13504 = n13455 ^ x62 ^ 1'b0 ;
  assign n13505 = x107 & ~n242 ;
  assign n13506 = x111 & n133 ;
  assign n13507 = x106 & n325 ;
  assign n13508 = ( x107 & ~n13505 ) | ( x107 & n13507 ) | ( ~n13505 & n13507 ) ;
  assign n13509 = ( x113 & n142 ) | ( x113 & n13506 ) | ( n142 & n13506 ) ;
  assign n13510 = n13506 | n13509 ;
  assign n13511 = ( n13406 & n13504 ) | ( n13406 & ~n13508 ) | ( n13504 & ~n13508 ) ;
  assign n13512 = n13508 ^ n13504 ^ n13406 ;
  assign n13513 = x112 & ~n134 ;
  assign n13514 = ( x112 & n13510 ) | ( x112 & ~n13513 ) | ( n13510 & ~n13513 ) ;
  assign n13515 = n140 & n9199 ;
  assign n13516 = n13514 | n13515 ;
  assign n13517 = n13516 ^ x59 ^ 1'b0 ;
  assign n13518 = ( n13407 & ~n13512 ) | ( n13407 & n13517 ) | ( ~n13512 & n13517 ) ;
  assign n13519 = n13517 ^ n13512 ^ n13407 ;
  assign n13520 = x114 & n263 ;
  assign n13521 = ( x116 & n264 ) | ( x116 & n13520 ) | ( n264 & n13520 ) ;
  assign n13522 = n13520 | n13521 ;
  assign n13523 = x115 & ~n260 ;
  assign n13524 = ( x115 & n13522 ) | ( x115 & ~n13523 ) | ( n13522 & ~n13523 ) ;
  assign n13525 = n272 & n9513 ;
  assign n13526 = n13524 | n13525 ;
  assign n13527 = n13526 ^ x56 ^ 1'b0 ;
  assign n13528 = ( n13417 & ~n13519 ) | ( n13417 & n13527 ) | ( ~n13519 & n13527 ) ;
  assign n13529 = n13527 ^ n13519 ^ n13417 ;
  assign n13530 = x117 & n408 ;
  assign n13531 = ( x119 & n403 ) | ( x119 & n13530 ) | ( n403 & n13530 ) ;
  assign n13532 = n13530 | n13531 ;
  assign n13533 = x118 & ~n410 ;
  assign n13534 = ( x118 & n13532 ) | ( x118 & ~n13533 ) | ( n13532 & ~n13533 ) ;
  assign n13535 = n402 & n9733 ;
  assign n13536 = n13534 | n13535 ;
  assign n13537 = n13536 ^ x53 ^ 1'b0 ;
  assign n13538 = ( n13428 & ~n13529 ) | ( n13428 & n13537 ) | ( ~n13529 & n13537 ) ;
  assign n13539 = n13537 ^ n13529 ^ n13428 ;
  assign n13540 = x120 & n561 ;
  assign n13541 = ( x122 & n551 ) | ( x122 & n13540 ) | ( n551 & n13540 ) ;
  assign n13542 = n13540 | n13541 ;
  assign n13543 = x121 & ~n550 ;
  assign n13544 = ( x121 & n13542 ) | ( x121 & ~n13543 ) | ( n13542 & ~n13543 ) ;
  assign n13545 = n553 & n9806 ;
  assign n13546 = n13544 | n13545 ;
  assign n13547 = n13546 ^ x50 ^ 1'b0 ;
  assign n13548 = ( n13438 & ~n13539 ) | ( n13438 & n13547 ) | ( ~n13539 & n13547 ) ;
  assign n13549 = n13547 ^ n13539 ^ n13438 ;
  assign n13550 = n13549 ^ n13502 ^ n13447 ;
  assign n13551 = ( n13447 & n13502 ) | ( n13447 & ~n13549 ) | ( n13502 & ~n13549 ) ;
  assign n13552 = n13550 ^ n13482 ^ n13466 ;
  assign n13553 = ( n13466 & n13482 ) | ( n13466 & ~n13550 ) | ( n13482 & ~n13550 ) ;
  assign n13554 = ( n13468 & ~n13469 ) | ( n13468 & n13552 ) | ( ~n13469 & n13552 ) ;
  assign n13555 = n13552 ^ n13469 ^ n13468 ;
  assign n13556 = x109 & n208 ;
  assign n13557 = x108 & ~n242 ;
  assign n13558 = x107 & n325 ;
  assign n13559 = ( x108 & ~n13557 ) | ( x108 & n13558 ) | ( ~n13557 & n13558 ) ;
  assign n13560 = ( x111 & n194 ) | ( x111 & n13556 ) | ( n194 & n13556 ) ;
  assign n13561 = n13556 | n13560 ;
  assign n13562 = x110 & ~n192 ;
  assign n13563 = ( x110 & n13561 ) | ( x110 & ~n13562 ) | ( n13561 & ~n13562 ) ;
  assign n13564 = ( n197 & n8946 ) | ( n197 & n13563 ) | ( n8946 & n13563 ) ;
  assign n13565 = n13563 | n13564 ;
  assign n13566 = n13565 ^ x62 ^ 1'b0 ;
  assign n13567 = n13566 ^ n13559 ^ n13508 ;
  assign n13568 = x112 & n133 ;
  assign n13569 = ( ~n13508 & n13559 ) | ( ~n13508 & n13566 ) | ( n13559 & n13566 ) ;
  assign n13570 = ( x114 & n142 ) | ( x114 & n13568 ) | ( n142 & n13568 ) ;
  assign n13571 = n13568 | n13570 ;
  assign n13572 = x113 & ~n134 ;
  assign n13573 = ( x113 & n13571 ) | ( x113 & ~n13572 ) | ( n13571 & ~n13572 ) ;
  assign n13574 = n140 & n9279 ;
  assign n13575 = n13573 | n13574 ;
  assign n13576 = n13575 ^ x59 ^ 1'b0 ;
  assign n13577 = n13576 ^ n13567 ^ n13511 ;
  assign n13578 = ( n13511 & ~n13567 ) | ( n13511 & n13576 ) | ( ~n13567 & n13576 ) ;
  assign n13579 = x115 & n263 ;
  assign n13580 = ( x117 & n264 ) | ( x117 & n13579 ) | ( n264 & n13579 ) ;
  assign n13581 = n13579 | n13580 ;
  assign n13582 = x116 & ~n260 ;
  assign n13583 = ( x116 & n13581 ) | ( x116 & ~n13582 ) | ( n13581 & ~n13582 ) ;
  assign n13584 = n272 & n9569 ;
  assign n13585 = n13583 | n13584 ;
  assign n13586 = n13585 ^ x56 ^ 1'b0 ;
  assign n13587 = n13586 ^ n13577 ^ n13518 ;
  assign n13588 = ( n13518 & ~n13577 ) | ( n13518 & n13586 ) | ( ~n13577 & n13586 ) ;
  assign n13589 = x118 & n408 ;
  assign n13590 = ( x120 & n403 ) | ( x120 & n13589 ) | ( n403 & n13589 ) ;
  assign n13591 = n13589 | n13590 ;
  assign n13592 = x119 & ~n410 ;
  assign n13593 = ( x119 & n13591 ) | ( x119 & ~n13592 ) | ( n13591 & ~n13592 ) ;
  assign n13594 = n402 & n9756 ;
  assign n13595 = n13593 | n13594 ;
  assign n13596 = n13595 ^ x53 ^ 1'b0 ;
  assign n13597 = ( n13528 & ~n13587 ) | ( n13528 & n13596 ) | ( ~n13587 & n13596 ) ;
  assign n13598 = n13596 ^ n13587 ^ n13528 ;
  assign n13599 = x121 & n561 ;
  assign n13600 = ( x123 & n551 ) | ( x123 & n13599 ) | ( n551 & n13599 ) ;
  assign n13601 = n13599 | n13600 ;
  assign n13602 = n13333 ^ x44 ^ 1'b0 ;
  assign n13603 = x122 & ~n550 ;
  assign n13604 = ( x122 & n13601 ) | ( x122 & ~n13603 ) | ( n13601 & ~n13603 ) ;
  assign n13605 = n553 & n9828 ;
  assign n13606 = n13604 | n13605 ;
  assign n13607 = n13606 ^ x50 ^ 1'b0 ;
  assign n13608 = n13607 ^ n13598 ^ n13538 ;
  assign n13609 = ( n13538 & ~n13598 ) | ( n13538 & n13607 ) | ( ~n13598 & n13607 ) ;
  assign n13610 = ( n13500 & n13548 ) | ( n13500 & ~n13608 ) | ( n13548 & ~n13608 ) ;
  assign n13611 = n13608 ^ n13548 ^ n13500 ;
  assign n13612 = n13611 ^ n13602 ^ n13551 ;
  assign n13613 = ( n13551 & n13602 ) | ( n13551 & ~n13611 ) | ( n13602 & ~n13611 ) ;
  assign n13614 = ( ~n13553 & n13554 ) | ( ~n13553 & n13612 ) | ( n13554 & n13612 ) ;
  assign n13615 = n13612 ^ n13554 ^ n13553 ;
  assign n13616 = x110 & n208 ;
  assign n13617 = ( x112 & n194 ) | ( x112 & n13616 ) | ( n194 & n13616 ) ;
  assign n13618 = n13616 | n13617 ;
  assign n13619 = x111 & ~n192 ;
  assign n13620 = ( x111 & n13618 ) | ( x111 & ~n13619 ) | ( n13618 & ~n13619 ) ;
  assign n13621 = x109 & ~n242 ;
  assign n13622 = n197 & n9080 ;
  assign n13623 = n13620 | n13622 ;
  assign n13624 = x108 & n325 ;
  assign n13625 = ( x109 & ~n13621 ) | ( x109 & n13624 ) | ( ~n13621 & n13624 ) ;
  assign n13626 = ( ~x44 & n13508 ) | ( ~x44 & n13625 ) | ( n13508 & n13625 ) ;
  assign n13627 = n13623 ^ x62 ^ 1'b0 ;
  assign n13628 = n13625 ^ n13508 ^ x44 ;
  assign n13629 = ( n13569 & n13627 ) | ( n13569 & ~n13628 ) | ( n13627 & ~n13628 ) ;
  assign n13630 = n13628 ^ n13627 ^ n13569 ;
  assign n13631 = x113 & n133 ;
  assign n13632 = ( x115 & n142 ) | ( x115 & n13631 ) | ( n142 & n13631 ) ;
  assign n13633 = n13631 | n13632 ;
  assign n13634 = x114 & ~n134 ;
  assign n13635 = ( x114 & n13633 ) | ( x114 & ~n13634 ) | ( n13633 & ~n13634 ) ;
  assign n13636 = n140 & n9414 ;
  assign n13637 = n13635 | n13636 ;
  assign n13638 = n13637 ^ x59 ^ 1'b0 ;
  assign n13639 = ( n13578 & ~n13630 ) | ( n13578 & n13638 ) | ( ~n13630 & n13638 ) ;
  assign n13640 = n13638 ^ n13630 ^ n13578 ;
  assign n13641 = x116 & n263 ;
  assign n13642 = n197 & n9199 ;
  assign n13643 = ( x118 & n264 ) | ( x118 & n13641 ) | ( n264 & n13641 ) ;
  assign n13644 = n13641 | n13643 ;
  assign n13645 = x117 & ~n260 ;
  assign n13646 = ( x117 & n13644 ) | ( x117 & ~n13645 ) | ( n13644 & ~n13645 ) ;
  assign n13647 = n272 & n9671 ;
  assign n13648 = n13646 | n13647 ;
  assign n13649 = n13648 ^ x56 ^ 1'b0 ;
  assign n13650 = n13649 ^ n13640 ^ n13588 ;
  assign n13651 = ( n13588 & ~n13640 ) | ( n13588 & n13649 ) | ( ~n13640 & n13649 ) ;
  assign n13652 = x119 & n408 ;
  assign n13653 = ( x121 & n403 ) | ( x121 & n13652 ) | ( n403 & n13652 ) ;
  assign n13654 = n13652 | n13653 ;
  assign n13655 = n13499 ^ x47 ^ 1'b0 ;
  assign n13656 = x120 & ~n410 ;
  assign n13657 = ( x120 & n13654 ) | ( x120 & ~n13656 ) | ( n13654 & ~n13656 ) ;
  assign n13658 = n402 & n9808 ;
  assign n13659 = n13657 | n13658 ;
  assign n13660 = n13659 ^ x53 ^ 1'b0 ;
  assign n13661 = ( n13597 & ~n13650 ) | ( n13597 & n13660 ) | ( ~n13650 & n13660 ) ;
  assign n13662 = n13660 ^ n13650 ^ n13597 ;
  assign n13663 = x122 & n561 ;
  assign n13664 = ( x124 & n551 ) | ( x124 & n13663 ) | ( n551 & n13663 ) ;
  assign n13665 = n13663 | n13664 ;
  assign n13666 = x123 & ~n550 ;
  assign n13667 = ( x123 & n13665 ) | ( x123 & ~n13666 ) | ( n13665 & ~n13666 ) ;
  assign n13668 = n553 & n9858 ;
  assign n13669 = n13667 | n13668 ;
  assign n13670 = n13669 ^ x50 ^ 1'b0 ;
  assign n13671 = ( n13609 & ~n13662 ) | ( n13609 & n13670 ) | ( ~n13662 & n13670 ) ;
  assign n13672 = n13670 ^ n13662 ^ n13609 ;
  assign n13673 = ( n13610 & n13655 ) | ( n13610 & ~n13672 ) | ( n13655 & ~n13672 ) ;
  assign n13674 = n13672 ^ n13655 ^ n13610 ;
  assign n13675 = ( ~n13613 & n13614 ) | ( ~n13613 & n13674 ) | ( n13614 & n13674 ) ;
  assign n13676 = n13674 ^ n13614 ^ n13613 ;
  assign n13677 = x111 & n208 ;
  assign n13678 = x110 & ~n242 ;
  assign n13679 = ( x113 & n194 ) | ( x113 & n13677 ) | ( n194 & n13677 ) ;
  assign n13680 = n13677 | n13679 ;
  assign n13681 = x112 & ~n192 ;
  assign n13682 = ( x112 & n13680 ) | ( x112 & ~n13681 ) | ( n13680 & ~n13681 ) ;
  assign n13683 = n13642 | n13682 ;
  assign n13684 = x114 & n133 ;
  assign n13685 = ( x116 & n142 ) | ( x116 & n13684 ) | ( n142 & n13684 ) ;
  assign n13686 = n13684 | n13685 ;
  assign n13687 = x109 & n325 ;
  assign n13688 = ( x110 & ~n13678 ) | ( x110 & n13687 ) | ( ~n13678 & n13687 ) ;
  assign n13689 = x115 & ~n134 ;
  assign n13690 = ( x115 & n13686 ) | ( x115 & ~n13689 ) | ( n13686 & ~n13689 ) ;
  assign n13691 = n13683 ^ x62 ^ 1'b0 ;
  assign n13692 = n140 & n9513 ;
  assign n13693 = n13690 | n13692 ;
  assign n13694 = n13693 ^ x59 ^ 1'b0 ;
  assign n13695 = ( n13626 & ~n13688 ) | ( n13626 & n13691 ) | ( ~n13688 & n13691 ) ;
  assign n13696 = n13691 ^ n13688 ^ n13626 ;
  assign n13697 = ( n13629 & n13694 ) | ( n13629 & ~n13696 ) | ( n13694 & ~n13696 ) ;
  assign n13698 = n13696 ^ n13694 ^ n13629 ;
  assign n13699 = x117 & n263 ;
  assign n13700 = ( x119 & n264 ) | ( x119 & n13699 ) | ( n264 & n13699 ) ;
  assign n13701 = n13699 | n13700 ;
  assign n13702 = x118 & ~n260 ;
  assign n13703 = ( x118 & n13701 ) | ( x118 & ~n13702 ) | ( n13701 & ~n13702 ) ;
  assign n13704 = n272 & n9733 ;
  assign n13705 = n13703 | n13704 ;
  assign n13706 = n13705 ^ x56 ^ 1'b0 ;
  assign n13707 = n13706 ^ n13698 ^ n13639 ;
  assign n13708 = ( n13639 & ~n13698 ) | ( n13639 & n13706 ) | ( ~n13698 & n13706 ) ;
  assign n13709 = x120 & n408 ;
  assign n13710 = n13503 ^ x47 ^ 1'b0 ;
  assign n13711 = ( x122 & n403 ) | ( x122 & n13709 ) | ( n403 & n13709 ) ;
  assign n13712 = n13709 | n13711 ;
  assign n13713 = x121 & ~n410 ;
  assign n13714 = ( x121 & n13712 ) | ( x121 & ~n13713 ) | ( n13712 & ~n13713 ) ;
  assign n13715 = n402 & n9806 ;
  assign n13716 = n13714 | n13715 ;
  assign n13717 = n13716 ^ x53 ^ 1'b0 ;
  assign n13718 = n13717 ^ n13707 ^ n13651 ;
  assign n13719 = ( n13651 & ~n13707 ) | ( n13651 & n13717 ) | ( ~n13707 & n13717 ) ;
  assign n13720 = x123 & n561 ;
  assign n13721 = ( x125 & n551 ) | ( x125 & n13720 ) | ( n551 & n13720 ) ;
  assign n13722 = n13720 | n13721 ;
  assign n13723 = x124 & ~n550 ;
  assign n13724 = ( x124 & n13722 ) | ( x124 & ~n13723 ) | ( n13722 & ~n13723 ) ;
  assign n13725 = n553 & n9883 ;
  assign n13726 = n13724 | n13725 ;
  assign n13727 = n13726 ^ x50 ^ 1'b0 ;
  assign n13728 = ( n13661 & ~n13718 ) | ( n13661 & n13727 ) | ( ~n13718 & n13727 ) ;
  assign n13729 = n13727 ^ n13718 ^ n13661 ;
  assign n13730 = ( n13671 & n13710 ) | ( n13671 & ~n13729 ) | ( n13710 & ~n13729 ) ;
  assign n13731 = n13729 ^ n13710 ^ n13671 ;
  assign n13732 = n13731 ^ n13675 ^ n13673 ;
  assign n13733 = ( ~n13673 & n13675 ) | ( ~n13673 & n13731 ) | ( n13675 & n13731 ) ;
  assign n13734 = x112 & n208 ;
  assign n13735 = ( x114 & n194 ) | ( x114 & n13734 ) | ( n194 & n13734 ) ;
  assign n13736 = n13734 | n13735 ;
  assign n13737 = x113 & ~n192 ;
  assign n13738 = ( x113 & n13736 ) | ( x113 & ~n13737 ) | ( n13736 & ~n13737 ) ;
  assign n13739 = x114 & n208 ;
  assign n13740 = n197 & n9279 ;
  assign n13741 = n13738 | n13740 ;
  assign n13742 = ( x116 & n194 ) | ( x116 & n13739 ) | ( n194 & n13739 ) ;
  assign n13743 = n13739 | n13742 ;
  assign n13744 = x115 & ~n192 ;
  assign n13745 = ( x115 & n13743 ) | ( x115 & ~n13744 ) | ( n13743 & ~n13744 ) ;
  assign n13746 = x124 & n561 ;
  assign n13747 = ( n197 & n9513 ) | ( n197 & n13745 ) | ( n9513 & n13745 ) ;
  assign n13748 = n197 & n9414 ;
  assign n13749 = n13745 | n13747 ;
  assign n13750 = ( x126 & n551 ) | ( x126 & n13746 ) | ( n551 & n13746 ) ;
  assign n13751 = n13746 | n13750 ;
  assign n13752 = x125 & ~n550 ;
  assign n13753 = ( x125 & n13751 ) | ( x125 & ~n13752 ) | ( n13751 & ~n13752 ) ;
  assign n13754 = x125 & n561 ;
  assign n13755 = ( x127 & n551 ) | ( x127 & n13754 ) | ( n551 & n13754 ) ;
  assign n13756 = n13754 | n13755 ;
  assign n13757 = x127 & ~n550 ;
  assign n13758 = x126 & ~n550 ;
  assign n13759 = ( x126 & n13756 ) | ( x126 & ~n13758 ) | ( n13756 & ~n13758 ) ;
  assign n13760 = n553 & n9917 ;
  assign n13761 = n13753 | n13760 ;
  assign n13762 = x127 & n561 ;
  assign n13763 = x126 & n561 ;
  assign n13764 = ( x127 & ~n13757 ) | ( x127 & n13763 ) | ( ~n13757 & n13763 ) ;
  assign n13765 = ( n553 & n9958 ) | ( n553 & n13763 ) | ( n9958 & n13763 ) ;
  assign n13766 = n13764 | n13765 ;
  assign n13767 = ( n553 & n9968 ) | ( n553 & n13762 ) | ( n9968 & n13762 ) ;
  assign n13768 = n13762 | n13767 ;
  assign n13769 = x113 & n208 ;
  assign n13770 = n553 & n9949 ;
  assign n13771 = n13759 | n13770 ;
  assign n13772 = ( x115 & n194 ) | ( x115 & n13769 ) | ( n194 & n13769 ) ;
  assign n13773 = n13769 | n13772 ;
  assign n13774 = x114 & ~n192 ;
  assign n13775 = ( x114 & n13773 ) | ( x114 & ~n13774 ) | ( n13773 & ~n13774 ) ;
  assign n13776 = n13748 | n13775 ;
  assign n13777 = x110 & n325 ;
  assign n13778 = x111 & ~n242 ;
  assign n13779 = ( x111 & n13777 ) | ( x111 & ~n13778 ) | ( n13777 & ~n13778 ) ;
  assign n13780 = n13779 ^ n13695 ^ n13688 ;
  assign n13781 = ( n13688 & n13695 ) | ( n13688 & ~n13779 ) | ( n13695 & ~n13779 ) ;
  assign n13782 = x115 & n133 ;
  assign n13783 = ( x117 & n142 ) | ( x117 & n13782 ) | ( n142 & n13782 ) ;
  assign n13784 = n13782 | n13783 ;
  assign n13785 = x116 & ~n134 ;
  assign n13786 = ( x116 & n13784 ) | ( x116 & ~n13785 ) | ( n13784 & ~n13785 ) ;
  assign n13787 = n13761 ^ x50 ^ 1'b0 ;
  assign n13788 = n140 & n9569 ;
  assign n13789 = n13786 | n13788 ;
  assign n13790 = n13741 ^ x62 ^ 1'b0 ;
  assign n13791 = n13789 ^ x59 ^ 1'b0 ;
  assign n13792 = ( ~n13780 & n13790 ) | ( ~n13780 & n13791 ) | ( n13790 & n13791 ) ;
  assign n13793 = n13791 ^ n13790 ^ n13780 ;
  assign n13794 = x118 & n263 ;
  assign n13795 = ( x120 & n264 ) | ( x120 & n13794 ) | ( n264 & n13794 ) ;
  assign n13796 = n13794 | n13795 ;
  assign n13797 = x119 & ~n260 ;
  assign n13798 = ( x119 & n13796 ) | ( x119 & ~n13797 ) | ( n13796 & ~n13797 ) ;
  assign n13799 = n272 & n9756 ;
  assign n13800 = n13798 | n13799 ;
  assign n13801 = n13800 ^ x56 ^ 1'b0 ;
  assign n13802 = ( n13697 & ~n13793 ) | ( n13697 & n13801 ) | ( ~n13793 & n13801 ) ;
  assign n13803 = n13801 ^ n13793 ^ n13697 ;
  assign n13804 = x121 & n408 ;
  assign n13805 = ( x123 & n403 ) | ( x123 & n13804 ) | ( n403 & n13804 ) ;
  assign n13806 = n13804 | n13805 ;
  assign n13807 = x122 & ~n410 ;
  assign n13808 = ( x122 & n13806 ) | ( x122 & ~n13807 ) | ( n13806 & ~n13807 ) ;
  assign n13809 = n402 & n9828 ;
  assign n13810 = n13808 | n13809 ;
  assign n13811 = n13810 ^ x53 ^ 1'b0 ;
  assign n13812 = n13776 ^ x62 ^ 1'b0 ;
  assign n13813 = ( n13708 & ~n13803 ) | ( n13708 & n13811 ) | ( ~n13803 & n13811 ) ;
  assign n13814 = n13811 ^ n13803 ^ n13708 ;
  assign n13815 = x111 & n325 ;
  assign n13816 = x112 & ~n242 ;
  assign n13817 = ( x112 & n13815 ) | ( x112 & ~n13816 ) | ( n13815 & ~n13816 ) ;
  assign n13818 = ( ~x47 & n13779 ) | ( ~x47 & n13817 ) | ( n13779 & n13817 ) ;
  assign n13819 = n13817 ^ n13779 ^ x47 ;
  assign n13820 = n13819 ^ n13812 ^ n13781 ;
  assign n13821 = ( n13781 & n13812 ) | ( n13781 & ~n13819 ) | ( n13812 & ~n13819 ) ;
  assign n13822 = n13814 ^ n13787 ^ n13719 ;
  assign n13823 = ( n13719 & n13787 ) | ( n13719 & ~n13814 ) | ( n13787 & ~n13814 ) ;
  assign n13824 = ( n13501 & n13728 ) | ( n13501 & ~n13822 ) | ( n13728 & ~n13822 ) ;
  assign n13825 = n13822 ^ n13728 ^ n13501 ;
  assign n13826 = n13825 ^ n13733 ^ n13730 ;
  assign n13827 = ( ~n13730 & n13733 ) | ( ~n13730 & n13825 ) | ( n13733 & n13825 ) ;
  assign n13828 = x116 & n133 ;
  assign n13829 = ( x118 & n142 ) | ( x118 & n13828 ) | ( n142 & n13828 ) ;
  assign n13830 = n13828 | n13829 ;
  assign n13831 = x117 & ~n134 ;
  assign n13832 = ( x117 & n13830 ) | ( x117 & ~n13831 ) | ( n13830 & ~n13831 ) ;
  assign n13833 = n140 & n9671 ;
  assign n13834 = n13832 | n13833 ;
  assign n13835 = n13834 ^ x59 ^ 1'b0 ;
  assign n13836 = ( n13792 & ~n13820 ) | ( n13792 & n13835 ) | ( ~n13820 & n13835 ) ;
  assign n13837 = n13835 ^ n13820 ^ n13792 ;
  assign n13838 = x119 & n263 ;
  assign n13839 = ( x121 & n264 ) | ( x121 & n13838 ) | ( n264 & n13838 ) ;
  assign n13840 = n13838 | n13839 ;
  assign n13841 = x120 & ~n260 ;
  assign n13842 = ( x120 & n13840 ) | ( x120 & ~n13841 ) | ( n13840 & ~n13841 ) ;
  assign n13843 = n272 & n9808 ;
  assign n13844 = n13842 | n13843 ;
  assign n13845 = n13844 ^ x56 ^ 1'b0 ;
  assign n13846 = ( n13802 & ~n13837 ) | ( n13802 & n13845 ) | ( ~n13837 & n13845 ) ;
  assign n13847 = n13845 ^ n13837 ^ n13802 ;
  assign n13848 = x115 & n208 ;
  assign n13849 = ( x117 & n194 ) | ( x117 & n13848 ) | ( n194 & n13848 ) ;
  assign n13850 = n13848 | n13849 ;
  assign n13851 = x116 & ~n192 ;
  assign n13852 = ( x116 & n13850 ) | ( x116 & ~n13851 ) | ( n13850 & ~n13851 ) ;
  assign n13853 = x122 & n408 ;
  assign n13854 = n13749 ^ x62 ^ 1'b0 ;
  assign n13855 = n197 & n9569 ;
  assign n13856 = n13852 | n13855 ;
  assign n13857 = n13856 ^ x62 ^ 1'b0 ;
  assign n13858 = ( x124 & n403 ) | ( x124 & n13853 ) | ( n403 & n13853 ) ;
  assign n13859 = n13853 | n13858 ;
  assign n13860 = x123 & ~n410 ;
  assign n13861 = ( x123 & n13859 ) | ( x123 & ~n13860 ) | ( n13859 & ~n13860 ) ;
  assign n13862 = n402 & n9858 ;
  assign n13863 = n13861 | n13862 ;
  assign n13864 = n13863 ^ x53 ^ 1'b0 ;
  assign n13865 = n13864 ^ n13847 ^ n13813 ;
  assign n13866 = ( n13813 & ~n13847 ) | ( n13813 & n13864 ) | ( ~n13847 & n13864 ) ;
  assign n13867 = n13771 ^ x50 ^ 1'b0 ;
  assign n13868 = n13867 ^ n13865 ^ n13823 ;
  assign n13869 = n13868 ^ n13827 ^ n13824 ;
  assign n13870 = ( ~n13824 & n13827 ) | ( ~n13824 & n13868 ) | ( n13827 & n13868 ) ;
  assign n13871 = ( n13823 & ~n13865 ) | ( n13823 & n13867 ) | ( ~n13865 & n13867 ) ;
  assign n13872 = x117 & n133 ;
  assign n13873 = ( x119 & n142 ) | ( x119 & n13872 ) | ( n142 & n13872 ) ;
  assign n13874 = n13872 | n13873 ;
  assign n13875 = x113 & ~n242 ;
  assign n13876 = x118 & ~n134 ;
  assign n13877 = ( x118 & n13874 ) | ( x118 & ~n13876 ) | ( n13874 & ~n13876 ) ;
  assign n13878 = x112 & n325 ;
  assign n13879 = ( x113 & ~n13875 ) | ( x113 & n13878 ) | ( ~n13875 & n13878 ) ;
  assign n13880 = n140 & n9733 ;
  assign n13881 = n13877 | n13880 ;
  assign n13882 = n13879 ^ n13854 ^ n13818 ;
  assign n13883 = n13768 ^ x50 ^ 1'b0 ;
  assign n13884 = n13881 ^ x59 ^ 1'b0 ;
  assign n13885 = ( n13818 & n13854 ) | ( n13818 & ~n13879 ) | ( n13854 & ~n13879 ) ;
  assign n13886 = ( n13821 & ~n13882 ) | ( n13821 & n13884 ) | ( ~n13882 & n13884 ) ;
  assign n13887 = n13884 ^ n13882 ^ n13821 ;
  assign n13888 = x120 & n263 ;
  assign n13889 = ( x122 & n264 ) | ( x122 & n13888 ) | ( n264 & n13888 ) ;
  assign n13890 = n13888 | n13889 ;
  assign n13891 = x121 & ~n260 ;
  assign n13892 = ( x121 & n13890 ) | ( x121 & ~n13891 ) | ( n13890 & ~n13891 ) ;
  assign n13893 = n272 & n9806 ;
  assign n13894 = n13892 | n13893 ;
  assign n13895 = n13894 ^ x56 ^ 1'b0 ;
  assign n13896 = n13895 ^ n13887 ^ n13836 ;
  assign n13897 = ( n13836 & ~n13887 ) | ( n13836 & n13895 ) | ( ~n13887 & n13895 ) ;
  assign n13898 = x123 & n408 ;
  assign n13899 = ( x125 & n403 ) | ( x125 & n13898 ) | ( n403 & n13898 ) ;
  assign n13900 = n13898 | n13899 ;
  assign n13901 = x124 & ~n410 ;
  assign n13902 = ( x124 & n13900 ) | ( x124 & ~n13901 ) | ( n13900 & ~n13901 ) ;
  assign n13903 = n402 & n9883 ;
  assign n13904 = n13902 | n13903 ;
  assign n13905 = n13904 ^ x53 ^ 1'b0 ;
  assign n13906 = n13905 ^ n13896 ^ n13846 ;
  assign n13907 = ( n13846 & ~n13896 ) | ( n13846 & n13905 ) | ( ~n13896 & n13905 ) ;
  assign n13908 = x127 & n408 ;
  assign n13909 = ( n402 & n9968 ) | ( n402 & n13908 ) | ( n9968 & n13908 ) ;
  assign n13910 = n13908 | n13909 ;
  assign n13911 = n13766 ^ x50 ^ 1'b0 ;
  assign n13912 = n13911 ^ n13906 ^ n13866 ;
  assign n13913 = ( n13866 & ~n13906 ) | ( n13866 & n13911 ) | ( ~n13906 & n13911 ) ;
  assign n13914 = ( n13870 & ~n13871 ) | ( n13870 & n13912 ) | ( ~n13871 & n13912 ) ;
  assign n13915 = n13912 ^ n13871 ^ n13870 ;
  assign n13916 = x125 & n408 ;
  assign n13917 = ( x127 & n403 ) | ( x127 & n13916 ) | ( n403 & n13916 ) ;
  assign n13918 = n13916 | n13917 ;
  assign n13919 = x124 & n408 ;
  assign n13920 = ( x126 & n403 ) | ( x126 & n13919 ) | ( n403 & n13919 ) ;
  assign n13921 = n13919 | n13920 ;
  assign n13922 = x126 & ~n410 ;
  assign n13923 = ( x126 & n13918 ) | ( x126 & ~n13922 ) | ( n13918 & ~n13922 ) ;
  assign n13924 = x125 & ~n410 ;
  assign n13925 = x127 & ~n410 ;
  assign n13926 = x126 & n408 ;
  assign n13927 = ( x127 & ~n13925 ) | ( x127 & n13926 ) | ( ~n13925 & n13926 ) ;
  assign n13928 = ( n402 & n9958 ) | ( n402 & n13926 ) | ( n9958 & n13926 ) ;
  assign n13929 = ( x125 & n13921 ) | ( x125 & ~n13924 ) | ( n13921 & ~n13924 ) ;
  assign n13930 = n13927 | n13928 ;
  assign n13931 = n402 & n9949 ;
  assign n13932 = n13923 | n13931 ;
  assign n13933 = x118 & n133 ;
  assign n13934 = ( x120 & n142 ) | ( x120 & n13933 ) | ( n142 & n13933 ) ;
  assign n13935 = n13933 | n13934 ;
  assign n13936 = n402 & n9917 ;
  assign n13937 = n13929 | n13936 ;
  assign n13938 = n140 & n9756 ;
  assign n13939 = x119 & ~n134 ;
  assign n13940 = ( x119 & n13935 ) | ( x119 & ~n13939 ) | ( n13935 & ~n13939 ) ;
  assign n13941 = n13938 | n13940 ;
  assign n13942 = x114 & ~n242 ;
  assign n13943 = x113 & n325 ;
  assign n13944 = ( x114 & ~n13942 ) | ( x114 & n13943 ) | ( ~n13942 & n13943 ) ;
  assign n13945 = n13944 ^ n13879 ^ n13857 ;
  assign n13946 = ( n13857 & ~n13879 ) | ( n13857 & n13944 ) | ( ~n13879 & n13944 ) ;
  assign n13947 = n13941 ^ x59 ^ 1'b0 ;
  assign n13948 = ( n13885 & ~n13945 ) | ( n13885 & n13947 ) | ( ~n13945 & n13947 ) ;
  assign n13949 = n13937 ^ x53 ^ 1'b0 ;
  assign n13950 = n13947 ^ n13945 ^ n13885 ;
  assign n13951 = x121 & n263 ;
  assign n13952 = ( x123 & n264 ) | ( x123 & n13951 ) | ( n264 & n13951 ) ;
  assign n13953 = n13951 | n13952 ;
  assign n13954 = x122 & ~n260 ;
  assign n13955 = ( x122 & n13953 ) | ( x122 & ~n13954 ) | ( n13953 & ~n13954 ) ;
  assign n13956 = n272 & n9828 ;
  assign n13957 = n13955 | n13956 ;
  assign n13958 = n13957 ^ x56 ^ 1'b0 ;
  assign n13959 = ( n13886 & ~n13950 ) | ( n13886 & n13958 ) | ( ~n13950 & n13958 ) ;
  assign n13960 = n13958 ^ n13950 ^ n13886 ;
  assign n13961 = n13960 ^ n13949 ^ n13897 ;
  assign n13962 = n13961 ^ n13907 ^ n13883 ;
  assign n13963 = ( n13883 & n13907 ) | ( n13883 & ~n13961 ) | ( n13907 & ~n13961 ) ;
  assign n13964 = n13962 ^ n13914 ^ n13913 ;
  assign n13965 = ( ~n13913 & n13914 ) | ( ~n13913 & n13962 ) | ( n13914 & n13962 ) ;
  assign n13966 = ( n13897 & n13949 ) | ( n13897 & ~n13960 ) | ( n13949 & ~n13960 ) ;
  assign n13967 = n197 & n9671 ;
  assign n13968 = x116 & n208 ;
  assign n13969 = ( x118 & n194 ) | ( x118 & n13968 ) | ( n194 & n13968 ) ;
  assign n13970 = n13968 | n13969 ;
  assign n13971 = x117 & ~n192 ;
  assign n13972 = ( x117 & n13970 ) | ( x117 & ~n13971 ) | ( n13970 & ~n13971 ) ;
  assign n13973 = n13967 | n13972 ;
  assign n13974 = x114 & n325 ;
  assign n13975 = x115 & ~n242 ;
  assign n13976 = ( x115 & n13974 ) | ( x115 & ~n13975 ) | ( n13974 & ~n13975 ) ;
  assign n13977 = n13973 ^ x62 ^ 1'b0 ;
  assign n13978 = n13976 ^ n13879 ^ x50 ;
  assign n13979 = ( ~x50 & n13879 ) | ( ~x50 & n13976 ) | ( n13879 & n13976 ) ;
  assign n13980 = n13978 ^ n13977 ^ n13946 ;
  assign n13981 = ( n13946 & n13977 ) | ( n13946 & ~n13978 ) | ( n13977 & ~n13978 ) ;
  assign n13982 = x119 & n133 ;
  assign n13983 = ( x121 & n142 ) | ( x121 & n13982 ) | ( n142 & n13982 ) ;
  assign n13984 = n13982 | n13983 ;
  assign n13985 = x120 & ~n134 ;
  assign n13986 = ( x120 & n13984 ) | ( x120 & ~n13985 ) | ( n13984 & ~n13985 ) ;
  assign n13987 = n140 & n9808 ;
  assign n13988 = n13986 | n13987 ;
  assign n13989 = n13988 ^ x59 ^ 1'b0 ;
  assign n13990 = ( n13948 & ~n13980 ) | ( n13948 & n13989 ) | ( ~n13980 & n13989 ) ;
  assign n13991 = n13989 ^ n13980 ^ n13948 ;
  assign n13992 = x122 & n263 ;
  assign n13993 = ( x124 & n264 ) | ( x124 & n13992 ) | ( n264 & n13992 ) ;
  assign n13994 = n13992 | n13993 ;
  assign n13995 = n197 & n9808 ;
  assign n13996 = x123 & ~n260 ;
  assign n13997 = ( x123 & n13994 ) | ( x123 & ~n13996 ) | ( n13994 & ~n13996 ) ;
  assign n13998 = n272 & n9858 ;
  assign n13999 = n13997 | n13998 ;
  assign n14000 = n13999 ^ x56 ^ 1'b0 ;
  assign n14001 = n14000 ^ n13991 ^ n13959 ;
  assign n14002 = n13932 ^ x53 ^ 1'b0 ;
  assign n14003 = ( n13959 & ~n13991 ) | ( n13959 & n14000 ) | ( ~n13991 & n14000 ) ;
  assign n14004 = n14002 ^ n14001 ^ n13966 ;
  assign n14005 = ( ~n13963 & n13965 ) | ( ~n13963 & n14004 ) | ( n13965 & n14004 ) ;
  assign n14006 = n14004 ^ n13965 ^ n13963 ;
  assign n14007 = ( n13966 & ~n14001 ) | ( n13966 & n14002 ) | ( ~n14001 & n14002 ) ;
  assign n14008 = x121 & ~n134 ;
  assign n14009 = x120 & n133 ;
  assign n14010 = ( x122 & n142 ) | ( x122 & n14009 ) | ( n142 & n14009 ) ;
  assign n14011 = n14009 | n14010 ;
  assign n14012 = ( x121 & ~n14008 ) | ( x121 & n14011 ) | ( ~n14008 & n14011 ) ;
  assign n14013 = x117 & n208 ;
  assign n14014 = n197 & n9733 ;
  assign n14015 = ( x119 & n194 ) | ( x119 & n14013 ) | ( n194 & n14013 ) ;
  assign n14016 = n14013 | n14015 ;
  assign n14017 = x118 & ~n192 ;
  assign n14018 = ( x118 & n14016 ) | ( x118 & ~n14017 ) | ( n14016 & ~n14017 ) ;
  assign n14019 = x115 & n325 ;
  assign n14020 = n14014 | n14018 ;
  assign n14021 = x116 & ~n242 ;
  assign n14022 = ( x116 & n14019 ) | ( x116 & ~n14021 ) | ( n14019 & ~n14021 ) ;
  assign n14023 = n14020 ^ x62 ^ 1'b0 ;
  assign n14024 = n14023 ^ n14022 ^ n13979 ;
  assign n14025 = ( n13979 & ~n14022 ) | ( n13979 & n14023 ) | ( ~n14022 & n14023 ) ;
  assign n14026 = n140 & n9806 ;
  assign n14027 = n14012 | n14026 ;
  assign n14028 = n14027 ^ x59 ^ 1'b0 ;
  assign n14029 = ( n13981 & ~n14024 ) | ( n13981 & n14028 ) | ( ~n14024 & n14028 ) ;
  assign n14030 = n13910 ^ x53 ^ 1'b0 ;
  assign n14031 = n14028 ^ n14024 ^ n13981 ;
  assign n14032 = x123 & n263 ;
  assign n14033 = n13930 ^ x53 ^ 1'b0 ;
  assign n14034 = ( x125 & n264 ) | ( x125 & n14032 ) | ( n264 & n14032 ) ;
  assign n14035 = n197 & n9756 ;
  assign n14036 = n14032 | n14034 ;
  assign n14037 = x124 & ~n260 ;
  assign n14038 = ( x124 & n14036 ) | ( x124 & ~n14037 ) | ( n14036 & ~n14037 ) ;
  assign n14039 = n272 & n9883 ;
  assign n14040 = n14038 | n14039 ;
  assign n14041 = n14040 ^ x56 ^ 1'b0 ;
  assign n14042 = n14041 ^ n14031 ^ n13990 ;
  assign n14043 = ( n13990 & ~n14031 ) | ( n13990 & n14041 ) | ( ~n14031 & n14041 ) ;
  assign n14044 = ( n14003 & n14033 ) | ( n14003 & ~n14042 ) | ( n14033 & ~n14042 ) ;
  assign n14045 = n14042 ^ n14033 ^ n14003 ;
  assign n14046 = n14045 ^ n14007 ^ n14005 ;
  assign n14047 = ( n14005 & ~n14007 ) | ( n14005 & n14045 ) | ( ~n14007 & n14045 ) ;
  assign n14048 = x118 & n208 ;
  assign n14049 = ( x120 & n194 ) | ( x120 & n14048 ) | ( n194 & n14048 ) ;
  assign n14050 = x119 & ~n192 ;
  assign n14051 = n14048 | n14049 ;
  assign n14052 = ( x119 & ~n14050 ) | ( x119 & n14051 ) | ( ~n14050 & n14051 ) ;
  assign n14053 = n14035 | n14052 ;
  assign n14054 = x117 & ~n242 ;
  assign n14055 = x121 & n133 ;
  assign n14056 = ( x123 & n142 ) | ( x123 & n14055 ) | ( n142 & n14055 ) ;
  assign n14057 = n14055 | n14056 ;
  assign n14058 = x122 & ~n134 ;
  assign n14059 = ( x122 & n14057 ) | ( x122 & ~n14058 ) | ( n14057 & ~n14058 ) ;
  assign n14060 = n140 & n9828 ;
  assign n14061 = n14059 | n14060 ;
  assign n14062 = x116 & n325 ;
  assign n14063 = ( x117 & ~n14054 ) | ( x117 & n14062 ) | ( ~n14054 & n14062 ) ;
  assign n14064 = n14053 ^ x62 ^ 1'b0 ;
  assign n14065 = n14063 ^ n14025 ^ n14022 ;
  assign n14066 = ( n14022 & n14025 ) | ( n14022 & ~n14063 ) | ( n14025 & ~n14063 ) ;
  assign n14067 = n14061 ^ x59 ^ 1'b0 ;
  assign n14068 = n14067 ^ n14065 ^ n14064 ;
  assign n14069 = ( n14064 & ~n14065 ) | ( n14064 & n14067 ) | ( ~n14065 & n14067 ) ;
  assign n14070 = x124 & n263 ;
  assign n14071 = ( x126 & n264 ) | ( x126 & n14070 ) | ( n264 & n14070 ) ;
  assign n14072 = n14070 | n14071 ;
  assign n14073 = x125 & ~n260 ;
  assign n14074 = ( x125 & n14072 ) | ( x125 & ~n14073 ) | ( n14072 & ~n14073 ) ;
  assign n14075 = n272 & n9917 ;
  assign n14076 = n14074 | n14075 ;
  assign n14077 = n14076 ^ x56 ^ 1'b0 ;
  assign n14078 = n14077 ^ n14068 ^ n14029 ;
  assign n14079 = ( n14029 & ~n14068 ) | ( n14029 & n14077 ) | ( ~n14068 & n14077 ) ;
  assign n14080 = ( n14030 & n14043 ) | ( n14030 & ~n14078 ) | ( n14043 & ~n14078 ) ;
  assign n14081 = n14078 ^ n14043 ^ n14030 ;
  assign n14082 = x119 & n208 ;
  assign n14083 = x125 & n263 ;
  assign n14084 = ( x121 & n194 ) | ( x121 & n14082 ) | ( n194 & n14082 ) ;
  assign n14085 = n14082 | n14084 ;
  assign n14086 = x120 & ~n192 ;
  assign n14087 = ( x120 & n14085 ) | ( x120 & ~n14086 ) | ( n14085 & ~n14086 ) ;
  assign n14088 = n13995 | n14087 ;
  assign n14089 = ( x127 & n264 ) | ( x127 & n14083 ) | ( n264 & n14083 ) ;
  assign n14090 = x118 & ~n242 ;
  assign n14091 = x117 & n325 ;
  assign n14092 = n14083 | n14089 ;
  assign n14093 = n14081 ^ n14047 ^ n14044 ;
  assign n14094 = ( ~n14044 & n14047 ) | ( ~n14044 & n14081 ) | ( n14047 & n14081 ) ;
  assign n14095 = n272 & n9949 ;
  assign n14096 = x126 & ~n260 ;
  assign n14097 = ( x126 & n14092 ) | ( x126 & ~n14096 ) | ( n14092 & ~n14096 ) ;
  assign n14098 = x127 & n263 ;
  assign n14099 = x126 & n263 ;
  assign n14100 = n14095 | n14097 ;
  assign n14101 = ( n272 & n9958 ) | ( n272 & n14099 ) | ( n9958 & n14099 ) ;
  assign n14102 = ( x118 & ~n14090 ) | ( x118 & n14091 ) | ( ~n14090 & n14091 ) ;
  assign n14103 = n140 & n9858 ;
  assign n14104 = n14088 ^ x62 ^ 1'b0 ;
  assign n14105 = x127 & ~n260 ;
  assign n14106 = ( x127 & n14099 ) | ( x127 & ~n14105 ) | ( n14099 & ~n14105 ) ;
  assign n14107 = ( ~x53 & n14063 ) | ( ~x53 & n14102 ) | ( n14063 & n14102 ) ;
  assign n14108 = n14102 ^ n14063 ^ x53 ;
  assign n14109 = x123 & ~n134 ;
  assign n14110 = n14101 | n14106 ;
  assign n14111 = ( n272 & n9968 ) | ( n272 & n14098 ) | ( n9968 & n14098 ) ;
  assign n14112 = ( n14066 & n14104 ) | ( n14066 & ~n14108 ) | ( n14104 & ~n14108 ) ;
  assign n14113 = n14100 ^ x56 ^ 1'b0 ;
  assign n14114 = n14108 ^ n14104 ^ n14066 ;
  assign n14115 = x122 & n133 ;
  assign n14116 = ( x124 & n142 ) | ( x124 & n14115 ) | ( n142 & n14115 ) ;
  assign n14117 = n14098 | n14111 ;
  assign n14118 = n14115 | n14116 ;
  assign n14119 = ( x123 & ~n14109 ) | ( x123 & n14118 ) | ( ~n14109 & n14118 ) ;
  assign n14120 = n14103 | n14119 ;
  assign n14121 = n14120 ^ x59 ^ 1'b0 ;
  assign n14122 = n14121 ^ n14114 ^ n14069 ;
  assign n14123 = ( n14069 & ~n14114 ) | ( n14069 & n14121 ) | ( ~n14114 & n14121 ) ;
  assign n14124 = n14122 ^ n14113 ^ n14079 ;
  assign n14125 = ( ~n14080 & n14094 ) | ( ~n14080 & n14124 ) | ( n14094 & n14124 ) ;
  assign n14126 = ( n14079 & n14113 ) | ( n14079 & ~n14122 ) | ( n14113 & ~n14122 ) ;
  assign n14127 = n14124 ^ n14094 ^ n14080 ;
  assign n14128 = x122 & n208 ;
  assign n14129 = x121 & n208 ;
  assign n14130 = n197 & n9828 ;
  assign n14131 = ( x123 & n194 ) | ( x123 & n14129 ) | ( n194 & n14129 ) ;
  assign n14132 = n14129 | n14131 ;
  assign n14133 = x122 & ~n192 ;
  assign n14134 = ( x122 & n14132 ) | ( x122 & ~n14133 ) | ( n14132 & ~n14133 ) ;
  assign n14135 = ( x124 & n194 ) | ( x124 & n14128 ) | ( n194 & n14128 ) ;
  assign n14136 = n14130 | n14134 ;
  assign n14137 = n14128 | n14135 ;
  assign n14138 = x123 & ~n192 ;
  assign n14139 = ( x123 & n14137 ) | ( x123 & ~n14138 ) | ( n14137 & ~n14138 ) ;
  assign n14140 = x123 & n133 ;
  assign n14141 = ( x125 & n142 ) | ( x125 & n14140 ) | ( n142 & n14140 ) ;
  assign n14142 = n14140 | n14141 ;
  assign n14143 = x124 & ~n134 ;
  assign n14144 = ( x124 & n14142 ) | ( x124 & ~n14143 ) | ( n14142 & ~n14143 ) ;
  assign n14145 = n140 & n9883 ;
  assign n14146 = n14144 | n14145 ;
  assign n14147 = x120 & n208 ;
  assign n14148 = n197 & n9858 ;
  assign n14149 = n14139 | n14148 ;
  assign n14150 = ( x122 & n194 ) | ( x122 & n14147 ) | ( n194 & n14147 ) ;
  assign n14151 = n14147 | n14150 ;
  assign n14152 = x121 & ~n192 ;
  assign n14153 = ( x121 & n14151 ) | ( x121 & ~n14152 ) | ( n14151 & ~n14152 ) ;
  assign n14154 = x119 & ~n242 ;
  assign n14155 = n14146 ^ x59 ^ 1'b0 ;
  assign n14156 = n14110 ^ x56 ^ 1'b0 ;
  assign n14157 = ( n197 & n9806 ) | ( n197 & n14153 ) | ( n9806 & n14153 ) ;
  assign n14158 = n14153 | n14157 ;
  assign n14159 = x118 & n325 ;
  assign n14160 = ( x119 & ~n14154 ) | ( x119 & n14159 ) | ( ~n14154 & n14159 ) ;
  assign n14161 = n14158 ^ x62 ^ 1'b0 ;
  assign n14162 = n14161 ^ n14160 ^ n14107 ;
  assign n14163 = ( n14107 & ~n14160 ) | ( n14107 & n14161 ) | ( ~n14160 & n14161 ) ;
  assign n14164 = ( n14112 & n14155 ) | ( n14112 & ~n14162 ) | ( n14155 & ~n14162 ) ;
  assign n14165 = n14162 ^ n14155 ^ n14112 ;
  assign n14166 = n14165 ^ n14156 ^ n14123 ;
  assign n14167 = ( n14123 & n14156 ) | ( n14123 & ~n14165 ) | ( n14156 & ~n14165 ) ;
  assign n14168 = n14166 ^ n14126 ^ n14125 ;
  assign n14169 = ( n14125 & ~n14126 ) | ( n14125 & n14166 ) | ( ~n14126 & n14166 ) ;
  assign n14170 = x124 & n133 ;
  assign n14171 = ( x126 & n142 ) | ( x126 & n14170 ) | ( n142 & n14170 ) ;
  assign n14172 = n14170 | n14171 ;
  assign n14173 = x125 & n133 ;
  assign n14174 = ( x127 & n142 ) | ( x127 & n14173 ) | ( n142 & n14173 ) ;
  assign n14175 = n14173 | n14174 ;
  assign n14176 = x126 & ~n134 ;
  assign n14177 = ( x126 & n14175 ) | ( x126 & ~n14176 ) | ( n14175 & ~n14176 ) ;
  assign n14178 = n140 & n9949 ;
  assign n14179 = n14177 | n14178 ;
  assign n14180 = x125 & ~n134 ;
  assign n14181 = ( x125 & n14172 ) | ( x125 & ~n14180 ) | ( n14172 & ~n14180 ) ;
  assign n14182 = x126 & n133 ;
  assign n14183 = x127 & ~n134 ;
  assign n14184 = ( x127 & n14182 ) | ( x127 & ~n14183 ) | ( n14182 & ~n14183 ) ;
  assign n14185 = ( n140 & n9958 ) | ( n140 & n14182 ) | ( n9958 & n14182 ) ;
  assign n14186 = n14149 ^ x62 ^ 1'b0 ;
  assign n14187 = n14184 | n14185 ;
  assign n14188 = n140 & n9917 ;
  assign n14189 = x127 & n133 ;
  assign n14190 = ( n140 & n9968 ) | ( n140 & n14189 ) | ( n9968 & n14189 ) ;
  assign n14191 = n14136 ^ x62 ^ 1'b0 ;
  assign n14192 = n14181 | n14188 ;
  assign n14193 = n14192 ^ x59 ^ 1'b0 ;
  assign n14194 = n14189 | n14190 ;
  assign n14195 = x119 & n325 ;
  assign n14196 = x120 & ~n242 ;
  assign n14197 = ( x120 & n14195 ) | ( x120 & ~n14196 ) | ( n14195 & ~n14196 ) ;
  assign n14198 = ( ~n14160 & n14191 ) | ( ~n14160 & n14197 ) | ( n14191 & n14197 ) ;
  assign n14199 = n14197 ^ n14191 ^ n14160 ;
  assign n14200 = ( n14163 & n14193 ) | ( n14163 & ~n14199 ) | ( n14193 & ~n14199 ) ;
  assign n14201 = n14199 ^ n14193 ^ n14163 ;
  assign n14202 = n14117 ^ x56 ^ 1'b0 ;
  assign n14203 = x121 & ~n242 ;
  assign n14204 = x120 & n325 ;
  assign n14205 = ( x121 & ~n14203 ) | ( x121 & n14204 ) | ( ~n14203 & n14204 ) ;
  assign n14206 = n14205 ^ n14160 ^ x56 ;
  assign n14207 = n14179 ^ x59 ^ 1'b0 ;
  assign n14208 = ( ~x56 & n14160 ) | ( ~x56 & n14205 ) | ( n14160 & n14205 ) ;
  assign n14209 = ( n14186 & n14198 ) | ( n14186 & ~n14206 ) | ( n14198 & ~n14206 ) ;
  assign n14210 = n14206 ^ n14198 ^ n14186 ;
  assign n14211 = n14202 ^ n14201 ^ n14164 ;
  assign n14212 = n14210 ^ n14207 ^ n14200 ;
  assign n14213 = ( n14200 & n14207 ) | ( n14200 & ~n14210 ) | ( n14207 & ~n14210 ) ;
  assign n14214 = ( ~n14167 & n14169 ) | ( ~n14167 & n14211 ) | ( n14169 & n14211 ) ;
  assign n14215 = n14211 ^ n14169 ^ n14167 ;
  assign n14216 = ( n14164 & ~n14201 ) | ( n14164 & n14202 ) | ( ~n14201 & n14202 ) ;
  assign n14217 = ( n14212 & n14214 ) | ( n14212 & ~n14216 ) | ( n14214 & ~n14216 ) ;
  assign n14218 = n14216 ^ n14214 ^ n14212 ;
  assign n14219 = x124 & n208 ;
  assign n14220 = ( x126 & n194 ) | ( x126 & n14219 ) | ( n194 & n14219 ) ;
  assign n14221 = n14219 | n14220 ;
  assign n14222 = x125 & ~n192 ;
  assign n14223 = ( x125 & n14221 ) | ( x125 & ~n14222 ) | ( n14221 & ~n14222 ) ;
  assign n14224 = n197 & n9917 ;
  assign n14225 = n14223 | n14224 ;
  assign n14226 = x125 & n208 ;
  assign n14227 = ( x127 & n194 ) | ( x127 & n14226 ) | ( n194 & n14226 ) ;
  assign n14228 = n14226 | n14227 ;
  assign n14229 = x126 & ~n192 ;
  assign n14230 = n197 & n9949 ;
  assign n14231 = ( x126 & n14228 ) | ( x126 & ~n14229 ) | ( n14228 & ~n14229 ) ;
  assign n14232 = x123 & n208 ;
  assign n14233 = ( x125 & n194 ) | ( x125 & n14232 ) | ( n194 & n14232 ) ;
  assign n14234 = n14232 | n14233 ;
  assign n14235 = x124 & ~n192 ;
  assign n14236 = x127 & ~n192 ;
  assign n14237 = ( x124 & n14234 ) | ( x124 & ~n14235 ) | ( n14234 & ~n14235 ) ;
  assign n14238 = x127 & n208 ;
  assign n14239 = ( n197 & n9968 ) | ( n197 & n14238 ) | ( n9968 & n14238 ) ;
  assign n14240 = x126 & n208 ;
  assign n14241 = ( n197 & n9958 ) | ( n197 & n14240 ) | ( n9958 & n14240 ) ;
  assign n14242 = ( x127 & ~n14236 ) | ( x127 & n14240 ) | ( ~n14236 & n14240 ) ;
  assign n14243 = x121 & n325 ;
  assign n14244 = n14238 | n14239 ;
  assign n14245 = x122 & ~n242 ;
  assign n14246 = n14187 ^ x59 ^ 1'b0 ;
  assign n14247 = ( n197 & n9883 ) | ( n197 & n14237 ) | ( n9883 & n14237 ) ;
  assign n14248 = n14237 | n14247 ;
  assign n14249 = n14248 ^ x62 ^ 1'b0 ;
  assign n14250 = n14241 | n14242 ;
  assign n14251 = ( x122 & n14243 ) | ( x122 & ~n14245 ) | ( n14243 & ~n14245 ) ;
  assign n14252 = n14251 ^ n14249 ^ n14208 ;
  assign n14253 = n14252 ^ n14246 ^ n14209 ;
  assign n14254 = ( ~n14213 & n14217 ) | ( ~n14213 & n14253 ) | ( n14217 & n14253 ) ;
  assign n14255 = ( n14208 & n14249 ) | ( n14208 & ~n14251 ) | ( n14249 & ~n14251 ) ;
  assign n14256 = n14253 ^ n14217 ^ n14213 ;
  assign n14257 = ( n14209 & n14246 ) | ( n14209 & ~n14252 ) | ( n14246 & ~n14252 ) ;
  assign n14258 = n14230 | n14231 ;
  assign n14259 = x123 & ~n242 ;
  assign n14260 = x122 & n325 ;
  assign n14261 = ( x123 & ~n14259 ) | ( x123 & n14260 ) | ( ~n14259 & n14260 ) ;
  assign n14262 = n14225 ^ x62 ^ 1'b0 ;
  assign n14263 = ( n14251 & n14255 ) | ( n14251 & ~n14261 ) | ( n14255 & ~n14261 ) ;
  assign n14264 = n14261 ^ n14255 ^ n14251 ;
  assign n14265 = n14194 ^ x59 ^ 1'b0 ;
  assign n14266 = n14265 ^ n14264 ^ n14262 ;
  assign n14267 = ( n14262 & ~n14264 ) | ( n14262 & n14265 ) | ( ~n14264 & n14265 ) ;
  assign n14268 = n14258 ^ x62 ^ 1'b0 ;
  assign n14269 = x123 & n325 ;
  assign n14270 = n14250 ^ x62 ^ 1'b0 ;
  assign n14271 = x124 & ~n242 ;
  assign n14272 = ( x124 & n14269 ) | ( x124 & ~n14271 ) | ( n14269 & ~n14271 ) ;
  assign n14273 = ( n14254 & ~n14257 ) | ( n14254 & n14266 ) | ( ~n14257 & n14266 ) ;
  assign n14274 = n14266 ^ n14257 ^ n14254 ;
  assign n14275 = n14272 ^ n14261 ^ x59 ;
  assign n14276 = n14275 ^ n14268 ^ n14263 ;
  assign n14277 = ( n14263 & n14268 ) | ( n14263 & ~n14275 ) | ( n14268 & ~n14275 ) ;
  assign n14278 = x125 & ~n242 ;
  assign n14279 = x126 & ~n242 ;
  assign n14280 = ( ~x59 & n14261 ) | ( ~x59 & n14272 ) | ( n14261 & n14272 ) ;
  assign n14281 = x124 & n325 ;
  assign n14282 = ( x125 & ~n14278 ) | ( x125 & n14281 ) | ( ~n14278 & n14281 ) ;
  assign n14283 = x125 & n325 ;
  assign n14284 = n14244 ^ x62 ^ 1'b0 ;
  assign n14285 = ( x126 & ~n14279 ) | ( x126 & n14283 ) | ( ~n14279 & n14283 ) ;
  assign n14286 = x126 & n325 ;
  assign n14287 = x127 & n325 ;
  assign n14288 = x127 & ~n242 ;
  assign n14289 = ( x127 & n14286 ) | ( x127 & ~n14288 ) | ( n14286 & ~n14288 ) ;
  assign n14290 = n14276 ^ n14273 ^ n14267 ;
  assign n14291 = ( ~n14267 & n14273 ) | ( ~n14267 & n14276 ) | ( n14273 & n14276 ) ;
  assign n14292 = n14285 ^ n14284 ^ n14282 ;
  assign n14293 = ( ~n14282 & n14284 ) | ( ~n14282 & n14285 ) | ( n14284 & n14285 ) ;
  assign n14294 = n14282 ^ n14280 ^ n14270 ;
  assign n14295 = n14294 ^ n14291 ^ n14277 ;
  assign n14296 = ( n14270 & n14280 ) | ( n14270 & ~n14282 ) | ( n14280 & ~n14282 ) ;
  assign n14297 = n14289 ^ n14282 ^ x62 ;
  assign n14298 = ( ~x62 & n14282 ) | ( ~x62 & n14289 ) | ( n14282 & n14289 ) ;
  assign n14299 = ( ~n14277 & n14291 ) | ( ~n14277 & n14294 ) | ( n14291 & n14294 ) ;
  assign n14300 = n14299 ^ n14296 ^ n14292 ;
  assign n14301 = ( n14292 & ~n14296 ) | ( n14292 & n14299 ) | ( ~n14296 & n14299 ) ;
  assign n14302 = ( ~n14293 & n14297 ) | ( ~n14293 & n14301 ) | ( n14297 & n14301 ) ;
  assign n14303 = n14301 ^ n14297 ^ n14293 ;
  assign n14304 = n14302 ^ n14298 ^ n14287 ;
  assign y0 = n6170 ;
  assign y1 = n6172 ;
  assign y2 = n6188 ;
  assign y3 = n6175 ;
  assign y4 = n6179 ;
  assign y5 = n6178 ;
  assign y6 = n6183 ;
  assign y7 = n6182 ;
  assign y8 = n6186 ;
  assign y9 = n6220 ;
  assign y10 = n6223 ;
  assign y11 = n6234 ;
  assign y12 = n6254 ;
  assign y13 = n6238 ;
  assign y14 = n6252 ;
  assign y15 = n6266 ;
  assign y16 = n6290 ;
  assign y17 = n6326 ;
  assign y18 = n6398 ;
  assign y19 = n6407 ;
  assign y20 = n6417 ;
  assign y21 = n6428 ;
  assign y22 = n6437 ;
  assign y23 = n6448 ;
  assign y24 = n6457 ;
  assign y25 = n6468 ;
  assign y26 = n6477 ;
  assign y27 = n6488 ;
  assign y28 = n6507 ;
  assign y29 = n7109 ;
  assign y30 = n7307 ;
  assign y31 = n7326 ;
  assign y32 = n7337 ;
  assign y33 = n7346 ;
  assign y34 = n7357 ;
  assign y35 = n7367 ;
  assign y36 = n7416 ;
  assign y37 = n7426 ;
  assign y38 = n7477 ;
  assign y39 = n8006 ;
  assign y40 = n8049 ;
  assign y41 = n8120 ;
  assign y42 = n8403 ;
  assign y43 = n8475 ;
  assign y44 = n8575 ;
  assign y45 = n8700 ;
  assign y46 = n8931 ;
  assign y47 = n8986 ;
  assign y48 = n9115 ;
  assign y49 = n9216 ;
  assign y50 = n9511 ;
  assign y51 = n9531 ;
  assign y52 = n9562 ;
  assign y53 = n9574 ;
  assign y54 = n9706 ;
  assign y55 = n9755 ;
  assign y56 = n9761 ;
  assign y57 = n9822 ;
  assign y58 = n9826 ;
  assign y59 = n9846 ;
  assign y60 = n9881 ;
  assign y61 = n9890 ;
  assign y62 = n9929 ;
  assign y63 = n9963 ;
  assign y64 = n9989 ;
  assign y65 = n10036 ;
  assign y66 = n10073 ;
  assign y67 = n10096 ;
  assign y68 = n10148 ;
  assign y69 = n10152 ;
  assign y70 = n10206 ;
  assign y71 = n10286 ;
  assign y72 = n10293 ;
  assign y73 = n10340 ;
  assign y74 = n10404 ;
  assign y75 = n10431 ;
  assign y76 = n10501 ;
  assign y77 = n10541 ;
  assign y78 = n10563 ;
  assign y79 = n10638 ;
  assign y80 = n10651 ;
  assign y81 = n10702 ;
  assign y82 = n10849 ;
  assign y83 = n11005 ;
  assign y84 = n11169 ;
  assign y85 = n11301 ;
  assign y86 = n11451 ;
  assign y87 = n11574 ;
  assign y88 = n11694 ;
  assign y89 = n11846 ;
  assign y90 = n11975 ;
  assign y91 = n12083 ;
  assign y92 = n12208 ;
  assign y93 = n12335 ;
  assign y94 = n12440 ;
  assign y95 = n12556 ;
  assign y96 = n12649 ;
  assign y97 = n12784 ;
  assign y98 = n12886 ;
  assign y99 = n12952 ;
  assign y100 = n13039 ;
  assign y101 = n13140 ;
  assign y102 = n13243 ;
  assign y103 = n13335 ;
  assign y104 = n13401 ;
  assign y105 = n13474 ;
  assign y106 = n13555 ;
  assign y107 = n13615 ;
  assign y108 = n13676 ;
  assign y109 = n13732 ;
  assign y110 = n13826 ;
  assign y111 = n13869 ;
  assign y112 = n13915 ;
  assign y113 = n13964 ;
  assign y114 = n14006 ;
  assign y115 = n14046 ;
  assign y116 = n14093 ;
  assign y117 = n14127 ;
  assign y118 = n14168 ;
  assign y119 = n14215 ;
  assign y120 = n14218 ;
  assign y121 = n14256 ;
  assign y122 = n14274 ;
  assign y123 = n14290 ;
  assign y124 = n14295 ;
  assign y125 = n14300 ;
  assign y126 = n14303 ;
  assign y127 = n14304 ;
endmodule
