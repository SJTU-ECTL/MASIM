module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 ;
  assign n129 = x30 ^ x29 ^ 1'b0 ;
  assign n130 = x27 | x28 ;
  assign n131 = ~x29 & n130 ;
  assign n132 = x25 | x26 ;
  assign n133 = x23 | x24 ;
  assign n134 = ( x30 & ~n129 ) | ( x30 & n130 ) | ( ~n129 & n130 ) ;
  assign n135 = n134 ^ x27 ^ 1'b0 ;
  assign n136 = x29 | x30 ;
  assign n137 = n130 ^ x29 ^ 1'b0 ;
  assign n138 = x30 & ~n137 ;
  assign n139 = ( x28 & x30 ) | ( x28 & ~n129 ) | ( x30 & ~n129 ) ;
  assign n140 = x27 | n139 ;
  assign n141 = n140 ^ x28 ^ x27 ;
  assign n142 = ( n132 & ~n134 ) | ( n132 & n135 ) | ( ~n134 & n135 ) ;
  assign n143 = ( ~n136 & n141 ) | ( ~n136 & n142 ) | ( n141 & n142 ) ;
  assign n144 = n138 | n143 ;
  assign n145 = ( n142 & n143 ) | ( n142 & n144 ) | ( n143 & n144 ) ;
  assign n146 = ( ~x30 & n141 ) | ( ~x30 & n142 ) | ( n141 & n142 ) ;
  assign n147 = n141 & ~n145 ;
  assign n148 = n147 ^ n145 ^ n143 ;
  assign n149 = n141 & ~n142 ;
  assign n150 = n136 & n146 ;
  assign n151 = ( n138 & n141 ) | ( n138 & ~n149 ) | ( n141 & ~n149 ) ;
  assign n152 = ~n136 & n146 ;
  assign n153 = n144 ^ x25 ^ 1'b0 ;
  assign n154 = x25 | n144 ;
  assign n155 = n154 ^ x26 ^ x25 ;
  assign n156 = ~n132 & n144 ;
  assign n157 = ~n138 & n149 ;
  assign n158 = ( n131 & n134 ) | ( n131 & n157 ) | ( n134 & n157 ) ;
  assign n159 = ( n146 & ~n150 ) | ( n146 & n158 ) | ( ~n150 & n158 ) ;
  assign n160 = ( ~n152 & n156 ) | ( ~n152 & n159 ) | ( n156 & n159 ) ;
  assign n161 = ( n133 & ~n144 ) | ( n133 & n153 ) | ( ~n144 & n153 ) ;
  assign n162 = ( ~n134 & n155 ) | ( ~n134 & n161 ) | ( n155 & n161 ) ;
  assign n163 = n160 ^ x27 ^ 1'b0 ;
  assign n164 = ( n136 & n162 ) | ( n136 & n163 ) | ( n162 & n163 ) ;
  assign n165 = n141 & ~n144 ;
  assign n166 = n161 ^ n134 ^ 1'b0 ;
  assign n167 = ~n136 & n162 ;
  assign n168 = ( ~n141 & n144 ) | ( ~n141 & n163 ) | ( n144 & n163 ) ;
  assign n169 = ( n141 & n142 ) | ( n141 & n163 ) | ( n142 & n163 ) ;
  assign n170 = ( ~n136 & n167 ) | ( ~n136 & n169 ) | ( n167 & n169 ) ;
  assign n171 = ( n136 & n142 ) | ( n136 & ~n170 ) | ( n142 & ~n170 ) ;
  assign n172 = n162 & n163 ;
  assign n173 = ( n168 & n170 ) | ( n168 & ~n171 ) | ( n170 & ~n171 ) ;
  assign n174 = n148 | n173 ;
  assign n175 = ( n162 & n172 ) | ( n162 & ~n174 ) | ( n172 & ~n174 ) ;
  assign n176 = n164 & ~n175 ;
  assign n177 = ( n148 & n163 ) | ( n148 & ~n165 ) | ( n163 & ~n165 ) ;
  assign n178 = n162 & ~n172 ;
  assign n179 = n172 | n174 ;
  assign n180 = ( ~n163 & n172 ) | ( ~n163 & n179 ) | ( n172 & n179 ) ;
  assign n181 = ( n172 & ~n178 ) | ( n172 & n180 ) | ( ~n178 & n180 ) ;
  assign n182 = n144 & ~n172 ;
  assign n183 = n165 | n179 ;
  assign n184 = ~n133 & n179 ;
  assign n185 = ( n148 & n173 ) | ( n148 & ~n184 ) | ( n173 & ~n184 ) ;
  assign n186 = n182 | n184 ;
  assign n187 = ~n176 & n179 ;
  assign n188 = ( n176 & n177 ) | ( n176 & ~n187 ) | ( n177 & ~n187 ) ;
  assign n189 = ( n184 & ~n185 ) | ( n184 & n186 ) | ( ~n185 & n186 ) ;
  assign n190 = ( n155 & n176 ) | ( n155 & n179 ) | ( n176 & n179 ) ;
  assign n191 = ~x23 & n179 ;
  assign n192 = n191 ^ x24 ^ 1'b0 ;
  assign n193 = x20 | x21 ;
  assign n194 = ( x23 & n144 ) | ( x23 & ~n193 ) | ( n144 & ~n193 ) ;
  assign n195 = ( ~n166 & n188 ) | ( ~n166 & n190 ) | ( n188 & n190 ) ;
  assign n196 = ( x23 & n152 ) | ( x23 & n179 ) | ( n152 & n179 ) ;
  assign n197 = ( x23 & ~n151 ) | ( x23 & n193 ) | ( ~n151 & n193 ) ;
  assign n198 = ~n151 & n197 ;
  assign n199 = ( ~x23 & n144 ) | ( ~x23 & n179 ) | ( n144 & n179 ) ;
  assign n200 = ( ~n152 & n196 ) | ( ~n152 & n198 ) | ( n196 & n198 ) ;
  assign n201 = ~n196 & n200 ;
  assign n202 = ~n166 & n179 ;
  assign n203 = n192 | n201 ;
  assign n204 = n194 & n199 ;
  assign n205 = n203 & ~n204 ;
  assign n206 = n189 ^ x25 ^ 1'b0 ;
  assign n207 = n202 ^ n155 ^ 1'b0 ;
  assign n208 = ( ~n134 & n205 ) | ( ~n134 & n206 ) | ( n205 & n206 ) ;
  assign n209 = ( n155 & ~n188 ) | ( n155 & n202 ) | ( ~n188 & n202 ) ;
  assign n210 = n207 | n208 ;
  assign n211 = ( ~x30 & n181 ) | ( ~x30 & n210 ) | ( n181 & n210 ) ;
  assign n212 = n207 & n208 ;
  assign n213 = ~n136 & n211 ;
  assign n214 = ( ~n188 & n195 ) | ( ~n188 & n209 ) | ( n195 & n209 ) ;
  assign n215 = ~n195 & n214 ;
  assign n216 = n212 | n213 ;
  assign n217 = n188 | n216 ;
  assign n218 = ( ~n210 & n212 ) | ( ~n210 & n217 ) | ( n212 & n217 ) ;
  assign n219 = ( n201 & ~n204 ) | ( n201 & n217 ) | ( ~n204 & n217 ) ;
  assign n220 = ~n201 & n219 ;
  assign n221 = ( ~n212 & n213 ) | ( ~n212 & n215 ) | ( n213 & n215 ) ;
  assign n222 = n220 ^ n191 ^ x24 ;
  assign n223 = ( n136 & n207 ) | ( n136 & n208 ) | ( n207 & n208 ) ;
  assign n224 = ( n208 & n212 ) | ( n208 & ~n217 ) | ( n212 & ~n217 ) ;
  assign n225 = n223 & ~n224 ;
  assign n226 = n213 & n221 ;
  assign n227 = ~n193 & n217 ;
  assign n228 = ( n176 & n213 ) | ( n176 & ~n227 ) | ( n213 & ~n227 ) ;
  assign n229 = ( n221 & n225 ) | ( n221 & ~n226 ) | ( n225 & ~n226 ) ;
  assign n230 = n179 & ~n212 ;
  assign n231 = n134 & n205 ;
  assign n232 = n227 | n230 ;
  assign n233 = ( n213 & n217 ) | ( n213 & ~n229 ) | ( n217 & ~n229 ) ;
  assign n234 = ( n134 & ~n205 ) | ( n134 & n217 ) | ( ~n205 & n217 ) ;
  assign n235 = ( n208 & n229 ) | ( n208 & n234 ) | ( n229 & n234 ) ;
  assign n236 = ( ~n134 & n231 ) | ( ~n134 & n234 ) | ( n231 & n234 ) ;
  assign n237 = n236 ^ n206 ^ 1'b0 ;
  assign n238 = ( n227 & ~n228 ) | ( n227 & n232 ) | ( ~n228 & n232 ) ;
  assign n239 = n229 | n235 ;
  assign n240 = n206 & ~n236 ;
  assign n241 = ( n236 & ~n239 ) | ( n236 & n240 ) | ( ~n239 & n240 ) ;
  assign n242 = x18 | x19 ;
  assign n243 = x20 & n217 ;
  assign n244 = x20 | n242 ;
  assign n245 = ( x20 & ~n148 ) | ( x20 & n242 ) | ( ~n148 & n242 ) ;
  assign n246 = n238 ^ x23 ^ 1'b0 ;
  assign n247 = ( n183 & ~n243 ) | ( n183 & n245 ) | ( ~n243 & n245 ) ;
  assign n248 = ~n183 & n247 ;
  assign n249 = n243 ^ n217 ^ x21 ;
  assign n250 = ( n179 & n243 ) | ( n179 & ~n244 ) | ( n243 & ~n244 ) ;
  assign n251 = n248 | n249 ;
  assign n252 = ~n250 & n251 ;
  assign n253 = ( ~n144 & n246 ) | ( ~n144 & n252 ) | ( n246 & n252 ) ;
  assign n254 = ( ~n134 & n222 ) | ( ~n134 & n253 ) | ( n222 & n253 ) ;
  assign n255 = n237 | n254 ;
  assign n256 = ( ~x30 & n218 ) | ( ~x30 & n255 ) | ( n218 & n255 ) ;
  assign n257 = ~n136 & n256 ;
  assign n258 = x16 | x17 ;
  assign n259 = n237 & n254 ;
  assign n260 = n257 | n259 ;
  assign n261 = n229 | n260 ;
  assign n262 = n261 ^ n253 ^ n134 ;
  assign n263 = n261 & n262 ;
  assign n264 = n261 ^ n252 ^ n144 ;
  assign n265 = n263 ^ n220 ^ n192 ;
  assign n266 = n248 & n261 ;
  assign n267 = ( n241 & n257 ) | ( n241 & ~n259 ) | ( n257 & ~n259 ) ;
  assign n268 = x18 & n261 ;
  assign n269 = ( ~x18 & n217 ) | ( ~x18 & n261 ) | ( n217 & n261 ) ;
  assign n270 = ( x18 & n217 ) | ( x18 & ~n258 ) | ( n217 & ~n258 ) ;
  assign n271 = n269 & n270 ;
  assign n272 = ~n242 & n261 ;
  assign n273 = ( n250 & n261 ) | ( n250 & ~n266 ) | ( n261 & ~n266 ) ;
  assign n274 = ( x18 & ~n216 ) | ( x18 & n258 ) | ( ~n216 & n258 ) ;
  assign n275 = ( ~n217 & n268 ) | ( ~n217 & n274 ) | ( n268 & n274 ) ;
  assign n276 = n260 & ~n272 ;
  assign n277 = ( n233 & n272 ) | ( n233 & ~n276 ) | ( n272 & ~n276 ) ;
  assign n278 = n277 ^ x20 ^ 1'b0 ;
  assign n279 = ~n268 & n275 ;
  assign n280 = n261 & n264 ;
  assign n281 = n257 & n267 ;
  assign n282 = ( ~n255 & n259 ) | ( ~n255 & n261 ) | ( n259 & n261 ) ;
  assign n283 = ( n136 & n237 ) | ( n136 & n254 ) | ( n237 & n254 ) ;
  assign n284 = ( n254 & n259 ) | ( n254 & ~n261 ) | ( n259 & ~n261 ) ;
  assign n285 = n283 & ~n284 ;
  assign n286 = ( n267 & ~n281 ) | ( n267 & n285 ) | ( ~n281 & n285 ) ;
  assign n287 = ( n257 & n261 ) | ( n257 & ~n286 ) | ( n261 & ~n286 ) ;
  assign n288 = n280 ^ n238 ^ x23 ;
  assign n289 = n268 ^ n261 ^ x19 ;
  assign n290 = n279 | n289 ;
  assign n291 = ~n271 & n290 ;
  assign n292 = n273 ^ n250 ^ n249 ;
  assign n293 = ( ~n179 & n278 ) | ( ~n179 & n291 ) | ( n278 & n291 ) ;
  assign n294 = ( ~n144 & n292 ) | ( ~n144 & n293 ) | ( n292 & n293 ) ;
  assign n295 = n293 ^ n144 ^ 1'b0 ;
  assign n296 = ( ~n134 & n288 ) | ( ~n134 & n294 ) | ( n288 & n294 ) ;
  assign n297 = n265 | n296 ;
  assign n298 = n265 & n296 ;
  assign n299 = ( ~x30 & n282 ) | ( ~x30 & n297 ) | ( n282 & n297 ) ;
  assign n300 = ~n136 & n299 ;
  assign n301 = n298 | n300 ;
  assign n302 = n286 | n301 ;
  assign n303 = n295 & n302 ;
  assign n304 = ~n258 & n302 ;
  assign n305 = n303 ^ n302 ^ n292 ;
  assign n306 = n301 & ~n304 ;
  assign n307 = n302 ^ n294 ^ n134 ;
  assign n308 = n302 & n307 ;
  assign n309 = n308 ^ n280 ^ n246 ;
  assign n310 = ( n287 & n304 ) | ( n287 & ~n306 ) | ( n304 & ~n306 ) ;
  assign n311 = n279 & n302 ;
  assign n312 = ( n271 & n302 ) | ( n271 & ~n311 ) | ( n302 & ~n311 ) ;
  assign n313 = n312 ^ n289 ^ n271 ;
  assign n314 = ( n265 & n297 ) | ( n265 & n302 ) | ( n297 & n302 ) ;
  assign n315 = x16 & n302 ;
  assign n316 = n315 ^ n302 ^ x17 ;
  assign n317 = x14 | x15 ;
  assign n318 = n310 ^ x18 ^ 1'b0 ;
  assign n319 = x16 | n317 ;
  assign n320 = ( n261 & n315 ) | ( n261 & ~n319 ) | ( n315 & ~n319 ) ;
  assign n321 = ( x16 & ~n260 ) | ( x16 & n317 ) | ( ~n260 & n317 ) ;
  assign n322 = n302 ^ n291 ^ n179 ;
  assign n323 = ~n302 & n314 ;
  assign n324 = ( ~n297 & n298 ) | ( ~n297 & n302 ) | ( n298 & n302 ) ;
  assign n325 = n302 & n322 ;
  assign n326 = ( ~n261 & n315 ) | ( ~n261 & n321 ) | ( n315 & n321 ) ;
  assign n327 = ( ~n136 & n298 ) | ( ~n136 & n324 ) | ( n298 & n324 ) ;
  assign n328 = n325 ^ n277 ^ x20 ;
  assign n329 = ( ~n136 & n265 ) | ( ~n136 & n296 ) | ( n265 & n296 ) ;
  assign n330 = ~n315 & n326 ;
  assign n331 = n316 | n330 ;
  assign n332 = ~n320 & n331 ;
  assign n333 = ( ~n217 & n318 ) | ( ~n217 & n332 ) | ( n318 & n332 ) ;
  assign n334 = ( ~n179 & n313 ) | ( ~n179 & n333 ) | ( n313 & n333 ) ;
  assign n335 = ( ~n144 & n328 ) | ( ~n144 & n334 ) | ( n328 & n334 ) ;
  assign n336 = ( ~n134 & n305 ) | ( ~n134 & n335 ) | ( n305 & n335 ) ;
  assign n337 = n309 | n336 ;
  assign n338 = n333 ^ n179 ^ 1'b0 ;
  assign n339 = ( ~x30 & n327 ) | ( ~x30 & n337 ) | ( n327 & n337 ) ;
  assign n340 = ( n314 & n323 ) | ( n314 & ~n329 ) | ( n323 & ~n329 ) ;
  assign n341 = n309 & n336 ;
  assign n342 = ( n300 & n302 ) | ( n300 & ~n340 ) | ( n302 & ~n340 ) ;
  assign n343 = ~n136 & n339 ;
  assign n344 = n341 | n343 ;
  assign n345 = n340 | n344 ;
  assign n346 = n345 ^ n332 ^ n217 ;
  assign n347 = n345 & n346 ;
  assign n348 = n347 ^ n310 ^ x18 ;
  assign n349 = n345 ^ n334 ^ n144 ;
  assign n350 = n345 & n349 ;
  assign n351 = n350 ^ n325 ^ n278 ;
  assign n352 = ( n134 & ~n335 ) | ( n134 & n345 ) | ( ~n335 & n345 ) ;
  assign n353 = n335 ^ n134 ^ 1'b0 ;
  assign n354 = ( n309 & n337 ) | ( n309 & n345 ) | ( n337 & n345 ) ;
  assign n355 = ( ~n337 & n341 ) | ( ~n337 & n345 ) | ( n341 & n345 ) ;
  assign n356 = ( ~n136 & n309 ) | ( ~n136 & n336 ) | ( n309 & n336 ) ;
  assign n357 = ~n345 & n354 ;
  assign n358 = ( n354 & ~n356 ) | ( n354 & n357 ) | ( ~n356 & n357 ) ;
  assign n359 = n336 | n358 ;
  assign n360 = ( n343 & n345 ) | ( n343 & ~n358 ) | ( n345 & ~n358 ) ;
  assign n361 = ~n317 & n345 ;
  assign n362 = n344 & ~n361 ;
  assign n363 = n338 & n345 ;
  assign n364 = n363 ^ n345 ^ n313 ;
  assign n365 = ( n342 & n361 ) | ( n342 & ~n362 ) | ( n361 & ~n362 ) ;
  assign n366 = n345 & ~n353 ;
  assign n367 = n366 ^ n305 ^ 1'b0 ;
  assign n368 = n330 & n345 ;
  assign n369 = ( n320 & n345 ) | ( n320 & ~n368 ) | ( n345 & ~n368 ) ;
  assign n370 = n369 ^ n320 ^ n316 ;
  assign n371 = ( n352 & n358 ) | ( n352 & n359 ) | ( n358 & n359 ) ;
  assign n372 = ( n305 & n366 ) | ( n305 & ~n371 ) | ( n366 & ~n371 ) ;
  assign n373 = ~n371 & n372 ;
  assign n374 = x12 | x13 ;
  assign n375 = ( ~x14 & n302 ) | ( ~x14 & n345 ) | ( n302 & n345 ) ;
  assign n376 = x14 & n345 ;
  assign n377 = ( x14 & ~n301 ) | ( x14 & n374 ) | ( ~n301 & n374 ) ;
  assign n378 = ( ~n302 & n376 ) | ( ~n302 & n377 ) | ( n376 & n377 ) ;
  assign n379 = n376 ^ n345 ^ x15 ;
  assign n380 = ~n376 & n378 ;
  assign n381 = n365 ^ x16 ^ 1'b0 ;
  assign n382 = n379 | n380 ;
  assign n383 = ( x14 & n302 ) | ( x14 & ~n374 ) | ( n302 & ~n374 ) ;
  assign n384 = n375 & n383 ;
  assign n385 = n382 & ~n384 ;
  assign n386 = ( ~n261 & n381 ) | ( ~n261 & n385 ) | ( n381 & n385 ) ;
  assign n387 = ( ~n217 & n370 ) | ( ~n217 & n386 ) | ( n370 & n386 ) ;
  assign n388 = ( ~n179 & n348 ) | ( ~n179 & n387 ) | ( n348 & n387 ) ;
  assign n389 = ( ~n144 & n364 ) | ( ~n144 & n388 ) | ( n364 & n388 ) ;
  assign n390 = ( ~n134 & n351 ) | ( ~n134 & n389 ) | ( n351 & n389 ) ;
  assign n391 = ( ~n136 & n367 ) | ( ~n136 & n390 ) | ( n367 & n390 ) ;
  assign n392 = ~n136 & n391 ;
  assign n393 = ( ~n136 & n355 ) | ( ~n136 & n392 ) | ( n355 & n392 ) ;
  assign n394 = n367 & n390 ;
  assign n395 = ( n373 & n393 ) | ( n373 & ~n394 ) | ( n393 & ~n394 ) ;
  assign n396 = ~n393 & n395 ;
  assign n397 = n386 ^ n217 ^ 1'b0 ;
  assign n398 = n393 | n394 ;
  assign n399 = n358 | n398 ;
  assign n400 = ~n374 & n399 ;
  assign n401 = n397 & n399 ;
  assign n402 = n401 ^ n399 ^ n370 ;
  assign n403 = n398 & ~n400 ;
  assign n404 = ( n360 & n400 ) | ( n360 & ~n403 ) | ( n400 & ~n403 ) ;
  assign n405 = n399 ^ n387 ^ n179 ;
  assign n406 = n399 & n405 ;
  assign n407 = ( n390 & n391 ) | ( n390 & n399 ) | ( n391 & n399 ) ;
  assign n408 = n399 ^ n385 ^ n261 ;
  assign n409 = n399 ^ n389 ^ n134 ;
  assign n410 = n399 & n408 ;
  assign n411 = n388 ^ n144 ^ 1'b0 ;
  assign n412 = n399 & n411 ;
  assign n413 = n380 & n399 ;
  assign n414 = ( n134 & ~n389 ) | ( n134 & n399 ) | ( ~n389 & n399 ) ;
  assign n415 = n412 ^ n399 ^ n364 ;
  assign n416 = n410 ^ n365 ^ x16 ;
  assign n417 = ( n384 & n399 ) | ( n384 & ~n413 ) | ( n399 & ~n413 ) ;
  assign n418 = n367 & ~n407 ;
  assign n419 = ( ~n367 & n394 ) | ( ~n367 & n399 ) | ( n394 & n399 ) ;
  assign n420 = n418 ^ n407 ^ n391 ;
  assign n421 = n406 ^ n347 ^ n318 ;
  assign n422 = n396 | n420 ;
  assign n423 = ( ~n390 & n394 ) | ( ~n390 & n419 ) | ( n394 & n419 ) ;
  assign n424 = n399 & n409 ;
  assign n425 = n424 ^ n351 ^ 1'b0 ;
  assign n426 = n390 | n422 ;
  assign n427 = ( n414 & n422 ) | ( n414 & n426 ) | ( n422 & n426 ) ;
  assign n428 = ( n351 & n424 ) | ( n351 & ~n427 ) | ( n424 & ~n427 ) ;
  assign n429 = n417 ^ n384 ^ n379 ;
  assign n430 = ~n427 & n428 ;
  assign n431 = x9 | x10 ;
  assign n432 = x12 & n399 ;
  assign n433 = ( x12 & n345 ) | ( x12 & ~n431 ) | ( n345 & ~n431 ) ;
  assign n434 = ( ~x12 & n345 ) | ( ~x12 & n399 ) | ( n345 & n399 ) ;
  assign n435 = n433 & n434 ;
  assign n436 = ( x12 & ~n344 ) | ( x12 & n431 ) | ( ~n344 & n431 ) ;
  assign n437 = n432 ^ n399 ^ x13 ;
  assign n438 = ( ~n345 & n432 ) | ( ~n345 & n436 ) | ( n432 & n436 ) ;
  assign n439 = ~n432 & n438 ;
  assign n440 = n437 | n439 ;
  assign n441 = ~n435 & n440 ;
  assign n442 = n404 ^ x14 ^ 1'b0 ;
  assign n443 = ( ~n302 & n441 ) | ( ~n302 & n442 ) | ( n441 & n442 ) ;
  assign n444 = n443 ^ n261 ^ 1'b0 ;
  assign n445 = ( ~n261 & n429 ) | ( ~n261 & n443 ) | ( n429 & n443 ) ;
  assign n446 = ( ~n217 & n416 ) | ( ~n217 & n445 ) | ( n416 & n445 ) ;
  assign n447 = n435 | n439 ;
  assign n448 = ( ~n179 & n402 ) | ( ~n179 & n446 ) | ( n402 & n446 ) ;
  assign n449 = ( ~n144 & n421 ) | ( ~n144 & n448 ) | ( n421 & n448 ) ;
  assign n450 = ( ~n134 & n415 ) | ( ~n134 & n449 ) | ( n415 & n449 ) ;
  assign n451 = n449 ^ n134 ^ 1'b0 ;
  assign n452 = n446 ^ n179 ^ 1'b0 ;
  assign n453 = n425 | n450 ;
  assign n454 = ( ~x30 & n423 ) | ( ~x30 & n453 ) | ( n423 & n453 ) ;
  assign n455 = ~n136 & n454 ;
  assign n456 = n425 & n450 ;
  assign n457 = n455 | n456 ;
  assign n458 = n422 | n457 ;
  assign n459 = n458 ^ n448 ^ n144 ;
  assign n460 = n458 & n459 ;
  assign n461 = ~n431 & n458 ;
  assign n462 = ( ~n453 & n456 ) | ( ~n453 & n458 ) | ( n456 & n458 ) ;
  assign n463 = n460 ^ n406 ^ n348 ;
  assign n464 = n458 ^ n445 ^ n217 ;
  assign n465 = n458 ^ n441 ^ n302 ;
  assign n466 = n444 & n458 ;
  assign n467 = n458 & n465 ;
  assign n468 = n467 ^ n404 ^ x14 ;
  assign n469 = n447 & n458 ;
  assign n470 = n469 ^ n458 ^ n437 ;
  assign n471 = n458 & n464 ;
  assign n472 = ( n430 & n455 ) | ( n430 & ~n456 ) | ( n455 & ~n456 ) ;
  assign n473 = n452 & n458 ;
  assign n474 = n471 ^ n410 ^ n381 ;
  assign n475 = n466 ^ n458 ^ n429 ;
  assign n476 = ~n455 & n472 ;
  assign n477 = ( n136 & n450 ) | ( n136 & n456 ) | ( n450 & n456 ) ;
  assign n478 = ( n456 & ~n458 ) | ( n456 & n477 ) | ( ~n458 & n477 ) ;
  assign n479 = ( n136 & n425 ) | ( n136 & n450 ) | ( n425 & n450 ) ;
  assign n480 = n451 & n458 ;
  assign n481 = n399 & ~n420 ;
  assign n482 = n479 ^ n478 ^ 1'b0 ;
  assign n483 = ( n396 & n457 ) | ( n396 & ~n461 ) | ( n457 & ~n461 ) ;
  assign n484 = n480 ^ n458 ^ n415 ;
  assign n485 = n473 ^ n458 ^ n402 ;
  assign n486 = n461 | n481 ;
  assign n487 = n476 | n482 ;
  assign n488 = ( n455 & n462 ) | ( n455 & ~n487 ) | ( n462 & ~n487 ) ;
  assign n489 = ( n461 & ~n483 ) | ( n461 & n486 ) | ( ~n483 & n486 ) ;
  assign n490 = n489 ^ x12 ^ 1'b0 ;
  assign n491 = x7 | x8 ;
  assign n492 = ( x9 & n399 ) | ( x9 & ~n491 ) | ( n399 & ~n491 ) ;
  assign n493 = ( ~x9 & n399 ) | ( ~x9 & n458 ) | ( n399 & n458 ) ;
  assign n494 = n492 & n493 ;
  assign n495 = x9 & n458 ;
  assign n496 = n495 ^ n458 ^ x10 ;
  assign n497 = ( x9 & ~n398 ) | ( x9 & n491 ) | ( ~n398 & n491 ) ;
  assign n498 = ( ~n399 & n495 ) | ( ~n399 & n497 ) | ( n495 & n497 ) ;
  assign n499 = ~n495 & n498 ;
  assign n500 = n496 | n499 ;
  assign n501 = ~n494 & n500 ;
  assign n502 = ( ~n345 & n490 ) | ( ~n345 & n501 ) | ( n490 & n501 ) ;
  assign n503 = ( ~n302 & n470 ) | ( ~n302 & n502 ) | ( n470 & n502 ) ;
  assign n504 = ( ~n261 & n468 ) | ( ~n261 & n503 ) | ( n468 & n503 ) ;
  assign n505 = ( ~n217 & n475 ) | ( ~n217 & n504 ) | ( n475 & n504 ) ;
  assign n506 = ( ~n179 & n474 ) | ( ~n179 & n505 ) | ( n474 & n505 ) ;
  assign n507 = ( ~n144 & n485 ) | ( ~n144 & n506 ) | ( n485 & n506 ) ;
  assign n508 = ( ~n134 & n463 ) | ( ~n134 & n507 ) | ( n463 & n507 ) ;
  assign n509 = n484 & n508 ;
  assign n510 = n484 | n508 ;
  assign n511 = ( ~x30 & n462 ) | ( ~x30 & n510 ) | ( n462 & n510 ) ;
  assign n512 = n136 & ~n509 ;
  assign n513 = ( n509 & n511 ) | ( n509 & ~n512 ) | ( n511 & ~n512 ) ;
  assign n514 = n487 | n513 ;
  assign n515 = ( n136 & n484 ) | ( n136 & n508 ) | ( n484 & n508 ) ;
  assign n516 = ( n136 & n508 ) | ( n136 & n509 ) | ( n508 & n509 ) ;
  assign n517 = ( n509 & ~n514 ) | ( n509 & n516 ) | ( ~n514 & n516 ) ;
  assign n518 = n517 ^ n515 ^ 1'b0 ;
  assign n519 = ( n484 & ~n514 ) | ( n484 & n518 ) | ( ~n514 & n518 ) ;
  assign n520 = ~n491 & n514 ;
  assign n521 = n513 & ~n520 ;
  assign n522 = ( n488 & n520 ) | ( n488 & ~n521 ) | ( n520 & ~n521 ) ;
  assign n523 = n499 & n514 ;
  assign n524 = ( n494 & n514 ) | ( n494 & ~n523 ) | ( n514 & ~n523 ) ;
  assign n525 = n524 ^ n496 ^ n494 ;
  assign n526 = n514 ^ n501 ^ n345 ;
  assign n527 = n514 & n526 ;
  assign n528 = n527 ^ n489 ^ x12 ;
  assign n529 = n502 ^ n302 ^ 1'b0 ;
  assign n530 = n514 & n529 ;
  assign n531 = n530 ^ n514 ^ n470 ;
  assign n532 = n514 ^ n503 ^ n261 ;
  assign n533 = n504 ^ n217 ^ 1'b0 ;
  assign n534 = n514 & n533 ;
  assign n535 = n534 ^ n514 ^ n475 ;
  assign n536 = n514 ^ n505 ^ n179 ;
  assign n537 = n514 & n536 ;
  assign n538 = n537 ^ n471 ^ n416 ;
  assign n539 = n506 ^ n144 ^ 1'b0 ;
  assign n540 = n514 & n539 ;
  assign n541 = n540 ^ n514 ^ n485 ;
  assign n542 = n514 ^ n507 ^ n134 ;
  assign n543 = n514 & n542 ;
  assign n544 = n543 ^ n460 ^ n421 ;
  assign n545 = n514 & n532 ;
  assign n546 = n545 ^ n467 ^ n442 ;
  assign n547 = ( n509 & ~n510 ) | ( n509 & n514 ) | ( ~n510 & n514 ) ;
  assign n548 = ( ~n136 & n509 ) | ( ~n136 & n547 ) | ( n509 & n547 ) ;
  assign n549 = n522 ^ x9 ^ 1'b0 ;
  assign n550 = x5 | x6 ;
  assign n551 = x7 | n550 ;
  assign n552 = x7 & n514 ;
  assign n553 = ( n458 & ~n551 ) | ( n458 & n552 ) | ( ~n551 & n552 ) ;
  assign n554 = n552 ^ n514 ^ x8 ;
  assign n555 = ( x7 & ~n457 ) | ( x7 & n550 ) | ( ~n457 & n550 ) ;
  assign n556 = ( ~n458 & n552 ) | ( ~n458 & n555 ) | ( n552 & n555 ) ;
  assign n557 = ~n552 & n556 ;
  assign n558 = n554 | n557 ;
  assign n559 = ~n553 & n558 ;
  assign n560 = ( ~n399 & n549 ) | ( ~n399 & n559 ) | ( n549 & n559 ) ;
  assign n561 = ( ~n345 & n525 ) | ( ~n345 & n560 ) | ( n525 & n560 ) ;
  assign n562 = ( ~n302 & n528 ) | ( ~n302 & n561 ) | ( n528 & n561 ) ;
  assign n563 = ( ~n261 & n531 ) | ( ~n261 & n562 ) | ( n531 & n562 ) ;
  assign n564 = ( ~n217 & n546 ) | ( ~n217 & n563 ) | ( n546 & n563 ) ;
  assign n565 = ( ~n179 & n535 ) | ( ~n179 & n564 ) | ( n535 & n564 ) ;
  assign n566 = ( ~n144 & n538 ) | ( ~n144 & n565 ) | ( n538 & n565 ) ;
  assign n567 = ( ~n134 & n541 ) | ( ~n134 & n566 ) | ( n541 & n566 ) ;
  assign n568 = ( ~n136 & n544 ) | ( ~n136 & n567 ) | ( n544 & n567 ) ;
  assign n569 = n136 & ~n568 ;
  assign n570 = ( n548 & n568 ) | ( n548 & ~n569 ) | ( n568 & ~n569 ) ;
  assign n571 = ( ~n518 & n519 ) | ( ~n518 & n570 ) | ( n519 & n570 ) ;
  assign n572 = n518 | n571 ;
  assign n573 = n566 ^ n134 ^ 1'b0 ;
  assign n574 = ~n550 & n572 ;
  assign n575 = ( n514 & ~n518 ) | ( n514 & n574 ) | ( ~n518 & n574 ) ;
  assign n576 = n570 & ~n574 ;
  assign n577 = ( n574 & n575 ) | ( n574 & ~n576 ) | ( n575 & ~n576 ) ;
  assign n578 = n557 & n572 ;
  assign n579 = ( n553 & n572 ) | ( n553 & ~n578 ) | ( n572 & ~n578 ) ;
  assign n580 = n579 ^ n554 ^ n553 ;
  assign n581 = n572 ^ n559 ^ n399 ;
  assign n582 = n560 ^ n345 ^ 1'b0 ;
  assign n583 = n572 & n582 ;
  assign n584 = n583 ^ n572 ^ n525 ;
  assign n585 = n572 ^ n561 ^ n302 ;
  assign n586 = n572 & n585 ;
  assign n587 = n586 ^ n527 ^ n490 ;
  assign n588 = n562 ^ n261 ^ 1'b0 ;
  assign n589 = n572 & n588 ;
  assign n590 = n589 ^ n572 ^ n531 ;
  assign n591 = n572 & n573 ;
  assign n592 = n591 ^ n572 ^ n541 ;
  assign n593 = n572 ^ n563 ^ n217 ;
  assign n594 = n572 & n593 ;
  assign n595 = n594 ^ n545 ^ n468 ;
  assign n596 = n564 ^ n179 ^ 1'b0 ;
  assign n597 = n572 & n596 ;
  assign n598 = n597 ^ n572 ^ n535 ;
  assign n599 = n572 ^ n565 ^ n144 ;
  assign n600 = n572 & n599 ;
  assign n601 = n600 ^ n537 ^ n474 ;
  assign n602 = x5 & n572 ;
  assign n603 = n577 ^ x7 ^ 1'b0 ;
  assign n604 = n602 ^ n572 ^ x6 ;
  assign n605 = n572 & n581 ;
  assign n606 = ( ~x5 & n514 ) | ( ~x5 & n572 ) | ( n514 & n572 ) ;
  assign n607 = x3 | x4 ;
  assign n608 = ( x5 & n514 ) | ( x5 & ~n607 ) | ( n514 & ~n607 ) ;
  assign n609 = n605 ^ n522 ^ x9 ;
  assign n610 = n606 & n608 ;
  assign n611 = ( x5 & ~n513 ) | ( x5 & n607 ) | ( ~n513 & n607 ) ;
  assign n612 = ( ~n514 & n602 ) | ( ~n514 & n611 ) | ( n602 & n611 ) ;
  assign n613 = ~n602 & n612 ;
  assign n614 = n604 | n613 ;
  assign n615 = ~n610 & n614 ;
  assign n616 = ( ~n458 & n603 ) | ( ~n458 & n615 ) | ( n603 & n615 ) ;
  assign n617 = ( ~n399 & n580 ) | ( ~n399 & n616 ) | ( n580 & n616 ) ;
  assign n618 = ( n136 & n544 ) | ( n136 & n567 ) | ( n544 & n567 ) ;
  assign n619 = ( ~n345 & n609 ) | ( ~n345 & n617 ) | ( n609 & n617 ) ;
  assign n620 = n572 ^ n567 ^ n544 ;
  assign n621 = ( ~n302 & n584 ) | ( ~n302 & n619 ) | ( n584 & n619 ) ;
  assign n622 = n544 & ~n572 ;
  assign n623 = ~n567 & n618 ;
  assign n624 = ( n544 & n567 ) | ( n544 & ~n572 ) | ( n567 & ~n572 ) ;
  assign n625 = n610 | n613 ;
  assign n626 = ( n618 & n623 ) | ( n618 & ~n624 ) | ( n623 & ~n624 ) ;
  assign n627 = n622 | n626 ;
  assign n628 = n616 ^ n399 ^ 1'b0 ;
  assign n629 = ( ~n261 & n587 ) | ( ~n261 & n621 ) | ( n587 & n621 ) ;
  assign n630 = ( ~n217 & n590 ) | ( ~n217 & n629 ) | ( n590 & n629 ) ;
  assign n631 = ( ~n179 & n595 ) | ( ~n179 & n630 ) | ( n595 & n630 ) ;
  assign n632 = ( ~n144 & n598 ) | ( ~n144 & n631 ) | ( n598 & n631 ) ;
  assign n633 = n572 & n620 ;
  assign n634 = ( ~n134 & n601 ) | ( ~n134 & n632 ) | ( n601 & n632 ) ;
  assign n635 = n592 | n634 ;
  assign n636 = ( ~x30 & n633 ) | ( ~x30 & n635 ) | ( n633 & n635 ) ;
  assign n637 = ~n136 & n636 ;
  assign n638 = n592 & n634 ;
  assign n639 = n637 | n638 ;
  assign n640 = n627 | n639 ;
  assign n641 = n625 & n640 ;
  assign n642 = n641 ^ n640 ^ n604 ;
  assign n643 = n640 ^ n617 ^ n345 ;
  assign n644 = n640 & n643 ;
  assign n645 = n640 ^ n621 ^ n261 ;
  assign n646 = n629 ^ n217 ^ 1'b0 ;
  assign n647 = n619 ^ n302 ^ 1'b0 ;
  assign n648 = n640 & n646 ;
  assign n649 = n640 & n647 ;
  assign n650 = n649 ^ n640 ^ n584 ;
  assign n651 = n640 & n645 ;
  assign n652 = n651 ^ n586 ^ n528 ;
  assign n653 = n644 ^ n605 ^ n549 ;
  assign n654 = n628 & n640 ;
  assign n655 = n654 ^ n640 ^ n580 ;
  assign n656 = n648 ^ n640 ^ n590 ;
  assign n657 = ~n607 & n640 ;
  assign n658 = x1 | x2 ;
  assign n659 = n626 & ~n657 ;
  assign n660 = ( x3 & ~n570 ) | ( x3 & n658 ) | ( ~n570 & n658 ) ;
  assign n661 = n640 ^ n615 ^ n458 ;
  assign n662 = ( n572 & ~n639 ) | ( n572 & n657 ) | ( ~n639 & n657 ) ;
  assign n663 = ( n136 & n592 ) | ( n136 & n634 ) | ( n592 & n634 ) ;
  assign n664 = ( n634 & n638 ) | ( n634 & ~n640 ) | ( n638 & ~n640 ) ;
  assign n665 = n640 ^ n632 ^ n134 ;
  assign n666 = n640 & n665 ;
  assign n667 = n666 ^ n601 ^ 1'b0 ;
  assign n668 = n663 & ~n664 ;
  assign n669 = ( n134 & ~n632 ) | ( n134 & n640 ) | ( ~n632 & n640 ) ;
  assign n670 = n592 & ~n640 ;
  assign n671 = n668 | n670 ;
  assign n672 = n634 | n671 ;
  assign n673 = ( n669 & n671 ) | ( n669 & n672 ) | ( n671 & n672 ) ;
  assign n674 = ( n601 & n666 ) | ( n601 & ~n673 ) | ( n666 & ~n673 ) ;
  assign n675 = ~n673 & n674 ;
  assign n676 = x3 & n640 ;
  assign n677 = n676 ^ n640 ^ x4 ;
  assign n678 = ( ~n572 & n660 ) | ( ~n572 & n676 ) | ( n660 & n676 ) ;
  assign n679 = ~n676 & n678 ;
  assign n680 = ( n657 & ~n659 ) | ( n657 & n662 ) | ( ~n659 & n662 ) ;
  assign n681 = n677 | n679 ;
  assign n682 = n680 ^ x5 ^ 1'b0 ;
  assign n683 = n640 & n661 ;
  assign n684 = n683 ^ n577 ^ x7 ;
  assign n685 = x3 | n658 ;
  assign n686 = ( n572 & n676 ) | ( n572 & ~n685 ) | ( n676 & ~n685 ) ;
  assign n687 = ( ~n635 & n638 ) | ( ~n635 & n640 ) | ( n638 & n640 ) ;
  assign n688 = n681 & ~n686 ;
  assign n689 = n640 ^ n630 ^ n179 ;
  assign n690 = ( ~n514 & n682 ) | ( ~n514 & n688 ) | ( n682 & n688 ) ;
  assign n691 = ( x1 & x125 ) | ( x1 & ~n639 ) | ( x125 & ~n639 ) ;
  assign n692 = ( ~n458 & n642 ) | ( ~n458 & n690 ) | ( n642 & n690 ) ;
  assign n693 = n640 & n689 ;
  assign n694 = n631 ^ n144 ^ 1'b0 ;
  assign n695 = n640 & n694 ;
  assign n696 = n693 ^ n594 ^ n546 ;
  assign n697 = n695 ^ n640 ^ n598 ;
  assign n698 = ( ~n399 & n684 ) | ( ~n399 & n692 ) | ( n684 & n692 ) ;
  assign n699 = ( ~n345 & n655 ) | ( ~n345 & n698 ) | ( n655 & n698 ) ;
  assign n700 = n698 ^ n345 ^ 1'b0 ;
  assign n701 = n690 ^ n458 ^ 1'b0 ;
  assign n702 = ( x126 & ~n639 ) | ( x126 & n691 ) | ( ~n639 & n691 ) ;
  assign n703 = ( ~n302 & n653 ) | ( ~n302 & n699 ) | ( n653 & n699 ) ;
  assign n704 = ( ~n261 & n650 ) | ( ~n261 & n703 ) | ( n650 & n703 ) ;
  assign n705 = ( ~n217 & n652 ) | ( ~n217 & n704 ) | ( n652 & n704 ) ;
  assign n706 = ( ~n179 & n656 ) | ( ~n179 & n705 ) | ( n656 & n705 ) ;
  assign n707 = ( ~n144 & n696 ) | ( ~n144 & n706 ) | ( n696 & n706 ) ;
  assign n708 = ( ~n134 & n697 ) | ( ~n134 & n707 ) | ( n697 & n707 ) ;
  assign n709 = n667 | n708 ;
  assign n710 = n707 ^ n134 ^ 1'b0 ;
  assign n711 = ( ~x30 & n687 ) | ( ~x30 & n709 ) | ( n687 & n709 ) ;
  assign n712 = ~n136 & n711 ;
  assign n713 = n705 ^ n179 ^ 1'b0 ;
  assign n714 = n667 & n708 ;
  assign n715 = n712 | n714 ;
  assign n716 = n671 | n715 ;
  assign n717 = n716 ^ n699 ^ n302 ;
  assign n718 = n716 & n717 ;
  assign n719 = n718 ^ n644 ^ n609 ;
  assign n720 = ( x1 & n639 ) | ( x1 & n716 ) | ( n639 & n716 ) ;
  assign n721 = n703 ^ n261 ^ 1'b0 ;
  assign n722 = n716 ^ n688 ^ n514 ;
  assign n723 = ( ~n709 & n714 ) | ( ~n709 & n716 ) | ( n714 & n716 ) ;
  assign n724 = ( n136 & n708 ) | ( n136 & n714 ) | ( n708 & n714 ) ;
  assign n725 = n716 ^ n704 ^ n217 ;
  assign n726 = n716 & n725 ;
  assign n727 = n716 & n722 ;
  assign n728 = n726 ^ n651 ^ n587 ;
  assign n729 = ~n658 & n716 ;
  assign n730 = ( n136 & n667 ) | ( n136 & n708 ) | ( n667 & n708 ) ;
  assign n731 = n701 & n716 ;
  assign n732 = n713 & n716 ;
  assign n733 = n727 ^ n680 ^ x5 ;
  assign n734 = n732 ^ n716 ^ n656 ;
  assign n735 = ~n136 & n723 ;
  assign n736 = n679 & n716 ;
  assign n737 = n731 ^ n716 ^ n642 ;
  assign n738 = ( n686 & n716 ) | ( n686 & ~n736 ) | ( n716 & ~n736 ) ;
  assign n739 = n738 ^ n686 ^ n677 ;
  assign n740 = n710 & n716 ;
  assign n741 = n716 ^ n706 ^ n144 ;
  assign n742 = n716 & n721 ;
  assign n743 = n700 & n716 ;
  assign n744 = n668 & ~n729 ;
  assign n745 = n740 ^ n716 ^ n697 ;
  assign n746 = ( n640 & ~n715 ) | ( n640 & n729 ) | ( ~n715 & n729 ) ;
  assign n747 = n716 & n741 ;
  assign n748 = ( n729 & ~n744 ) | ( n729 & n746 ) | ( ~n744 & n746 ) ;
  assign n749 = n742 ^ n716 ^ n650 ;
  assign n750 = ( n675 & n712 ) | ( n675 & ~n714 ) | ( n712 & ~n714 ) ;
  assign n751 = ~n712 & n750 ;
  assign n752 = n747 ^ n693 ^ n595 ;
  assign n753 = n716 ^ n692 ^ n399 ;
  assign n754 = ( n714 & ~n716 ) | ( n714 & n724 ) | ( ~n716 & n724 ) ;
  assign n755 = n716 & n753 ;
  assign n756 = ( ~n627 & n702 ) | ( ~n627 & n720 ) | ( n702 & n720 ) ;
  assign n757 = n743 ^ n716 ^ n655 ;
  assign n758 = n754 ^ n730 ^ 1'b0 ;
  assign n759 = n751 | n758 ;
  assign n760 = ( n712 & n723 ) | ( n712 & ~n759 ) | ( n723 & ~n759 ) ;
  assign n761 = n755 ^ n683 ^ n603 ;
  assign n762 = ~n720 & n756 ;
  assign n763 = n748 ^ x3 ^ 1'b0 ;
  assign n764 = x125 | x126 ;
  assign n765 = ( x1 & n640 ) | ( x1 & ~n764 ) | ( n640 & ~n764 ) ;
  assign n766 = ( ~x1 & n640 ) | ( ~x1 & n716 ) | ( n640 & n716 ) ;
  assign n767 = n765 & n766 ;
  assign n768 = ~x1 & n716 ;
  assign n769 = n768 ^ x2 ^ 1'b0 ;
  assign n770 = n762 | n769 ;
  assign n771 = ~n767 & n770 ;
  assign n772 = ( ~n572 & n763 ) | ( ~n572 & n771 ) | ( n763 & n771 ) ;
  assign n773 = ( ~n514 & n739 ) | ( ~n514 & n772 ) | ( n739 & n772 ) ;
  assign n774 = ( ~n458 & n733 ) | ( ~n458 & n773 ) | ( n733 & n773 ) ;
  assign n775 = ( ~n399 & n737 ) | ( ~n399 & n774 ) | ( n737 & n774 ) ;
  assign n776 = ( ~n345 & n761 ) | ( ~n345 & n775 ) | ( n761 & n775 ) ;
  assign n777 = ( ~n302 & n757 ) | ( ~n302 & n776 ) | ( n757 & n776 ) ;
  assign n778 = ( ~n261 & n719 ) | ( ~n261 & n777 ) | ( n719 & n777 ) ;
  assign n779 = ( ~n217 & n749 ) | ( ~n217 & n778 ) | ( n749 & n778 ) ;
  assign n780 = ( ~n179 & n728 ) | ( ~n179 & n779 ) | ( n728 & n779 ) ;
  assign n781 = ( ~n144 & n734 ) | ( ~n144 & n780 ) | ( n734 & n780 ) ;
  assign n782 = ( ~n134 & n752 ) | ( ~n134 & n781 ) | ( n752 & n781 ) ;
  assign n783 = ( ~n136 & n745 ) | ( ~n136 & n782 ) | ( n745 & n782 ) ;
  assign n784 = n735 | n783 ;
  assign n785 = n759 | n784 ;
  assign n786 = ~n764 & n785 ;
  assign n787 = n784 & ~n786 ;
  assign n788 = ( n760 & n786 ) | ( n760 & ~n787 ) | ( n786 & ~n787 ) ;
  assign n789 = ( n762 & ~n767 ) | ( n762 & n785 ) | ( ~n767 & n785 ) ;
  assign n790 = ~n762 & n789 ;
  assign n791 = n790 ^ n768 ^ x2 ;
  assign n792 = n785 ^ n771 ^ n572 ;
  assign n793 = n785 & n792 ;
  assign n794 = n793 ^ n748 ^ x3 ;
  assign n795 = n772 ^ n514 ^ 1'b0 ;
  assign n796 = n785 & n795 ;
  assign n797 = n796 ^ n785 ^ n739 ;
  assign n798 = n785 ^ n773 ^ n458 ;
  assign n799 = n785 & n798 ;
  assign n800 = n799 ^ n727 ^ n682 ;
  assign n801 = n774 ^ n399 ^ 1'b0 ;
  assign n802 = n785 & n801 ;
  assign n803 = n802 ^ n785 ^ n737 ;
  assign n804 = n785 ^ n775 ^ n345 ;
  assign n805 = n785 & n804 ;
  assign n806 = n805 ^ n755 ^ n684 ;
  assign n807 = n776 ^ n302 ^ 1'b0 ;
  assign n808 = n785 & n807 ;
  assign n809 = n808 ^ n785 ^ n757 ;
  assign n810 = n785 ^ n777 ^ n261 ;
  assign n811 = n785 & n810 ;
  assign n812 = n811 ^ n718 ^ n653 ;
  assign n813 = n778 ^ n217 ^ 1'b0 ;
  assign n814 = n785 & n813 ;
  assign n815 = n814 ^ n785 ^ n749 ;
  assign n816 = n785 ^ n779 ^ n179 ;
  assign n817 = n785 & n816 ;
  assign n818 = n817 ^ n726 ^ n652 ;
  assign n819 = n780 ^ n144 ^ 1'b0 ;
  assign n820 = n785 & n819 ;
  assign n821 = n820 ^ n785 ^ n734 ;
  assign n822 = n785 ^ n781 ^ n134 ;
  assign n823 = n785 & n822 ;
  assign n824 = n823 ^ n747 ^ n696 ;
  assign n825 = x125 & n785 ;
  assign n826 = n788 ^ x1 ^ 1'b0 ;
  assign n827 = x123 | x124 ;
  assign n828 = ( x125 & ~n715 ) | ( x125 & n827 ) | ( ~n715 & n827 ) ;
  assign n829 = ( ~n716 & n825 ) | ( ~n716 & n828 ) | ( n825 & n828 ) ;
  assign n830 = ~n825 & n829 ;
  assign n831 = ~n745 & n782 ;
  assign n832 = n825 ^ n785 ^ x126 ;
  assign n833 = n830 | n832 ;
  assign n834 = x125 | n827 ;
  assign n835 = ( ~n745 & n782 ) | ( ~n745 & n785 ) | ( n782 & n785 ) ;
  assign n836 = ( n716 & n825 ) | ( n716 & ~n834 ) | ( n825 & ~n834 ) ;
  assign n837 = n833 & ~n836 ;
  assign n838 = n830 | n836 ;
  assign n839 = ( ~n640 & n826 ) | ( ~n640 & n837 ) | ( n826 & n837 ) ;
  assign n840 = ( ~n572 & n791 ) | ( ~n572 & n839 ) | ( n791 & n839 ) ;
  assign n841 = ( ~n514 & n794 ) | ( ~n514 & n840 ) | ( n794 & n840 ) ;
  assign n842 = ( ~n458 & n797 ) | ( ~n458 & n841 ) | ( n797 & n841 ) ;
  assign n843 = ( ~n399 & n800 ) | ( ~n399 & n842 ) | ( n800 & n842 ) ;
  assign n844 = ( ~n345 & n803 ) | ( ~n345 & n843 ) | ( n803 & n843 ) ;
  assign n845 = ( ~n302 & n806 ) | ( ~n302 & n844 ) | ( n806 & n844 ) ;
  assign n846 = ( ~n261 & n809 ) | ( ~n261 & n845 ) | ( n809 & n845 ) ;
  assign n847 = ( ~n217 & n812 ) | ( ~n217 & n846 ) | ( n812 & n846 ) ;
  assign n848 = ( ~n179 & n815 ) | ( ~n179 & n847 ) | ( n815 & n847 ) ;
  assign n849 = ( ~n144 & n818 ) | ( ~n144 & n848 ) | ( n818 & n848 ) ;
  assign n850 = ( ~n134 & n821 ) | ( ~n134 & n849 ) | ( n821 & n849 ) ;
  assign n851 = ( ~n136 & n824 ) | ( ~n136 & n850 ) | ( n824 & n850 ) ;
  assign n852 = ( ~n136 & n835 ) | ( ~n136 & n851 ) | ( n835 & n851 ) ;
  assign n853 = ( ~n831 & n851 ) | ( ~n831 & n852 ) | ( n851 & n852 ) ;
  assign n854 = ( n745 & ~n785 ) | ( n745 & n853 ) | ( ~n785 & n853 ) ;
  assign n855 = ( ~n745 & n785 ) | ( ~n745 & n853 ) | ( n785 & n853 ) ;
  assign n856 = n782 & ~n855 ;
  assign n857 = ( n136 & n745 ) | ( n136 & n782 ) | ( n745 & n782 ) ;
  assign n858 = ( n853 & ~n856 ) | ( n853 & n857 ) | ( ~n856 & n857 ) ;
  assign n859 = n854 | n858 ;
  assign n860 = n859 ^ n839 ^ n572 ;
  assign n861 = n859 & n860 ;
  assign n862 = n859 ^ n848 ^ n144 ;
  assign n863 = n859 & n862 ;
  assign n864 = n863 ^ n817 ^ n728 ;
  assign n865 = n859 ^ n844 ^ n302 ;
  assign n866 = n859 & n865 ;
  assign n867 = n866 ^ n805 ^ n761 ;
  assign n868 = n859 ^ n842 ^ n399 ;
  assign n869 = n859 & n868 ;
  assign n870 = n869 ^ n799 ^ n733 ;
  assign n871 = n859 ^ n840 ^ n514 ;
  assign n872 = n859 & n871 ;
  assign n873 = n827 & n859 ;
  assign n874 = n872 ^ n793 ^ n763 ;
  assign n875 = n861 ^ n790 ^ n769 ;
  assign n876 = n859 ^ n846 ^ n217 ;
  assign n877 = n859 & n876 ;
  assign n878 = n859 ^ n837 ^ n640 ;
  assign n879 = n877 ^ n811 ^ n719 ;
  assign n880 = n859 & n878 ;
  assign n881 = n841 ^ n458 ^ 1'b0 ;
  assign n882 = n880 ^ n788 ^ x1 ;
  assign n883 = n843 ^ n345 ^ 1'b0 ;
  assign n884 = n845 ^ n261 ^ 1'b0 ;
  assign n885 = n859 & n884 ;
  assign n886 = n847 ^ n179 ^ 1'b0 ;
  assign n887 = n859 & n886 ;
  assign n888 = n887 ^ n859 ^ n815 ;
  assign n889 = n849 ^ n134 ^ 1'b0 ;
  assign n890 = n885 ^ n859 ^ n809 ;
  assign n891 = n859 & n883 ;
  assign n892 = n891 ^ n859 ^ n803 ;
  assign n893 = n859 & n881 ;
  assign n894 = n893 ^ n859 ^ n797 ;
  assign n895 = n838 & n859 ;
  assign n896 = n785 & ~n858 ;
  assign n897 = n895 ^ n859 ^ n832 ;
  assign n898 = n859 & n889 ;
  assign n899 = n898 ^ n859 ^ n821 ;
  assign n900 = ( n859 & ~n873 ) | ( n859 & n896 ) | ( ~n873 & n896 ) ;
  assign n901 = ( ~x123 & n785 ) | ( ~x123 & n859 ) | ( n785 & n859 ) ;
  assign n902 = x121 | x122 ;
  assign n903 = ( x123 & n785 ) | ( x123 & ~n902 ) | ( n785 & ~n902 ) ;
  assign n904 = n901 & n903 ;
  assign n905 = x123 & n859 ;
  assign n906 = ( x123 & ~n784 ) | ( x123 & n902 ) | ( ~n784 & n902 ) ;
  assign n907 = n905 ^ n859 ^ x124 ;
  assign n908 = ( n824 & n850 ) | ( n824 & ~n859 ) | ( n850 & ~n859 ) ;
  assign n909 = ( n136 & n824 ) | ( n136 & n850 ) | ( n824 & n850 ) ;
  assign n910 = ~n850 & n909 ;
  assign n911 = ( ~n908 & n909 ) | ( ~n908 & n910 ) | ( n909 & n910 ) ;
  assign n912 = n900 ^ x125 ^ 1'b0 ;
  assign n913 = ( ~n785 & n905 ) | ( ~n785 & n906 ) | ( n905 & n906 ) ;
  assign n914 = ~n905 & n913 ;
  assign n915 = n907 | n914 ;
  assign n916 = ~n904 & n915 ;
  assign n917 = ( ~n716 & n912 ) | ( ~n716 & n916 ) | ( n912 & n916 ) ;
  assign n918 = ( ~n640 & n897 ) | ( ~n640 & n917 ) | ( n897 & n917 ) ;
  assign n919 = ~n824 & n850 ;
  assign n920 = ( ~n572 & n882 ) | ( ~n572 & n918 ) | ( n882 & n918 ) ;
  assign n921 = ( ~n824 & n850 ) | ( ~n824 & n859 ) | ( n850 & n859 ) ;
  assign n922 = ( n899 & ~n919 ) | ( n899 & n921 ) | ( ~n919 & n921 ) ;
  assign n923 = n904 | n914 ;
  assign n924 = ( ~n514 & n875 ) | ( ~n514 & n920 ) | ( n875 & n920 ) ;
  assign n925 = ( ~n458 & n874 ) | ( ~n458 & n924 ) | ( n874 & n924 ) ;
  assign n926 = ( ~n399 & n894 ) | ( ~n399 & n925 ) | ( n894 & n925 ) ;
  assign n927 = ( ~n345 & n870 ) | ( ~n345 & n926 ) | ( n870 & n926 ) ;
  assign n928 = ( ~n302 & n892 ) | ( ~n302 & n927 ) | ( n892 & n927 ) ;
  assign n929 = ( ~n261 & n867 ) | ( ~n261 & n928 ) | ( n867 & n928 ) ;
  assign n930 = ( ~n217 & n890 ) | ( ~n217 & n929 ) | ( n890 & n929 ) ;
  assign n931 = ( ~n179 & n879 ) | ( ~n179 & n930 ) | ( n879 & n930 ) ;
  assign n932 = ( ~n144 & n888 ) | ( ~n144 & n931 ) | ( n888 & n931 ) ;
  assign n933 = ( ~n134 & n864 ) | ( ~n134 & n932 ) | ( n864 & n932 ) ;
  assign n934 = ( ~x30 & n922 ) | ( ~x30 & n933 ) | ( n922 & n933 ) ;
  assign n935 = ~n136 & n934 ;
  assign n936 = n917 ^ n640 ^ 1'b0 ;
  assign n937 = ( n824 & ~n859 ) | ( n824 & n911 ) | ( ~n859 & n911 ) ;
  assign n938 = n899 & n933 ;
  assign n939 = n935 | n938 ;
  assign n940 = ( ~n911 & n937 ) | ( ~n911 & n939 ) | ( n937 & n939 ) ;
  assign n941 = n911 | n940 ;
  assign n942 = n929 ^ n217 ^ 1'b0 ;
  assign n943 = n941 & n942 ;
  assign n944 = n923 & n941 ;
  assign n945 = n943 ^ n941 ^ n890 ;
  assign n946 = n936 & n941 ;
  assign n947 = n941 ^ n932 ^ n134 ;
  assign n948 = n941 & n947 ;
  assign n949 = n941 ^ n926 ^ n345 ;
  assign n950 = n941 ^ n928 ^ n261 ;
  assign n951 = n941 & n950 ;
  assign n952 = n951 ^ n866 ^ n806 ;
  assign n953 = n941 & n949 ;
  assign n954 = n948 ^ n863 ^ n818 ;
  assign n955 = n941 ^ n920 ^ n514 ;
  assign n956 = n941 & n955 ;
  assign n957 = n956 ^ n861 ^ n791 ;
  assign n958 = n941 ^ n918 ^ n572 ;
  assign n959 = n941 ^ n924 ^ n458 ;
  assign n960 = n941 & n959 ;
  assign n961 = n953 ^ n869 ^ n800 ;
  assign n962 = n941 & n958 ;
  assign n963 = n962 ^ n880 ^ n826 ;
  assign n964 = n960 ^ n872 ^ n794 ;
  assign n965 = n946 ^ n941 ^ n897 ;
  assign n966 = n944 ^ n941 ^ n907 ;
  assign n967 = x119 | x120 ;
  assign n968 = ~n902 & n941 ;
  assign n969 = n939 & ~n968 ;
  assign n970 = ( x121 & ~n853 ) | ( x121 & n967 ) | ( ~n853 & n967 ) ;
  assign n971 = ( n859 & ~n911 ) | ( n859 & n968 ) | ( ~n911 & n968 ) ;
  assign n972 = ( n968 & ~n969 ) | ( n968 & n971 ) | ( ~n969 & n971 ) ;
  assign n973 = n925 ^ n399 ^ 1'b0 ;
  assign n974 = n972 ^ x123 ^ 1'b0 ;
  assign n975 = n941 & n973 ;
  assign n976 = x121 & n941 ;
  assign n977 = n941 ^ n916 ^ n716 ;
  assign n978 = n975 ^ n941 ^ n894 ;
  assign n979 = ( ~n859 & n970 ) | ( ~n859 & n976 ) | ( n970 & n976 ) ;
  assign n980 = n976 ^ n941 ^ x122 ;
  assign n981 = ~n976 & n979 ;
  assign n982 = n980 | n981 ;
  assign n983 = n941 & n977 ;
  assign n984 = n983 ^ n900 ^ x125 ;
  assign n985 = n931 ^ n144 ^ 1'b0 ;
  assign n986 = n941 & n985 ;
  assign n987 = ( n899 & ~n933 ) | ( n899 & n941 ) | ( ~n933 & n941 ) ;
  assign n988 = ( n933 & n938 ) | ( n933 & ~n941 ) | ( n938 & ~n941 ) ;
  assign n989 = ( n136 & n899 ) | ( n136 & n933 ) | ( n899 & n933 ) ;
  assign n990 = n899 & ~n933 ;
  assign n991 = n986 ^ n941 ^ n888 ;
  assign n992 = ( ~x121 & n859 ) | ( ~x121 & n941 ) | ( n859 & n941 ) ;
  assign n993 = n927 ^ n302 ^ 1'b0 ;
  assign n994 = ( x121 & n859 ) | ( x121 & ~n967 ) | ( n859 & ~n967 ) ;
  assign n995 = ~n988 & n989 ;
  assign n996 = n992 & n994 ;
  assign n997 = n982 & ~n996 ;
  assign n998 = ( ~n785 & n974 ) | ( ~n785 & n997 ) | ( n974 & n997 ) ;
  assign n999 = ( ~n716 & n966 ) | ( ~n716 & n998 ) | ( n966 & n998 ) ;
  assign n1000 = n941 & n993 ;
  assign n1001 = n1000 ^ n941 ^ n892 ;
  assign n1002 = ( ~n640 & n984 ) | ( ~n640 & n999 ) | ( n984 & n999 ) ;
  assign n1003 = ( ~n572 & n965 ) | ( ~n572 & n1002 ) | ( n965 & n1002 ) ;
  assign n1004 = n998 ^ n716 ^ 1'b0 ;
  assign n1005 = ( ~n514 & n963 ) | ( ~n514 & n1003 ) | ( n963 & n1003 ) ;
  assign n1006 = n981 | n996 ;
  assign n1007 = ( ~n458 & n957 ) | ( ~n458 & n1005 ) | ( n957 & n1005 ) ;
  assign n1008 = ( ~n399 & n964 ) | ( ~n399 & n1007 ) | ( n964 & n1007 ) ;
  assign n1009 = ( n954 & n987 ) | ( n954 & ~n990 ) | ( n987 & ~n990 ) ;
  assign n1010 = n1008 ^ n345 ^ 1'b0 ;
  assign n1011 = ( ~n345 & n978 ) | ( ~n345 & n1008 ) | ( n978 & n1008 ) ;
  assign n1012 = ( ~n302 & n961 ) | ( ~n302 & n1011 ) | ( n961 & n1011 ) ;
  assign n1013 = n941 ^ n930 ^ n179 ;
  assign n1014 = n1002 ^ n572 ^ 1'b0 ;
  assign n1015 = n941 & n1013 ;
  assign n1016 = n899 & ~n941 ;
  assign n1017 = n1015 ^ n877 ^ n812 ;
  assign n1018 = ( x114 & x115 ) | ( x114 & ~n1016 ) | ( x115 & ~n1016 ) ;
  assign n1019 = ( x117 & ~n1016 ) | ( x117 & n1018 ) | ( ~n1016 & n1018 ) ;
  assign n1020 = ( ~n261 & n1001 ) | ( ~n261 & n1012 ) | ( n1001 & n1012 ) ;
  assign n1021 = ( ~n217 & n952 ) | ( ~n217 & n1020 ) | ( n952 & n1020 ) ;
  assign n1022 = ( ~n179 & n945 ) | ( ~n179 & n1021 ) | ( n945 & n1021 ) ;
  assign n1023 = ( ~n144 & n1017 ) | ( ~n144 & n1022 ) | ( n1017 & n1022 ) ;
  assign n1024 = ( ~n134 & n991 ) | ( ~n134 & n1023 ) | ( n991 & n1023 ) ;
  assign n1025 = n954 & n1024 ;
  assign n1026 = n1016 | n1025 ;
  assign n1027 = ( ~n995 & n1019 ) | ( ~n995 & n1026 ) | ( n1019 & n1026 ) ;
  assign n1028 = ~n1026 & n1027 ;
  assign n1029 = ( n954 & n995 ) | ( n954 & ~n1016 ) | ( n995 & ~n1016 ) ;
  assign n1030 = n995 | n1025 ;
  assign n1031 = ( ~x30 & n1009 ) | ( ~x30 & n1024 ) | ( n1009 & n1024 ) ;
  assign n1032 = ~n136 & n1031 ;
  assign n1033 = n1030 | n1032 ;
  assign n1034 = n1016 | n1033 ;
  assign n1035 = n1014 & n1034 ;
  assign n1036 = n1021 ^ n179 ^ 1'b0 ;
  assign n1037 = ~n967 & n1034 ;
  assign n1038 = n1034 ^ n1022 ^ n144 ;
  assign n1039 = n1034 & n1038 ;
  assign n1040 = n1039 ^ n1015 ^ n879 ;
  assign n1041 = n1004 & n1034 ;
  assign n1042 = ( n136 & n954 ) | ( n136 & n1024 ) | ( n954 & n1024 ) ;
  assign n1043 = n1034 ^ n999 ^ n640 ;
  assign n1044 = n1034 ^ n1005 ^ n458 ;
  assign n1045 = n1035 ^ n1034 ^ n965 ;
  assign n1046 = n1034 & n1044 ;
  assign n1047 = n1023 ^ n134 ^ 1'b0 ;
  assign n1048 = n1034 ^ n1003 ^ n514 ;
  assign n1049 = n941 & ~n1033 ;
  assign n1050 = n1006 & n1034 ;
  assign n1051 = n1034 & n1043 ;
  assign n1052 = ( n1024 & n1025 ) | ( n1024 & ~n1034 ) | ( n1025 & ~n1034 ) ;
  assign n1053 = n1034 & n1036 ;
  assign n1054 = n1034 ^ n1011 ^ n302 ;
  assign n1055 = n1053 ^ n1034 ^ n945 ;
  assign n1056 = n1034 ^ n1020 ^ n217 ;
  assign n1057 = n1034 & n1048 ;
  assign n1058 = n1057 ^ n962 ^ n882 ;
  assign n1059 = n1029 & ~n1033 ;
  assign n1060 = ~n954 & n1024 ;
  assign n1061 = n1034 & n1056 ;
  assign n1062 = n1041 ^ n1034 ^ n966 ;
  assign n1063 = n1046 ^ n956 ^ n875 ;
  assign n1064 = n1034 & n1054 ;
  assign n1065 = n1061 ^ n951 ^ n867 ;
  assign n1066 = n1050 ^ n1034 ^ n980 ;
  assign n1067 = n1051 ^ n983 ^ n912 ;
  assign n1068 = n1012 ^ n261 ^ 1'b0 ;
  assign n1069 = n1064 ^ n953 ^ n870 ;
  assign n1070 = n1034 & n1047 ;
  assign n1071 = n1034 ^ n1007 ^ n399 ;
  assign n1072 = n1010 & n1034 ;
  assign n1073 = n1070 ^ n1034 ^ n991 ;
  assign n1074 = ( ~n954 & n1024 ) | ( ~n954 & n1034 ) | ( n1024 & n1034 ) ;
  assign n1075 = ( ~n1060 & n1073 ) | ( ~n1060 & n1074 ) | ( n1073 & n1074 ) ;
  assign n1076 = n1042 & ~n1052 ;
  assign n1077 = n1034 & n1068 ;
  assign n1078 = n1072 ^ n1034 ^ n978 ;
  assign n1079 = n1077 ^ n1034 ^ n1001 ;
  assign n1080 = n1034 ^ n997 ^ n785 ;
  assign n1081 = n1034 & n1071 ;
  assign n1082 = n1037 | n1049 ;
  assign n1083 = n1081 ^ n960 ^ n874 ;
  assign n1084 = n1034 & n1080 ;
  assign n1085 = x117 | x118 ;
  assign n1086 = x119 | n1085 ;
  assign n1087 = x119 & n1034 ;
  assign n1088 = n1087 ^ n1034 ^ x120 ;
  assign n1089 = ( x119 & ~n939 ) | ( x119 & n1085 ) | ( ~n939 & n1085 ) ;
  assign n1090 = n1084 ^ n972 ^ x123 ;
  assign n1091 = ( n941 & ~n1086 ) | ( n941 & n1087 ) | ( ~n1086 & n1087 ) ;
  assign n1092 = ( ~n941 & n1087 ) | ( ~n941 & n1089 ) | ( n1087 & n1089 ) ;
  assign n1093 = ~n1087 & n1092 ;
  assign n1094 = n1082 ^ x121 ^ 1'b0 ;
  assign n1095 = n1088 | n1093 ;
  assign n1096 = ~n1091 & n1095 ;
  assign n1097 = ( ~n859 & n1094 ) | ( ~n859 & n1096 ) | ( n1094 & n1096 ) ;
  assign n1098 = ( ~n785 & n1066 ) | ( ~n785 & n1097 ) | ( n1066 & n1097 ) ;
  assign n1099 = ( ~n716 & n1090 ) | ( ~n716 & n1098 ) | ( n1090 & n1098 ) ;
  assign n1100 = ( ~n640 & n1062 ) | ( ~n640 & n1099 ) | ( n1062 & n1099 ) ;
  assign n1101 = ( ~n572 & n1067 ) | ( ~n572 & n1100 ) | ( n1067 & n1100 ) ;
  assign n1102 = ( ~n514 & n1045 ) | ( ~n514 & n1101 ) | ( n1045 & n1101 ) ;
  assign n1103 = ( ~n458 & n1058 ) | ( ~n458 & n1102 ) | ( n1058 & n1102 ) ;
  assign n1104 = ( ~n399 & n1063 ) | ( ~n399 & n1103 ) | ( n1063 & n1103 ) ;
  assign n1105 = ( ~n345 & n1083 ) | ( ~n345 & n1104 ) | ( n1083 & n1104 ) ;
  assign n1106 = ( ~n302 & n1078 ) | ( ~n302 & n1105 ) | ( n1078 & n1105 ) ;
  assign n1107 = ( ~n261 & n1069 ) | ( ~n261 & n1106 ) | ( n1069 & n1106 ) ;
  assign n1108 = ( ~n217 & n1079 ) | ( ~n217 & n1107 ) | ( n1079 & n1107 ) ;
  assign n1109 = ( ~n179 & n1065 ) | ( ~n179 & n1108 ) | ( n1065 & n1108 ) ;
  assign n1110 = ( ~n144 & n1055 ) | ( ~n144 & n1109 ) | ( n1055 & n1109 ) ;
  assign n1111 = ( ~n134 & n1040 ) | ( ~n134 & n1110 ) | ( n1040 & n1110 ) ;
  assign n1112 = n1073 & n1111 ;
  assign n1113 = ( ~x30 & n1075 ) | ( ~x30 & n1111 ) | ( n1075 & n1111 ) ;
  assign n1114 = n1059 | n1112 ;
  assign n1115 = n1091 | n1093 ;
  assign n1116 = ~n136 & n1113 ;
  assign n1117 = n1114 | n1116 ;
  assign n1118 = n1076 | n1117 ;
  assign n1119 = n1118 ^ n1103 ^ n399 ;
  assign n1120 = n1105 ^ n302 ^ 1'b0 ;
  assign n1121 = n1118 ^ n1102 ^ n458 ;
  assign n1122 = n1118 & n1119 ;
  assign n1123 = n1122 ^ n1046 ^ n957 ;
  assign n1124 = n1118 & n1121 ;
  assign n1125 = n1124 ^ n1057 ^ n963 ;
  assign n1126 = n1118 ^ n1110 ^ n134 ;
  assign n1127 = n1118 & n1126 ;
  assign n1128 = n1127 ^ n1039 ^ n1017 ;
  assign n1129 = n1099 ^ n640 ^ 1'b0 ;
  assign n1130 = n1118 & n1120 ;
  assign n1131 = n1097 ^ n785 ^ 1'b0 ;
  assign n1132 = n1107 ^ n217 ^ 1'b0 ;
  assign n1133 = n1118 ^ n1108 ^ n179 ;
  assign n1134 = n1118 ^ n1106 ^ n261 ;
  assign n1135 = n1118 ^ n1104 ^ n345 ;
  assign n1136 = n1130 ^ n1118 ^ n1078 ;
  assign n1137 = ( x117 & n1032 ) | ( x117 & n1118 ) | ( n1032 & n1118 ) ;
  assign n1138 = ( n1028 & ~n1032 ) | ( n1028 & n1137 ) | ( ~n1032 & n1137 ) ;
  assign n1139 = n1118 ^ n1098 ^ n716 ;
  assign n1140 = n1118 ^ n1100 ^ n572 ;
  assign n1141 = n1118 & n1139 ;
  assign n1142 = ~n1137 & n1138 ;
  assign n1143 = n1109 ^ n144 ^ 1'b0 ;
  assign n1144 = n1101 ^ n514 ^ 1'b0 ;
  assign n1145 = n1115 & n1118 ;
  assign n1146 = n1118 & n1143 ;
  assign n1147 = n1118 & n1140 ;
  assign n1148 = n1145 ^ n1118 ^ n1088 ;
  assign n1149 = n1118 & n1135 ;
  assign n1150 = n1147 ^ n1051 ^ n984 ;
  assign n1151 = n1118 & n1134 ;
  assign n1152 = n1118 & n1144 ;
  assign n1153 = n1118 & n1132 ;
  assign n1154 = n1118 & n1129 ;
  assign n1155 = n1118 & n1131 ;
  assign n1156 = n1149 ^ n1081 ^ n964 ;
  assign n1157 = n1141 ^ n1084 ^ n974 ;
  assign n1158 = n1151 ^ n1064 ^ n961 ;
  assign n1159 = n1118 & n1133 ;
  assign n1160 = n1159 ^ n1061 ^ n952 ;
  assign n1161 = n1155 ^ n1118 ^ n1066 ;
  assign n1162 = n1154 ^ n1118 ^ n1062 ;
  assign n1163 = n1152 ^ n1118 ^ n1045 ;
  assign n1164 = n1153 ^ n1118 ^ n1079 ;
  assign n1165 = n1146 ^ n1118 ^ n1055 ;
  assign n1166 = ~n1085 & n1118 ;
  assign n1167 = ~x117 & n1118 ;
  assign n1168 = ( ~x117 & n1034 ) | ( ~x117 & n1118 ) | ( n1034 & n1118 ) ;
  assign n1169 = x114 | x115 ;
  assign n1170 = ( x117 & n1034 ) | ( x117 & ~n1169 ) | ( n1034 & ~n1169 ) ;
  assign n1171 = n1167 ^ x118 ^ 1'b0 ;
  assign n1172 = n1168 & n1170 ;
  assign n1173 = ( n1034 & n1059 ) | ( n1034 & ~n1076 ) | ( n1059 & ~n1076 ) ;
  assign n1174 = n1117 & ~n1166 ;
  assign n1175 = n1118 ^ n1096 ^ n859 ;
  assign n1176 = n1118 & n1175 ;
  assign n1177 = n1142 | n1171 ;
  assign n1178 = ~n1172 & n1177 ;
  assign n1179 = n1076 | n1112 ;
  assign n1180 = ( x112 & x113 ) | ( x112 & ~n1076 ) | ( x113 & ~n1076 ) ;
  assign n1181 = n1176 ^ n1082 ^ x121 ;
  assign n1182 = ( x114 & ~n1076 ) | ( x114 & n1180 ) | ( ~n1076 & n1180 ) ;
  assign n1183 = ( ~n1059 & n1179 ) | ( ~n1059 & n1182 ) | ( n1179 & n1182 ) ;
  assign n1184 = ( n1166 & n1173 ) | ( n1166 & ~n1174 ) | ( n1173 & ~n1174 ) ;
  assign n1185 = n1184 ^ x119 ^ 1'b0 ;
  assign n1186 = ( n1059 & n1073 ) | ( n1059 & ~n1076 ) | ( n1073 & ~n1076 ) ;
  assign n1187 = ( ~n941 & n1178 ) | ( ~n941 & n1185 ) | ( n1178 & n1185 ) ;
  assign n1188 = ( ~n859 & n1148 ) | ( ~n859 & n1187 ) | ( n1148 & n1187 ) ;
  assign n1189 = ( ~n785 & n1181 ) | ( ~n785 & n1188 ) | ( n1181 & n1188 ) ;
  assign n1190 = ( ~n716 & n1161 ) | ( ~n716 & n1189 ) | ( n1161 & n1189 ) ;
  assign n1191 = ( ~n640 & n1157 ) | ( ~n640 & n1190 ) | ( n1157 & n1190 ) ;
  assign n1192 = ~n1117 & n1186 ;
  assign n1193 = ( ~n572 & n1162 ) | ( ~n572 & n1191 ) | ( n1162 & n1191 ) ;
  assign n1194 = ( ~n514 & n1150 ) | ( ~n514 & n1193 ) | ( n1150 & n1193 ) ;
  assign n1195 = ( ~n458 & n1163 ) | ( ~n458 & n1194 ) | ( n1163 & n1194 ) ;
  assign n1196 = ( ~n399 & n1125 ) | ( ~n399 & n1195 ) | ( n1125 & n1195 ) ;
  assign n1197 = ( ~n345 & n1123 ) | ( ~n345 & n1196 ) | ( n1123 & n1196 ) ;
  assign n1198 = ( ~n302 & n1156 ) | ( ~n302 & n1197 ) | ( n1156 & n1197 ) ;
  assign n1199 = ~n1179 & n1183 ;
  assign n1200 = ( ~n261 & n1136 ) | ( ~n261 & n1198 ) | ( n1136 & n1198 ) ;
  assign n1201 = ( ~n217 & n1158 ) | ( ~n217 & n1200 ) | ( n1158 & n1200 ) ;
  assign n1202 = ( ~n179 & n1164 ) | ( ~n179 & n1201 ) | ( n1164 & n1201 ) ;
  assign n1203 = ( ~n144 & n1160 ) | ( ~n144 & n1202 ) | ( n1160 & n1202 ) ;
  assign n1204 = n1198 ^ n261 ^ 1'b0 ;
  assign n1205 = ( n136 & n1073 ) | ( n136 & n1111 ) | ( n1073 & n1111 ) ;
  assign n1206 = ( n1111 & n1112 ) | ( n1111 & ~n1118 ) | ( n1112 & ~n1118 ) ;
  assign n1207 = n1187 ^ n859 ^ 1'b0 ;
  assign n1208 = ( ~n1073 & n1111 ) | ( ~n1073 & n1118 ) | ( n1111 & n1118 ) ;
  assign n1209 = ~n1073 & n1111 ;
  assign n1210 = ( ~n134 & n1165 ) | ( ~n134 & n1203 ) | ( n1165 & n1203 ) ;
  assign n1211 = n1205 & ~n1206 ;
  assign n1212 = n1203 ^ n134 ^ 1'b0 ;
  assign n1213 = ( n1128 & n1208 ) | ( n1128 & ~n1209 ) | ( n1208 & ~n1209 ) ;
  assign n1214 = n1201 ^ n179 ^ 1'b0 ;
  assign n1215 = ( ~x30 & n1210 ) | ( ~x30 & n1213 ) | ( n1210 & n1213 ) ;
  assign n1216 = ~n136 & n1215 ;
  assign n1217 = n1128 & n1210 ;
  assign n1218 = n1216 | n1217 ;
  assign n1219 = n1211 | n1218 ;
  assign n1220 = n1192 | n1219 ;
  assign n1221 = n1220 ^ n1190 ^ n640 ;
  assign n1222 = n1220 & n1221 ;
  assign n1223 = n1222 ^ n1141 ^ n1090 ;
  assign n1224 = n1207 & n1220 ;
  assign n1225 = n1212 & n1220 ;
  assign n1226 = n1220 ^ n1202 ^ n144 ;
  assign n1227 = ~n1169 & n1220 ;
  assign n1228 = n1220 & n1226 ;
  assign n1229 = n1220 ^ n1196 ^ n345 ;
  assign n1230 = ( x114 & n1116 ) | ( x114 & n1220 ) | ( n1116 & n1220 ) ;
  assign n1231 = n1220 & n1229 ;
  assign n1232 = ( ~n1116 & n1199 ) | ( ~n1116 & n1230 ) | ( n1199 & n1230 ) ;
  assign n1233 = n1214 & n1220 ;
  assign n1234 = n1204 & n1220 ;
  assign n1235 = n1225 ^ n1220 ^ n1165 ;
  assign n1236 = n1220 ^ n1195 ^ n399 ;
  assign n1237 = n1234 ^ n1220 ^ n1136 ;
  assign n1238 = n1224 ^ n1220 ^ n1148 ;
  assign n1239 = n1228 ^ n1159 ^ n1065 ;
  assign n1240 = n1233 ^ n1220 ^ n1164 ;
  assign n1241 = ( n1192 & n1211 ) | ( n1192 & ~n1227 ) | ( n1211 & ~n1227 ) ;
  assign n1242 = ~n1230 & n1232 ;
  assign n1243 = n1231 ^ n1122 ^ n1063 ;
  assign n1244 = ( n1128 & ~n1210 ) | ( n1128 & n1220 ) | ( ~n1210 & n1220 ) ;
  assign n1245 = n1118 & ~n1218 ;
  assign n1246 = n1227 | n1245 ;
  assign n1247 = ( n1227 & ~n1241 ) | ( n1227 & n1246 ) | ( ~n1241 & n1246 ) ;
  assign n1248 = n1220 ^ n1188 ^ n785 ;
  assign n1249 = ~x114 & n1220 ;
  assign n1250 = n1220 & n1236 ;
  assign n1251 = n1128 & ~n1210 ;
  assign n1252 = n1250 ^ n1124 ^ n1058 ;
  assign n1253 = ( n136 & n1128 ) | ( n136 & n1210 ) | ( n1128 & n1210 ) ;
  assign n1254 = n1247 ^ x117 ^ 1'b0 ;
  assign n1255 = ( n1142 & ~n1172 ) | ( n1142 & n1220 ) | ( ~n1172 & n1220 ) ;
  assign n1256 = n1189 ^ n716 ^ 1'b0 ;
  assign n1257 = ~n1142 & n1255 ;
  assign n1258 = n1220 ^ n1200 ^ n217 ;
  assign n1259 = n1220 ^ n1178 ^ n941 ;
  assign n1260 = x112 | x113 ;
  assign n1261 = n1257 ^ n1167 ^ x118 ;
  assign n1262 = n1220 & n1259 ;
  assign n1263 = n1262 ^ n1184 ^ x119 ;
  assign n1264 = n1191 ^ n572 ^ 1'b0 ;
  assign n1265 = ( x114 & n1118 ) | ( x114 & ~n1260 ) | ( n1118 & ~n1260 ) ;
  assign n1266 = n1220 ^ n1193 ^ n514 ;
  assign n1267 = n1194 ^ n458 ^ 1'b0 ;
  assign n1268 = n1220 ^ n1197 ^ n302 ;
  assign n1269 = n1220 & n1256 ;
  assign n1270 = n1249 ^ x115 ^ 1'b0 ;
  assign n1271 = n1220 & n1264 ;
  assign n1272 = n1269 ^ n1220 ^ n1161 ;
  assign n1273 = n1220 & n1258 ;
  assign n1274 = ( ~x114 & n1118 ) | ( ~x114 & n1220 ) | ( n1118 & n1220 ) ;
  assign n1275 = ( n1210 & n1217 ) | ( n1210 & ~n1220 ) | ( n1217 & ~n1220 ) ;
  assign n1276 = n1220 & n1266 ;
  assign n1277 = n1242 | n1270 ;
  assign n1278 = n1265 & n1274 ;
  assign n1279 = n1271 ^ n1220 ^ n1162 ;
  assign n1280 = n1276 ^ n1147 ^ n1067 ;
  assign n1281 = n1277 & ~n1278 ;
  assign n1282 = ( ~n1034 & n1254 ) | ( ~n1034 & n1281 ) | ( n1254 & n1281 ) ;
  assign n1283 = n1220 & n1268 ;
  assign n1284 = n1220 & n1248 ;
  assign n1285 = ( ~n941 & n1261 ) | ( ~n941 & n1282 ) | ( n1261 & n1282 ) ;
  assign n1286 = n1284 ^ n1176 ^ n1094 ;
  assign n1287 = ( ~n859 & n1263 ) | ( ~n859 & n1285 ) | ( n1263 & n1285 ) ;
  assign n1288 = ( ~n785 & n1238 ) | ( ~n785 & n1287 ) | ( n1238 & n1287 ) ;
  assign n1289 = n1273 ^ n1151 ^ n1069 ;
  assign n1290 = ( ~n716 & n1286 ) | ( ~n716 & n1288 ) | ( n1286 & n1288 ) ;
  assign n1291 = ( ~n640 & n1272 ) | ( ~n640 & n1290 ) | ( n1272 & n1290 ) ;
  assign n1292 = ( n1235 & n1244 ) | ( n1235 & ~n1251 ) | ( n1244 & ~n1251 ) ;
  assign n1293 = ( ~n572 & n1223 ) | ( ~n572 & n1291 ) | ( n1223 & n1291 ) ;
  assign n1294 = n1253 & ~n1275 ;
  assign n1295 = n1293 ^ n514 ^ 1'b0 ;
  assign n1296 = ( ~n514 & n1279 ) | ( ~n514 & n1293 ) | ( n1279 & n1293 ) ;
  assign n1297 = n1290 ^ n640 ^ 1'b0 ;
  assign n1298 = n1220 & n1267 ;
  assign n1299 = n1287 ^ n785 ^ 1'b0 ;
  assign n1300 = n1298 ^ n1220 ^ n1163 ;
  assign n1301 = ( ~n458 & n1280 ) | ( ~n458 & n1296 ) | ( n1280 & n1296 ) ;
  assign n1302 = n1283 ^ n1149 ^ n1083 ;
  assign n1303 = n1301 ^ n399 ^ 1'b0 ;
  assign n1304 = ( ~n399 & n1300 ) | ( ~n399 & n1301 ) | ( n1300 & n1301 ) ;
  assign n1305 = ( ~n345 & n1252 ) | ( ~n345 & n1304 ) | ( n1252 & n1304 ) ;
  assign n1306 = ( ~n302 & n1243 ) | ( ~n302 & n1305 ) | ( n1243 & n1305 ) ;
  assign n1307 = ( ~n261 & n1302 ) | ( ~n261 & n1306 ) | ( n1302 & n1306 ) ;
  assign n1308 = ( ~n217 & n1237 ) | ( ~n217 & n1307 ) | ( n1237 & n1307 ) ;
  assign n1309 = ( ~n179 & n1289 ) | ( ~n179 & n1308 ) | ( n1289 & n1308 ) ;
  assign n1310 = ( ~n144 & n1240 ) | ( ~n144 & n1309 ) | ( n1240 & n1309 ) ;
  assign n1311 = ( ~n134 & n1239 ) | ( ~n134 & n1310 ) | ( n1239 & n1310 ) ;
  assign n1312 = n1235 & n1311 ;
  assign n1313 = ( n1128 & ~n1220 ) | ( n1128 & n1312 ) | ( ~n1220 & n1312 ) ;
  assign n1314 = ( ~x30 & n1292 ) | ( ~x30 & n1311 ) | ( n1292 & n1311 ) ;
  assign n1315 = ~n136 & n1314 ;
  assign n1316 = n1312 | n1315 ;
  assign n1317 = ( n1294 & ~n1313 ) | ( n1294 & n1316 ) | ( ~n1313 & n1316 ) ;
  assign n1318 = n1313 | n1317 ;
  assign n1319 = n1318 ^ n1310 ^ n134 ;
  assign n1320 = n1318 & n1319 ;
  assign n1321 = n1320 ^ n1228 ^ n1160 ;
  assign n1322 = ~n1260 & n1318 ;
  assign n1323 = ( n1220 & ~n1316 ) | ( n1220 & n1322 ) | ( ~n1316 & n1322 ) ;
  assign n1324 = n1294 & ~n1322 ;
  assign n1325 = ( n1322 & n1323 ) | ( n1322 & ~n1324 ) | ( n1323 & ~n1324 ) ;
  assign n1326 = n1318 ^ n1281 ^ n1034 ;
  assign n1327 = n1318 & n1326 ;
  assign n1328 = n1327 ^ n1247 ^ x117 ;
  assign n1329 = n1318 ^ n1282 ^ n941 ;
  assign n1330 = n1318 & n1329 ;
  assign n1331 = n1330 ^ n1257 ^ n1171 ;
  assign n1332 = n1318 ^ n1285 ^ n859 ;
  assign n1333 = n1318 & n1332 ;
  assign n1334 = n1333 ^ n1262 ^ n1185 ;
  assign n1335 = n1299 & n1318 ;
  assign n1336 = n1335 ^ n1318 ^ n1238 ;
  assign n1337 = n1318 ^ n1288 ^ n716 ;
  assign n1338 = n1318 & n1337 ;
  assign n1339 = n1338 ^ n1284 ^ n1181 ;
  assign n1340 = n1297 & n1318 ;
  assign n1341 = n1340 ^ n1318 ^ n1272 ;
  assign n1342 = n1318 ^ n1291 ^ n572 ;
  assign n1343 = n1318 & n1342 ;
  assign n1344 = n1343 ^ n1222 ^ n1157 ;
  assign n1345 = n1295 & n1318 ;
  assign n1346 = n1345 ^ n1318 ^ n1279 ;
  assign n1347 = n1318 ^ n1296 ^ n458 ;
  assign n1348 = n1318 & n1347 ;
  assign n1349 = n1348 ^ n1276 ^ n1150 ;
  assign n1350 = n1303 & n1318 ;
  assign n1351 = n1350 ^ n1318 ^ n1300 ;
  assign n1352 = n1318 ^ n1304 ^ n345 ;
  assign n1353 = n1318 & n1352 ;
  assign n1354 = n1353 ^ n1250 ^ n1125 ;
  assign n1355 = n1318 ^ n1305 ^ n302 ;
  assign n1356 = n1318 & n1355 ;
  assign n1357 = n1356 ^ n1231 ^ n1123 ;
  assign n1358 = n1318 ^ n1306 ^ n261 ;
  assign n1359 = n1318 & n1358 ;
  assign n1360 = ( n1242 & ~n1278 ) | ( n1242 & n1318 ) | ( ~n1278 & n1318 ) ;
  assign n1361 = ~n1242 & n1360 ;
  assign n1362 = n1361 ^ n1249 ^ x115 ;
  assign n1363 = n1359 ^ n1283 ^ n1156 ;
  assign n1364 = n1307 ^ n217 ^ 1'b0 ;
  assign n1365 = n1318 & n1364 ;
  assign n1366 = n1365 ^ n1318 ^ n1237 ;
  assign n1367 = n1318 ^ n1308 ^ n179 ;
  assign n1368 = n1318 & n1367 ;
  assign n1369 = n1368 ^ n1273 ^ n1158 ;
  assign n1370 = n1309 ^ n144 ^ 1'b0 ;
  assign n1371 = n1318 & n1370 ;
  assign n1372 = n1371 ^ n1318 ^ n1240 ;
  assign n1373 = ( n136 & n1235 ) | ( n136 & n1311 ) | ( n1235 & n1311 ) ;
  assign n1374 = ( n1311 & n1312 ) | ( n1311 & ~n1318 ) | ( n1312 & ~n1318 ) ;
  assign n1375 = n1373 & ~n1374 ;
  assign n1376 = x110 | x111 ;
  assign n1377 = ( ~x112 & n1220 ) | ( ~x112 & n1318 ) | ( n1220 & n1318 ) ;
  assign n1378 = ( x112 & n1220 ) | ( x112 & ~n1376 ) | ( n1220 & ~n1376 ) ;
  assign n1379 = n1377 & n1378 ;
  assign n1380 = x112 & n1318 ;
  assign n1381 = n1380 ^ n1318 ^ x113 ;
  assign n1382 = ( x112 & ~n1218 ) | ( x112 & n1376 ) | ( ~n1218 & n1376 ) ;
  assign n1383 = ( ~n1220 & n1380 ) | ( ~n1220 & n1382 ) | ( n1380 & n1382 ) ;
  assign n1384 = ~n1380 & n1383 ;
  assign n1385 = n1381 | n1384 ;
  assign n1386 = n1325 ^ x114 ^ 1'b0 ;
  assign n1387 = ~n1379 & n1385 ;
  assign n1388 = ( ~n1118 & n1386 ) | ( ~n1118 & n1387 ) | ( n1386 & n1387 ) ;
  assign n1389 = ( ~n1034 & n1362 ) | ( ~n1034 & n1388 ) | ( n1362 & n1388 ) ;
  assign n1390 = ( ~n941 & n1328 ) | ( ~n941 & n1389 ) | ( n1328 & n1389 ) ;
  assign n1391 = ( ~n859 & n1331 ) | ( ~n859 & n1390 ) | ( n1331 & n1390 ) ;
  assign n1392 = ( ~n785 & n1334 ) | ( ~n785 & n1391 ) | ( n1334 & n1391 ) ;
  assign n1393 = ( ~n716 & n1336 ) | ( ~n716 & n1392 ) | ( n1336 & n1392 ) ;
  assign n1394 = ( ~n640 & n1339 ) | ( ~n640 & n1393 ) | ( n1339 & n1393 ) ;
  assign n1395 = ( ~n572 & n1341 ) | ( ~n572 & n1394 ) | ( n1341 & n1394 ) ;
  assign n1396 = ( ~n514 & n1344 ) | ( ~n514 & n1395 ) | ( n1344 & n1395 ) ;
  assign n1397 = ( ~n458 & n1346 ) | ( ~n458 & n1396 ) | ( n1346 & n1396 ) ;
  assign n1398 = ( ~n399 & n1349 ) | ( ~n399 & n1397 ) | ( n1349 & n1397 ) ;
  assign n1399 = ( ~n345 & n1351 ) | ( ~n345 & n1398 ) | ( n1351 & n1398 ) ;
  assign n1400 = ( ~n302 & n1354 ) | ( ~n302 & n1399 ) | ( n1354 & n1399 ) ;
  assign n1401 = ( ~n261 & n1357 ) | ( ~n261 & n1400 ) | ( n1357 & n1400 ) ;
  assign n1402 = ( ~n217 & n1363 ) | ( ~n217 & n1401 ) | ( n1363 & n1401 ) ;
  assign n1403 = n1235 & ~n1318 ;
  assign n1404 = ( ~n179 & n1366 ) | ( ~n179 & n1402 ) | ( n1366 & n1402 ) ;
  assign n1405 = ( ~n144 & n1369 ) | ( ~n144 & n1404 ) | ( n1369 & n1404 ) ;
  assign n1406 = ( ~n134 & n1372 ) | ( ~n134 & n1405 ) | ( n1372 & n1405 ) ;
  assign n1407 = ( n1235 & ~n1311 ) | ( n1235 & n1318 ) | ( ~n1311 & n1318 ) ;
  assign n1408 = ( n136 & n1235 ) | ( n136 & ~n1311 ) | ( n1235 & ~n1311 ) ;
  assign n1409 = ( n1321 & n1407 ) | ( n1321 & ~n1408 ) | ( n1407 & ~n1408 ) ;
  assign n1410 = ~n136 & n1406 ;
  assign n1411 = ( ~n136 & n1409 ) | ( ~n136 & n1410 ) | ( n1409 & n1410 ) ;
  assign n1412 = n1375 | n1411 ;
  assign n1413 = n1379 | n1384 ;
  assign n1414 = n1321 & n1406 ;
  assign n1415 = n1412 | n1414 ;
  assign n1416 = n1403 | n1415 ;
  assign n1417 = n1416 ^ n1399 ^ n302 ;
  assign n1418 = n1416 & n1417 ;
  assign n1419 = n1418 ^ n1353 ^ n1252 ;
  assign n1420 = n1413 & n1416 ;
  assign n1421 = n1420 ^ n1416 ^ n1381 ;
  assign n1422 = n1416 ^ n1400 ^ n261 ;
  assign n1423 = n1416 ^ n1390 ^ n859 ;
  assign n1424 = n1416 & n1423 ;
  assign n1425 = n1424 ^ n1330 ^ n1261 ;
  assign n1426 = n1416 & n1422 ;
  assign n1427 = n1426 ^ n1356 ^ n1243 ;
  assign n1428 = n1416 ^ n1401 ^ n217 ;
  assign n1429 = n1416 & n1428 ;
  assign n1430 = n1429 ^ n1359 ^ n1302 ;
  assign n1431 = n1402 ^ n179 ^ 1'b0 ;
  assign n1432 = n1416 & n1431 ;
  assign n1433 = n1432 ^ n1416 ^ n1366 ;
  assign n1434 = n1416 ^ n1404 ^ n144 ;
  assign n1435 = n1416 & n1434 ;
  assign n1436 = n1435 ^ n1368 ^ n1289 ;
  assign n1437 = n1416 ^ n1387 ^ n1118 ;
  assign n1438 = n1416 ^ n1393 ^ n640 ;
  assign n1439 = n1398 ^ n345 ^ 1'b0 ;
  assign n1440 = n1392 ^ n716 ^ 1'b0 ;
  assign n1441 = n1405 ^ n134 ^ 1'b0 ;
  assign n1442 = n1416 ^ n1389 ^ n941 ;
  assign n1443 = n1416 ^ n1388 ^ n1034 ;
  assign n1444 = n1416 & n1443 ;
  assign n1445 = n1416 & n1438 ;
  assign n1446 = n1445 ^ n1338 ^ n1286 ;
  assign n1447 = ~n1376 & n1416 ;
  assign n1448 = ( n1321 & n1375 ) | ( n1321 & ~n1403 ) | ( n1375 & ~n1403 ) ;
  assign n1449 = n1416 & n1437 ;
  assign n1450 = ~n1415 & n1448 ;
  assign n1451 = n1416 & n1440 ;
  assign n1452 = n1416 ^ n1391 ^ n785 ;
  assign n1453 = n1416 ^ n1397 ^ n399 ;
  assign n1454 = n1416 & n1442 ;
  assign n1455 = n1449 ^ n1325 ^ x114 ;
  assign n1456 = n1416 & n1453 ;
  assign n1457 = n1416 ^ n1395 ^ n514 ;
  assign n1458 = n1416 & n1457 ;
  assign n1459 = n1454 ^ n1327 ^ n1254 ;
  assign n1460 = ( n1321 & ~n1406 ) | ( n1321 & n1416 ) | ( ~n1406 & n1416 ) ;
  assign n1461 = n1416 & n1452 ;
  assign n1462 = n1461 ^ n1333 ^ n1263 ;
  assign n1463 = n1394 ^ n572 ^ 1'b0 ;
  assign n1464 = n1416 & n1463 ;
  assign n1465 = n1464 ^ n1416 ^ n1341 ;
  assign n1466 = ( n136 & n1321 ) | ( n136 & n1406 ) | ( n1321 & n1406 ) ;
  assign n1467 = n1396 ^ n458 ^ 1'b0 ;
  assign n1468 = n1416 & n1467 ;
  assign n1469 = n1468 ^ n1416 ^ n1346 ;
  assign n1470 = ( n1406 & n1414 ) | ( n1406 & ~n1416 ) | ( n1414 & ~n1416 ) ;
  assign n1471 = n1416 & n1439 ;
  assign n1472 = ( x106 & x107 ) | ( x106 & ~n1403 ) | ( x107 & ~n1403 ) ;
  assign n1473 = n1471 ^ n1416 ^ n1351 ;
  assign n1474 = n1466 & ~n1470 ;
  assign n1475 = ( x108 & ~n1403 ) | ( x108 & n1472 ) | ( ~n1403 & n1472 ) ;
  assign n1476 = n1444 ^ n1361 ^ n1270 ;
  assign n1477 = n1456 ^ n1348 ^ n1280 ;
  assign n1478 = n1458 ^ n1343 ^ n1223 ;
  assign n1479 = n1375 | n1403 ;
  assign n1480 = n1318 & ~n1415 ;
  assign n1481 = n1321 & ~n1406 ;
  assign n1482 = n1416 & n1441 ;
  assign n1483 = n1451 ^ n1416 ^ n1336 ;
  assign n1484 = n1482 ^ n1416 ^ n1372 ;
  assign n1485 = ( n1460 & ~n1481 ) | ( n1460 & n1484 ) | ( ~n1481 & n1484 ) ;
  assign n1486 = ( ~n1414 & n1475 ) | ( ~n1414 & n1479 ) | ( n1475 & n1479 ) ;
  assign n1487 = ~n1479 & n1486 ;
  assign n1488 = n1447 | n1480 ;
  assign n1489 = x108 | x109 ;
  assign n1490 = x110 & n1416 ;
  assign n1491 = x110 | n1489 ;
  assign n1492 = ( n1318 & n1490 ) | ( n1318 & ~n1491 ) | ( n1490 & ~n1491 ) ;
  assign n1493 = ( x110 & ~n1316 ) | ( x110 & n1489 ) | ( ~n1316 & n1489 ) ;
  assign n1494 = ( ~n1318 & n1490 ) | ( ~n1318 & n1493 ) | ( n1490 & n1493 ) ;
  assign n1495 = n1490 ^ n1416 ^ x111 ;
  assign n1496 = n1488 ^ x112 ^ 1'b0 ;
  assign n1497 = ~n1490 & n1494 ;
  assign n1498 = n1495 | n1497 ;
  assign n1499 = ~n1492 & n1498 ;
  assign n1500 = ( ~n1220 & n1496 ) | ( ~n1220 & n1499 ) | ( n1496 & n1499 ) ;
  assign n1501 = ( ~n1118 & n1421 ) | ( ~n1118 & n1500 ) | ( n1421 & n1500 ) ;
  assign n1502 = ( ~n1034 & n1455 ) | ( ~n1034 & n1501 ) | ( n1455 & n1501 ) ;
  assign n1503 = n941 & n1502 ;
  assign n1504 = ( n1476 & n1502 ) | ( n1476 & ~n1503 ) | ( n1502 & ~n1503 ) ;
  assign n1505 = n941 & ~n1502 ;
  assign n1506 = ( n859 & ~n1504 ) | ( n859 & n1505 ) | ( ~n1504 & n1505 ) ;
  assign n1507 = ( ~n859 & n1504 ) | ( ~n859 & n1505 ) | ( n1504 & n1505 ) ;
  assign n1508 = ~n1505 & n1507 ;
  assign n1509 = n859 & n1506 ;
  assign n1510 = ( n1459 & n1508 ) | ( n1459 & ~n1509 ) | ( n1508 & ~n1509 ) ;
  assign n1511 = ~n1509 & n1510 ;
  assign n1512 = ( ~n785 & n1425 ) | ( ~n785 & n1511 ) | ( n1425 & n1511 ) ;
  assign n1513 = ( ~n716 & n1462 ) | ( ~n716 & n1512 ) | ( n1462 & n1512 ) ;
  assign n1514 = ( ~n640 & n1483 ) | ( ~n640 & n1513 ) | ( n1483 & n1513 ) ;
  assign n1515 = ( ~n572 & n1446 ) | ( ~n572 & n1514 ) | ( n1446 & n1514 ) ;
  assign n1516 = ( ~n514 & n1465 ) | ( ~n514 & n1515 ) | ( n1465 & n1515 ) ;
  assign n1517 = ( ~n458 & n1478 ) | ( ~n458 & n1516 ) | ( n1478 & n1516 ) ;
  assign n1518 = ( ~n399 & n1469 ) | ( ~n399 & n1517 ) | ( n1469 & n1517 ) ;
  assign n1519 = n1513 ^ n640 ^ 1'b0 ;
  assign n1520 = ( ~n345 & n1477 ) | ( ~n345 & n1518 ) | ( n1477 & n1518 ) ;
  assign n1521 = ( ~n302 & n1473 ) | ( ~n302 & n1520 ) | ( n1473 & n1520 ) ;
  assign n1522 = ( ~n261 & n1419 ) | ( ~n261 & n1521 ) | ( n1419 & n1521 ) ;
  assign n1523 = ( ~n217 & n1427 ) | ( ~n217 & n1522 ) | ( n1427 & n1522 ) ;
  assign n1524 = ( ~n179 & n1430 ) | ( ~n179 & n1523 ) | ( n1430 & n1523 ) ;
  assign n1525 = ( ~n144 & n1433 ) | ( ~n144 & n1524 ) | ( n1433 & n1524 ) ;
  assign n1526 = n1492 | n1497 ;
  assign n1527 = ( ~n134 & n1436 ) | ( ~n134 & n1525 ) | ( n1436 & n1525 ) ;
  assign n1528 = n1520 ^ n302 ^ 1'b0 ;
  assign n1529 = n1484 & n1527 ;
  assign n1530 = ( ~x30 & n1485 ) | ( ~x30 & n1527 ) | ( n1485 & n1527 ) ;
  assign n1531 = ~n136 & n1530 ;
  assign n1532 = n1474 | n1529 ;
  assign n1533 = n1531 | n1532 ;
  assign n1534 = n1450 | n1533 ;
  assign n1535 = n1519 & n1534 ;
  assign n1536 = n1534 ^ n1525 ^ n134 ;
  assign n1537 = n1528 & n1534 ;
  assign n1538 = n1526 & n1534 ;
  assign n1539 = n1534 ^ n1522 ^ n217 ;
  assign n1540 = n1515 ^ n514 ^ 1'b0 ;
  assign n1541 = n1534 ^ n1512 ^ n716 ;
  assign n1542 = n1534 & n1541 ;
  assign n1543 = n1537 ^ n1534 ^ n1473 ;
  assign n1544 = n1535 ^ n1534 ^ n1483 ;
  assign n1545 = n1534 & n1539 ;
  assign n1546 = n1534 & n1540 ;
  assign n1547 = n1542 ^ n1461 ^ n1334 ;
  assign n1548 = n1545 ^ n1426 ^ n1357 ;
  assign n1549 = n1534 ^ n1502 ^ n941 ;
  assign n1550 = n1534 & n1549 ;
  assign n1551 = n1508 | n1510 ;
  assign n1552 = n1550 ^ n1444 ^ n1362 ;
  assign n1553 = n1546 ^ n1534 ^ n1465 ;
  assign n1554 = ( n1508 & ~n1509 ) | ( n1508 & n1534 ) | ( ~n1509 & n1534 ) ;
  assign n1555 = ~n1508 & n1554 ;
  assign n1556 = n1555 ^ n1454 ^ n1328 ;
  assign n1557 = n1534 & n1536 ;
  assign n1558 = n1557 ^ n1435 ^ n1369 ;
  assign n1559 = n1538 ^ n1534 ^ n1495 ;
  assign n1560 = n1534 ^ n1521 ^ n261 ;
  assign n1561 = n1517 ^ n399 ^ 1'b0 ;
  assign n1562 = n1500 ^ n1118 ^ 1'b0 ;
  assign n1563 = n1534 ^ n1501 ^ n1034 ;
  assign n1564 = n1534 ^ n1514 ^ n572 ;
  assign n1565 = n1534 & n1561 ;
  assign n1566 = n1565 ^ n1534 ^ n1469 ;
  assign n1567 = n1534 ^ n1518 ^ n345 ;
  assign n1568 = n1534 & n1567 ;
  assign n1569 = n1534 & n1562 ;
  assign n1570 = n1511 ^ n1425 ^ n785 ;
  assign n1571 = n1569 ^ n1534 ^ n1421 ;
  assign n1572 = n1534 ^ n1516 ^ n458 ;
  assign n1573 = n1534 & n1560 ;
  assign n1574 = n1534 ^ n1523 ^ n179 ;
  assign n1575 = n1534 & n1574 ;
  assign n1576 = n1425 | n1570 ;
  assign n1577 = n1576 ^ n1551 ^ n785 ;
  assign n1578 = n1524 ^ n144 ^ 1'b0 ;
  assign n1579 = n1534 & n1578 ;
  assign n1580 = ( x103 & x104 ) | ( x103 & ~n1450 ) | ( x104 & ~n1450 ) ;
  assign n1581 = ( x108 & n1411 ) | ( x108 & n1534 ) | ( n1411 & n1534 ) ;
  assign n1582 = ( ~n1411 & n1487 ) | ( ~n1411 & n1581 ) | ( n1487 & n1581 ) ;
  assign n1583 = n1579 ^ n1534 ^ n1433 ;
  assign n1584 = ~n1581 & n1582 ;
  assign n1585 = ( x106 & ~n1450 ) | ( x106 & n1580 ) | ( ~n1450 & n1580 ) ;
  assign n1586 = n1534 & ~n1577 ;
  assign n1587 = n1568 ^ n1456 ^ n1349 ;
  assign n1588 = n1575 ^ n1429 ^ n1363 ;
  assign n1589 = n1534 & n1572 ;
  assign n1590 = n1589 ^ n1458 ^ n1344 ;
  assign n1591 = n1534 & n1564 ;
  assign n1592 = n1591 ^ n1445 ^ n1339 ;
  assign n1593 = n1534 ^ n1499 ^ n1220 ;
  assign n1594 = n785 & ~n1551 ;
  assign n1595 = ( n1416 & ~n1450 ) | ( n1416 & n1474 ) | ( ~n1450 & n1474 ) ;
  assign n1596 = ( ~n1450 & n1474 ) | ( ~n1450 & n1484 ) | ( n1474 & n1484 ) ;
  assign n1597 = n1450 | n1529 ;
  assign n1598 = n1534 & n1593 ;
  assign n1599 = n1598 ^ n1488 ^ x112 ;
  assign n1600 = ( ~n1484 & n1527 ) | ( ~n1484 & n1534 ) | ( n1527 & n1534 ) ;
  assign n1601 = ( n136 & n1484 ) | ( n136 & n1527 ) | ( n1484 & n1527 ) ;
  assign n1602 = ~n1484 & n1527 ;
  assign n1603 = ( n785 & n1534 ) | ( n785 & ~n1551 ) | ( n1534 & ~n1551 ) ;
  assign n1604 = ~n1489 & n1534 ;
  assign n1605 = n1533 & ~n1604 ;
  assign n1606 = ( n1595 & n1604 ) | ( n1595 & ~n1605 ) | ( n1604 & ~n1605 ) ;
  assign n1607 = n1573 ^ n1418 ^ n1354 ;
  assign n1608 = ( n1425 & ~n1594 ) | ( n1425 & n1603 ) | ( ~n1594 & n1603 ) ;
  assign n1609 = ( ~n1474 & n1585 ) | ( ~n1474 & n1597 ) | ( n1585 & n1597 ) ;
  assign n1610 = n1534 & n1563 ;
  assign n1611 = ( n1558 & n1600 ) | ( n1558 & ~n1602 ) | ( n1600 & ~n1602 ) ;
  assign n1612 = n1610 ^ n1449 ^ n1386 ;
  assign n1613 = ~n1597 & n1609 ;
  assign n1614 = ( n1527 & n1529 ) | ( n1527 & ~n1534 ) | ( n1529 & ~n1534 ) ;
  assign n1615 = n1601 & ~n1614 ;
  assign n1616 = ~n1533 & n1596 ;
  assign n1617 = ( ~n1534 & n1586 ) | ( ~n1534 & n1608 ) | ( n1586 & n1608 ) ;
  assign n1618 = n1606 ^ x110 ^ 1'b0 ;
  assign n1619 = x106 | x107 ;
  assign n1620 = ( x108 & n1416 ) | ( x108 & ~n1619 ) | ( n1416 & ~n1619 ) ;
  assign n1621 = ( ~x108 & n1416 ) | ( ~x108 & n1534 ) | ( n1416 & n1534 ) ;
  assign n1622 = n1620 & n1621 ;
  assign n1623 = ~x108 & n1534 ;
  assign n1624 = n1623 ^ x109 ^ 1'b0 ;
  assign n1625 = n1584 | n1624 ;
  assign n1626 = ~n1622 & n1625 ;
  assign n1627 = ( ~n1318 & n1618 ) | ( ~n1318 & n1626 ) | ( n1618 & n1626 ) ;
  assign n1628 = ( ~n1220 & n1559 ) | ( ~n1220 & n1627 ) | ( n1559 & n1627 ) ;
  assign n1629 = ( ~n1118 & n1599 ) | ( ~n1118 & n1628 ) | ( n1599 & n1628 ) ;
  assign n1630 = ( ~n1034 & n1571 ) | ( ~n1034 & n1629 ) | ( n1571 & n1629 ) ;
  assign n1631 = ( ~n941 & n1612 ) | ( ~n941 & n1630 ) | ( n1612 & n1630 ) ;
  assign n1632 = ( ~n859 & n1552 ) | ( ~n859 & n1631 ) | ( n1552 & n1631 ) ;
  assign n1633 = ( ~n785 & n1556 ) | ( ~n785 & n1632 ) | ( n1556 & n1632 ) ;
  assign n1634 = ( ~n716 & n1617 ) | ( ~n716 & n1633 ) | ( n1617 & n1633 ) ;
  assign n1635 = ( ~n640 & n1547 ) | ( ~n640 & n1634 ) | ( n1547 & n1634 ) ;
  assign n1636 = ( ~n572 & n1544 ) | ( ~n572 & n1635 ) | ( n1544 & n1635 ) ;
  assign n1637 = ( ~n514 & n1592 ) | ( ~n514 & n1636 ) | ( n1592 & n1636 ) ;
  assign n1638 = ( ~n458 & n1553 ) | ( ~n458 & n1637 ) | ( n1553 & n1637 ) ;
  assign n1639 = ( ~n399 & n1590 ) | ( ~n399 & n1638 ) | ( n1590 & n1638 ) ;
  assign n1640 = ( ~n345 & n1566 ) | ( ~n345 & n1639 ) | ( n1566 & n1639 ) ;
  assign n1641 = ( ~n302 & n1587 ) | ( ~n302 & n1640 ) | ( n1587 & n1640 ) ;
  assign n1642 = ( ~n261 & n1543 ) | ( ~n261 & n1641 ) | ( n1543 & n1641 ) ;
  assign n1643 = ( ~n217 & n1607 ) | ( ~n217 & n1642 ) | ( n1607 & n1642 ) ;
  assign n1644 = ( ~n179 & n1548 ) | ( ~n179 & n1643 ) | ( n1548 & n1643 ) ;
  assign n1645 = ( ~n144 & n1588 ) | ( ~n144 & n1644 ) | ( n1588 & n1644 ) ;
  assign n1646 = ( ~n134 & n1583 ) | ( ~n134 & n1645 ) | ( n1583 & n1645 ) ;
  assign n1647 = n1558 & n1646 ;
  assign n1648 = ( ~x30 & n1611 ) | ( ~x30 & n1646 ) | ( n1611 & n1646 ) ;
  assign n1649 = ~n136 & n1648 ;
  assign n1650 = n1647 | n1649 ;
  assign n1651 = n1615 | n1650 ;
  assign n1652 = n1616 | n1651 ;
  assign n1653 = n1645 ^ n134 ^ 1'b0 ;
  assign n1654 = n1652 & n1653 ;
  assign n1655 = n1654 ^ n1652 ^ n1583 ;
  assign n1656 = n1627 ^ n1220 ^ 1'b0 ;
  assign n1657 = n1652 & n1656 ;
  assign n1658 = n1657 ^ n1652 ^ n1559 ;
  assign n1659 = n1629 ^ n1034 ^ 1'b0 ;
  assign n1660 = n1652 & n1659 ;
  assign n1661 = n1660 ^ n1652 ^ n1571 ;
  assign n1662 = n1633 ^ n716 ^ 1'b0 ;
  assign n1663 = n1652 & n1662 ;
  assign n1664 = n1663 ^ n1652 ^ n1617 ;
  assign n1665 = n1635 ^ n572 ^ 1'b0 ;
  assign n1666 = n1652 & n1665 ;
  assign n1667 = n1666 ^ n1652 ^ n1544 ;
  assign n1668 = n1637 ^ n458 ^ 1'b0 ;
  assign n1669 = n1652 & n1668 ;
  assign n1670 = n1669 ^ n1652 ^ n1553 ;
  assign n1671 = n1639 ^ n345 ^ 1'b0 ;
  assign n1672 = n1652 & n1671 ;
  assign n1673 = n1672 ^ n1652 ^ n1566 ;
  assign n1674 = n1641 ^ n261 ^ 1'b0 ;
  assign n1675 = n1652 & n1674 ;
  assign n1676 = n1675 ^ n1652 ^ n1543 ;
  assign n1677 = ~n1619 & n1652 ;
  assign n1678 = ( n1615 & n1616 ) | ( n1615 & ~n1677 ) | ( n1616 & ~n1677 ) ;
  assign n1679 = n1534 & ~n1650 ;
  assign n1680 = n1677 | n1679 ;
  assign n1681 = ( n1677 & ~n1678 ) | ( n1677 & n1680 ) | ( ~n1678 & n1680 ) ;
  assign n1682 = ( x106 & n1531 ) | ( x106 & n1652 ) | ( n1531 & n1652 ) ;
  assign n1683 = ( ~n1531 & n1613 ) | ( ~n1531 & n1682 ) | ( n1613 & n1682 ) ;
  assign n1684 = ~n1682 & n1683 ;
  assign n1685 = ( n1584 & ~n1622 ) | ( n1584 & n1652 ) | ( ~n1622 & n1652 ) ;
  assign n1686 = ~n1584 & n1685 ;
  assign n1687 = n1686 ^ n1623 ^ x109 ;
  assign n1688 = n1652 ^ n1626 ^ n1318 ;
  assign n1689 = n1652 & n1688 ;
  assign n1690 = n1689 ^ n1606 ^ x110 ;
  assign n1691 = n1652 ^ n1628 ^ n1118 ;
  assign n1692 = n1652 & n1691 ;
  assign n1693 = n1692 ^ n1598 ^ n1496 ;
  assign n1694 = n1652 ^ n1630 ^ n941 ;
  assign n1695 = n1652 & n1694 ;
  assign n1696 = n1695 ^ n1610 ^ n1455 ;
  assign n1697 = n1652 ^ n1631 ^ n859 ;
  assign n1698 = n1652 & n1697 ;
  assign n1699 = n1698 ^ n1550 ^ n1476 ;
  assign n1700 = n1652 ^ n1632 ^ n785 ;
  assign n1701 = n1652 & n1700 ;
  assign n1702 = n1701 ^ n1555 ^ n1459 ;
  assign n1703 = n1652 ^ n1634 ^ n640 ;
  assign n1704 = n1652 & n1703 ;
  assign n1705 = n1704 ^ n1542 ^ n1462 ;
  assign n1706 = n1652 ^ n1636 ^ n514 ;
  assign n1707 = n1652 & n1706 ;
  assign n1708 = n1707 ^ n1591 ^ n1446 ;
  assign n1709 = n1652 ^ n1638 ^ n399 ;
  assign n1710 = n1652 & n1709 ;
  assign n1711 = n1710 ^ n1589 ^ n1478 ;
  assign n1712 = n1652 ^ n1640 ^ n302 ;
  assign n1713 = n1652 & n1712 ;
  assign n1714 = n1713 ^ n1568 ^ n1477 ;
  assign n1715 = n1652 ^ n1642 ^ n217 ;
  assign n1716 = n1652 & n1715 ;
  assign n1717 = n1716 ^ n1573 ^ n1419 ;
  assign n1718 = n1652 ^ n1643 ^ n179 ;
  assign n1719 = n1652 & n1718 ;
  assign n1720 = n1719 ^ n1545 ^ n1427 ;
  assign n1721 = n1652 ^ n1644 ^ n144 ;
  assign n1722 = n1652 & n1721 ;
  assign n1723 = n1722 ^ n1575 ^ n1430 ;
  assign n1724 = ( n136 & n1558 ) | ( n136 & n1646 ) | ( n1558 & n1646 ) ;
  assign n1725 = ( n1646 & n1647 ) | ( n1646 & ~n1652 ) | ( n1647 & ~n1652 ) ;
  assign n1726 = n1724 & ~n1725 ;
  assign n1727 = ~x106 & n1652 ;
  assign n1728 = x103 | x104 ;
  assign n1729 = n1727 ^ x107 ^ 1'b0 ;
  assign n1730 = ( x106 & n1534 ) | ( x106 & ~n1728 ) | ( n1534 & ~n1728 ) ;
  assign n1731 = ( ~x106 & n1534 ) | ( ~x106 & n1652 ) | ( n1534 & n1652 ) ;
  assign n1732 = n1730 & n1731 ;
  assign n1733 = n1681 ^ x108 ^ 1'b0 ;
  assign n1734 = n1558 & ~n1646 ;
  assign n1735 = n1684 | n1729 ;
  assign n1736 = ( n1558 & ~n1646 ) | ( n1558 & n1652 ) | ( ~n1646 & n1652 ) ;
  assign n1737 = ( n1655 & ~n1734 ) | ( n1655 & n1736 ) | ( ~n1734 & n1736 ) ;
  assign n1738 = ~n1732 & n1735 ;
  assign n1739 = ( ~n1416 & n1733 ) | ( ~n1416 & n1738 ) | ( n1733 & n1738 ) ;
  assign n1740 = ( ~n1318 & n1687 ) | ( ~n1318 & n1739 ) | ( n1687 & n1739 ) ;
  assign n1741 = ( ~n1220 & n1690 ) | ( ~n1220 & n1740 ) | ( n1690 & n1740 ) ;
  assign n1742 = ( ~n1118 & n1658 ) | ( ~n1118 & n1741 ) | ( n1658 & n1741 ) ;
  assign n1743 = ( ~n1034 & n1693 ) | ( ~n1034 & n1742 ) | ( n1693 & n1742 ) ;
  assign n1744 = ( ~n941 & n1661 ) | ( ~n941 & n1743 ) | ( n1661 & n1743 ) ;
  assign n1745 = ( ~n859 & n1696 ) | ( ~n859 & n1744 ) | ( n1696 & n1744 ) ;
  assign n1746 = ( ~n785 & n1699 ) | ( ~n785 & n1745 ) | ( n1699 & n1745 ) ;
  assign n1747 = ( ~n716 & n1702 ) | ( ~n716 & n1746 ) | ( n1702 & n1746 ) ;
  assign n1748 = ( ~n640 & n1664 ) | ( ~n640 & n1747 ) | ( n1664 & n1747 ) ;
  assign n1749 = ( ~n572 & n1705 ) | ( ~n572 & n1748 ) | ( n1705 & n1748 ) ;
  assign n1750 = ( ~n514 & n1667 ) | ( ~n514 & n1749 ) | ( n1667 & n1749 ) ;
  assign n1751 = ( ~n458 & n1708 ) | ( ~n458 & n1750 ) | ( n1708 & n1750 ) ;
  assign n1752 = ( ~n399 & n1670 ) | ( ~n399 & n1751 ) | ( n1670 & n1751 ) ;
  assign n1753 = ( ~n345 & n1711 ) | ( ~n345 & n1752 ) | ( n1711 & n1752 ) ;
  assign n1754 = ( ~n302 & n1673 ) | ( ~n302 & n1753 ) | ( n1673 & n1753 ) ;
  assign n1755 = ( ~n261 & n1714 ) | ( ~n261 & n1754 ) | ( n1714 & n1754 ) ;
  assign n1756 = ( ~n217 & n1676 ) | ( ~n217 & n1755 ) | ( n1676 & n1755 ) ;
  assign n1757 = ( ~n179 & n1717 ) | ( ~n179 & n1756 ) | ( n1717 & n1756 ) ;
  assign n1758 = ( ~n144 & n1720 ) | ( ~n144 & n1757 ) | ( n1720 & n1757 ) ;
  assign n1759 = ( ~n134 & n1723 ) | ( ~n134 & n1758 ) | ( n1723 & n1758 ) ;
  assign n1760 = n1655 & n1759 ;
  assign n1761 = ( n1558 & ~n1652 ) | ( n1558 & n1760 ) | ( ~n1652 & n1760 ) ;
  assign n1762 = ( ~x30 & n1737 ) | ( ~x30 & n1759 ) | ( n1737 & n1759 ) ;
  assign n1763 = ~n136 & n1762 ;
  assign n1764 = n1760 | n1763 ;
  assign n1765 = ( n1726 & ~n1761 ) | ( n1726 & n1764 ) | ( ~n1761 & n1764 ) ;
  assign n1766 = n1761 | n1765 ;
  assign n1767 = n1766 ^ n1756 ^ n179 ;
  assign n1768 = n1766 ^ n1750 ^ n458 ;
  assign n1769 = n1766 & n1767 ;
  assign n1770 = n1766 & n1768 ;
  assign n1771 = n1769 ^ n1716 ^ n1607 ;
  assign n1772 = n1770 ^ n1707 ^ n1592 ;
  assign n1773 = ( n1684 & ~n1732 ) | ( n1684 & n1766 ) | ( ~n1732 & n1766 ) ;
  assign n1774 = ~n1684 & n1773 ;
  assign n1775 = n1766 ^ n1742 ^ n1034 ;
  assign n1776 = n1766 ^ n1754 ^ n261 ;
  assign n1777 = n1766 & n1776 ;
  assign n1778 = n1766 & n1775 ;
  assign n1779 = n1778 ^ n1692 ^ n1599 ;
  assign n1780 = n1766 ^ n1748 ^ n572 ;
  assign n1781 = n1766 & n1780 ;
  assign n1782 = n1781 ^ n1704 ^ n1547 ;
  assign n1783 = n1766 ^ n1758 ^ n134 ;
  assign n1784 = n1766 & n1783 ;
  assign n1785 = n1784 ^ n1722 ^ n1588 ;
  assign n1786 = n1766 ^ n1739 ^ n1318 ;
  assign n1787 = n1766 & n1786 ;
  assign n1788 = n1787 ^ n1686 ^ n1624 ;
  assign n1789 = n1777 ^ n1713 ^ n1587 ;
  assign n1790 = n1766 ^ n1744 ^ n859 ;
  assign n1791 = n1766 ^ n1740 ^ n1220 ;
  assign n1792 = n1743 ^ n941 ^ 1'b0 ;
  assign n1793 = n1766 & n1792 ;
  assign n1794 = ~n1728 & n1766 ;
  assign n1795 = n1741 ^ n1118 ^ 1'b0 ;
  assign n1796 = n1766 & n1791 ;
  assign n1797 = n1747 ^ n640 ^ 1'b0 ;
  assign n1798 = n1796 ^ n1689 ^ n1618 ;
  assign n1799 = ( n1652 & ~n1764 ) | ( n1652 & n1794 ) | ( ~n1764 & n1794 ) ;
  assign n1800 = n1726 & ~n1794 ;
  assign n1801 = ( n1794 & n1799 ) | ( n1794 & ~n1800 ) | ( n1799 & ~n1800 ) ;
  assign n1802 = n1749 ^ n514 ^ 1'b0 ;
  assign n1803 = n1416 & n1738 ;
  assign n1804 = ( ~n1416 & n1766 ) | ( ~n1416 & n1803 ) | ( n1766 & n1803 ) ;
  assign n1805 = n1766 & n1802 ;
  assign n1806 = n1766 & n1797 ;
  assign n1807 = n1766 & n1795 ;
  assign n1808 = n1751 ^ n399 ^ 1'b0 ;
  assign n1809 = n1774 ^ n1727 ^ x107 ;
  assign n1810 = n1755 ^ n217 ^ 1'b0 ;
  assign n1811 = n1766 ^ n1757 ^ n144 ;
  assign n1812 = n1766 ^ n1746 ^ n716 ;
  assign n1813 = n1766 ^ n1752 ^ n345 ;
  assign n1814 = n1766 & n1808 ;
  assign n1815 = ( ~n1738 & n1803 ) | ( ~n1738 & n1804 ) | ( n1803 & n1804 ) ;
  assign n1816 = n1766 & n1790 ;
  assign n1817 = n1753 ^ n302 ^ 1'b0 ;
  assign n1818 = n1766 & n1817 ;
  assign n1819 = n1766 ^ n1745 ^ n785 ;
  assign n1820 = ( n136 & n1655 ) | ( n136 & n1759 ) | ( n1655 & n1759 ) ;
  assign n1821 = n1766 & n1819 ;
  assign n1822 = n1815 ^ n1681 ^ x108 ;
  assign n1823 = n1816 ^ n1695 ^ n1612 ;
  assign n1824 = n1821 ^ n1698 ^ n1552 ;
  assign n1825 = n1766 & n1812 ;
  assign n1826 = n1825 ^ n1701 ^ n1556 ;
  assign n1827 = ( n1759 & n1760 ) | ( n1759 & ~n1766 ) | ( n1760 & ~n1766 ) ;
  assign n1828 = n1766 & n1813 ;
  assign n1829 = n1766 & n1811 ;
  assign n1830 = n1828 ^ n1710 ^ n1590 ;
  assign n1831 = n1829 ^ n1719 ^ n1548 ;
  assign n1832 = n1766 & n1810 ;
  assign n1833 = n1793 ^ n1766 ^ n1661 ;
  assign n1834 = n1806 ^ n1766 ^ n1664 ;
  assign n1835 = n1805 ^ n1766 ^ n1667 ;
  assign n1836 = n1814 ^ n1766 ^ n1670 ;
  assign n1837 = n1818 ^ n1766 ^ n1673 ;
  assign n1838 = n1832 ^ n1766 ^ n1676 ;
  assign n1839 = n1807 ^ n1766 ^ n1658 ;
  assign n1840 = n1820 & ~n1827 ;
  assign n1841 = x103 & n1766 ;
  assign n1842 = x101 | x102 ;
  assign n1843 = n1841 ^ n1766 ^ x104 ;
  assign n1844 = ( x103 & ~n1650 ) | ( x103 & n1842 ) | ( ~n1650 & n1842 ) ;
  assign n1845 = ( ~n1652 & n1841 ) | ( ~n1652 & n1844 ) | ( n1841 & n1844 ) ;
  assign n1846 = ~n1841 & n1845 ;
  assign n1847 = n1843 | n1846 ;
  assign n1848 = ( n1655 & ~n1759 ) | ( n1655 & n1766 ) | ( ~n1759 & n1766 ) ;
  assign n1849 = n1655 & ~n1759 ;
  assign n1850 = ( n1785 & n1848 ) | ( n1785 & ~n1849 ) | ( n1848 & ~n1849 ) ;
  assign n1851 = n1801 ^ x106 ^ 1'b0 ;
  assign n1852 = ( ~x103 & n1652 ) | ( ~x103 & n1766 ) | ( n1652 & n1766 ) ;
  assign n1853 = ( x103 & n1652 ) | ( x103 & ~n1842 ) | ( n1652 & ~n1842 ) ;
  assign n1854 = n1852 & n1853 ;
  assign n1855 = n1847 & ~n1854 ;
  assign n1856 = ( ~n1534 & n1851 ) | ( ~n1534 & n1855 ) | ( n1851 & n1855 ) ;
  assign n1857 = ( ~n1416 & n1809 ) | ( ~n1416 & n1856 ) | ( n1809 & n1856 ) ;
  assign n1858 = ( ~n1318 & n1822 ) | ( ~n1318 & n1857 ) | ( n1822 & n1857 ) ;
  assign n1859 = ( ~n1220 & n1788 ) | ( ~n1220 & n1858 ) | ( n1788 & n1858 ) ;
  assign n1860 = ( ~n1118 & n1798 ) | ( ~n1118 & n1859 ) | ( n1798 & n1859 ) ;
  assign n1861 = ( ~n1034 & n1839 ) | ( ~n1034 & n1860 ) | ( n1839 & n1860 ) ;
  assign n1862 = ( ~n941 & n1779 ) | ( ~n941 & n1861 ) | ( n1779 & n1861 ) ;
  assign n1863 = ( ~n859 & n1833 ) | ( ~n859 & n1862 ) | ( n1833 & n1862 ) ;
  assign n1864 = ( ~n785 & n1823 ) | ( ~n785 & n1863 ) | ( n1823 & n1863 ) ;
  assign n1865 = ( ~n716 & n1824 ) | ( ~n716 & n1864 ) | ( n1824 & n1864 ) ;
  assign n1866 = ( ~n640 & n1826 ) | ( ~n640 & n1865 ) | ( n1826 & n1865 ) ;
  assign n1867 = ( ~n572 & n1834 ) | ( ~n572 & n1866 ) | ( n1834 & n1866 ) ;
  assign n1868 = ( ~n514 & n1782 ) | ( ~n514 & n1867 ) | ( n1782 & n1867 ) ;
  assign n1869 = ( ~n458 & n1835 ) | ( ~n458 & n1868 ) | ( n1835 & n1868 ) ;
  assign n1870 = ( ~n399 & n1772 ) | ( ~n399 & n1869 ) | ( n1772 & n1869 ) ;
  assign n1871 = ( ~n345 & n1836 ) | ( ~n345 & n1870 ) | ( n1836 & n1870 ) ;
  assign n1872 = ( ~n302 & n1830 ) | ( ~n302 & n1871 ) | ( n1830 & n1871 ) ;
  assign n1873 = ( ~n261 & n1837 ) | ( ~n261 & n1872 ) | ( n1837 & n1872 ) ;
  assign n1874 = ( ~n217 & n1789 ) | ( ~n217 & n1873 ) | ( n1789 & n1873 ) ;
  assign n1875 = ( ~n179 & n1838 ) | ( ~n179 & n1874 ) | ( n1838 & n1874 ) ;
  assign n1876 = n1655 & ~n1766 ;
  assign n1877 = ( ~n144 & n1771 ) | ( ~n144 & n1875 ) | ( n1771 & n1875 ) ;
  assign n1878 = ( ~n134 & n1831 ) | ( ~n134 & n1877 ) | ( n1831 & n1877 ) ;
  assign n1879 = ( ~x30 & n1850 ) | ( ~x30 & n1878 ) | ( n1850 & n1878 ) ;
  assign n1880 = ~n136 & n1879 ;
  assign n1881 = n1846 | n1854 ;
  assign n1882 = n1785 & n1878 ;
  assign n1883 = n1876 | n1882 ;
  assign n1884 = n1880 | n1883 ;
  assign n1885 = n1840 | n1884 ;
  assign n1886 = n1885 ^ n1875 ^ n144 ;
  assign n1887 = n1885 ^ n1858 ^ n1220 ;
  assign n1888 = n1885 & n1887 ;
  assign n1889 = n1885 ^ n1869 ^ n399 ;
  assign n1890 = n1885 & n1889 ;
  assign n1891 = n1881 & n1885 ;
  assign n1892 = n1891 ^ n1885 ^ n1843 ;
  assign n1893 = n1888 ^ n1787 ^ n1687 ;
  assign n1894 = n1885 ^ n1857 ^ n1318 ;
  assign n1895 = n1885 ^ n1859 ^ n1118 ;
  assign n1896 = n1885 & n1894 ;
  assign n1897 = n1896 ^ n1815 ^ n1733 ;
  assign n1898 = n1885 & n1895 ;
  assign n1899 = n1898 ^ n1796 ^ n1690 ;
  assign n1900 = n1885 & n1886 ;
  assign n1901 = n1885 ^ n1856 ^ n1416 ;
  assign n1902 = n1885 ^ n1877 ^ n134 ;
  assign n1903 = n1900 ^ n1769 ^ n1717 ;
  assign n1904 = n1885 & n1901 ;
  assign n1905 = n1885 ^ n1863 ^ n785 ;
  assign n1906 = n1890 ^ n1770 ^ n1708 ;
  assign n1907 = n1885 & n1905 ;
  assign n1908 = n1907 ^ n1816 ^ n1696 ;
  assign n1909 = n1885 & n1902 ;
  assign n1910 = n1909 ^ n1829 ^ n1720 ;
  assign n1911 = n1904 ^ n1774 ^ n1729 ;
  assign n1912 = n1885 ^ n1865 ^ n640 ;
  assign n1913 = n1885 & n1912 ;
  assign n1914 = n1913 ^ n1825 ^ n1702 ;
  assign n1915 = ( n1766 & n1876 ) | ( n1766 & ~n1885 ) | ( n1876 & ~n1885 ) ;
  assign n1916 = n1860 ^ n1034 ^ 1'b0 ;
  assign n1917 = n1885 & n1916 ;
  assign n1918 = n1885 ^ n1867 ^ n514 ;
  assign n1919 = n1885 & n1918 ;
  assign n1920 = n1917 ^ n1885 ^ n1839 ;
  assign n1921 = n1885 ^ n1873 ^ n217 ;
  assign n1922 = n1870 ^ n345 ^ 1'b0 ;
  assign n1923 = n1885 ^ n1861 ^ n941 ;
  assign n1924 = n1885 & n1923 ;
  assign n1925 = ( n1878 & n1882 ) | ( n1878 & ~n1885 ) | ( n1882 & ~n1885 ) ;
  assign n1926 = n1885 ^ n1871 ^ n302 ;
  assign n1927 = ( x97 & x98 ) | ( x97 & ~n1876 ) | ( x98 & ~n1876 ) ;
  assign n1928 = n1885 ^ n1864 ^ n716 ;
  assign n1929 = n1885 & n1928 ;
  assign n1930 = ( x99 & ~n1876 ) | ( x99 & n1927 ) | ( ~n1876 & n1927 ) ;
  assign n1931 = n1924 ^ n1778 ^ n1693 ;
  assign n1932 = ( n136 & n1785 ) | ( n136 & n1878 ) | ( n1785 & n1878 ) ;
  assign n1933 = ( ~n1840 & n1883 ) | ( ~n1840 & n1930 ) | ( n1883 & n1930 ) ;
  assign n1934 = n1868 ^ n458 ^ 1'b0 ;
  assign n1935 = n1929 ^ n1821 ^ n1699 ;
  assign n1936 = n1862 ^ n859 ^ 1'b0 ;
  assign n1937 = n1885 & n1934 ;
  assign n1938 = n1937 ^ n1885 ^ n1835 ;
  assign n1939 = ~n1785 & n1878 ;
  assign n1940 = ( ~n1785 & n1878 ) | ( ~n1785 & n1885 ) | ( n1878 & n1885 ) ;
  assign n1941 = ( n1785 & ~n1840 ) | ( n1785 & n1876 ) | ( ~n1840 & n1876 ) ;
  assign n1942 = n1885 & n1922 ;
  assign n1943 = n1866 ^ n572 ^ 1'b0 ;
  assign n1944 = n1942 ^ n1885 ^ n1836 ;
  assign n1945 = n1874 ^ n179 ^ 1'b0 ;
  assign n1946 = n1885 & n1945 ;
  assign n1947 = ~n1925 & n1932 ;
  assign n1948 = n1885 & n1936 ;
  assign n1949 = n1885 ^ n1855 ^ n1534 ;
  assign n1950 = n1842 & n1885 ;
  assign n1951 = n1885 & n1949 ;
  assign n1952 = n1872 ^ n261 ^ 1'b0 ;
  assign n1953 = n1948 ^ n1885 ^ n1833 ;
  assign n1954 = n1885 & n1952 ;
  assign n1955 = ( n1885 & n1915 ) | ( n1885 & ~n1950 ) | ( n1915 & ~n1950 ) ;
  assign n1956 = n1951 ^ n1801 ^ x106 ;
  assign n1957 = n1885 & n1921 ;
  assign n1958 = n1885 & n1943 ;
  assign n1959 = n1885 & n1926 ;
  assign n1960 = n1954 ^ n1885 ^ n1837 ;
  assign n1961 = n1958 ^ n1885 ^ n1834 ;
  assign n1962 = n1959 ^ n1828 ^ n1711 ;
  assign n1963 = n1919 ^ n1781 ^ n1705 ;
  assign n1964 = n1946 ^ n1885 ^ n1838 ;
  assign n1965 = ( n1910 & ~n1939 ) | ( n1910 & n1940 ) | ( ~n1939 & n1940 ) ;
  assign n1966 = ~n1884 & n1941 ;
  assign n1967 = ~n1883 & n1933 ;
  assign n1968 = n1957 ^ n1777 ^ n1714 ;
  assign n1969 = x99 | x100 ;
  assign n1970 = ( x101 & ~n1764 ) | ( x101 & n1969 ) | ( ~n1764 & n1969 ) ;
  assign n1971 = x101 & n1885 ;
  assign n1972 = ( ~n1766 & n1970 ) | ( ~n1766 & n1971 ) | ( n1970 & n1971 ) ;
  assign n1973 = x101 | n1969 ;
  assign n1974 = ( n1766 & n1971 ) | ( n1766 & ~n1973 ) | ( n1971 & ~n1973 ) ;
  assign n1975 = ~n1971 & n1972 ;
  assign n1976 = n1971 ^ n1885 ^ x102 ;
  assign n1977 = n1975 | n1976 ;
  assign n1978 = ~n1974 & n1977 ;
  assign n1979 = n1955 ^ x103 ^ 1'b0 ;
  assign n1980 = ( ~n1652 & n1978 ) | ( ~n1652 & n1979 ) | ( n1978 & n1979 ) ;
  assign n1981 = ( ~n1534 & n1892 ) | ( ~n1534 & n1980 ) | ( n1892 & n1980 ) ;
  assign n1982 = ( ~n1416 & n1956 ) | ( ~n1416 & n1981 ) | ( n1956 & n1981 ) ;
  assign n1983 = ( ~n1318 & n1911 ) | ( ~n1318 & n1982 ) | ( n1911 & n1982 ) ;
  assign n1984 = ( ~n1220 & n1897 ) | ( ~n1220 & n1983 ) | ( n1897 & n1983 ) ;
  assign n1985 = ( ~n1118 & n1893 ) | ( ~n1118 & n1984 ) | ( n1893 & n1984 ) ;
  assign n1986 = ( ~n1034 & n1899 ) | ( ~n1034 & n1985 ) | ( n1899 & n1985 ) ;
  assign n1987 = ( ~n941 & n1920 ) | ( ~n941 & n1986 ) | ( n1920 & n1986 ) ;
  assign n1988 = ( ~n859 & n1931 ) | ( ~n859 & n1987 ) | ( n1931 & n1987 ) ;
  assign n1989 = ( ~n785 & n1953 ) | ( ~n785 & n1988 ) | ( n1953 & n1988 ) ;
  assign n1990 = ( ~n716 & n1908 ) | ( ~n716 & n1989 ) | ( n1908 & n1989 ) ;
  assign n1991 = ( ~n640 & n1935 ) | ( ~n640 & n1990 ) | ( n1935 & n1990 ) ;
  assign n1992 = ( ~n572 & n1914 ) | ( ~n572 & n1991 ) | ( n1914 & n1991 ) ;
  assign n1993 = ( ~n514 & n1961 ) | ( ~n514 & n1992 ) | ( n1961 & n1992 ) ;
  assign n1994 = ( ~n458 & n1963 ) | ( ~n458 & n1993 ) | ( n1963 & n1993 ) ;
  assign n1995 = ( ~n399 & n1938 ) | ( ~n399 & n1994 ) | ( n1938 & n1994 ) ;
  assign n1996 = ( ~n345 & n1906 ) | ( ~n345 & n1995 ) | ( n1906 & n1995 ) ;
  assign n1997 = ( ~n302 & n1944 ) | ( ~n302 & n1996 ) | ( n1944 & n1996 ) ;
  assign n1998 = ( ~n261 & n1962 ) | ( ~n261 & n1997 ) | ( n1962 & n1997 ) ;
  assign n1999 = ( ~n217 & n1960 ) | ( ~n217 & n1998 ) | ( n1960 & n1998 ) ;
  assign n2000 = ( ~n179 & n1968 ) | ( ~n179 & n1999 ) | ( n1968 & n1999 ) ;
  assign n2001 = ( ~n144 & n1964 ) | ( ~n144 & n2000 ) | ( n1964 & n2000 ) ;
  assign n2002 = ( ~n134 & n1903 ) | ( ~n134 & n2001 ) | ( n1903 & n2001 ) ;
  assign n2003 = n1910 & n2002 ;
  assign n2004 = ( ~x30 & n1965 ) | ( ~x30 & n2002 ) | ( n1965 & n2002 ) ;
  assign n2005 = ~n136 & n2004 ;
  assign n2006 = n1966 | n2003 ;
  assign n2007 = n2005 | n2006 ;
  assign n2008 = n1974 | n1975 ;
  assign n2009 = n1947 | n2007 ;
  assign n2010 = n2009 ^ n1984 ^ n1118 ;
  assign n2011 = n2009 & n2010 ;
  assign n2012 = n2009 ^ n1997 ^ n261 ;
  assign n2013 = n2009 & n2012 ;
  assign n2014 = n2013 ^ n1959 ^ n1830 ;
  assign n2015 = n2009 ^ n1995 ^ n345 ;
  assign n2016 = n2011 ^ n1888 ^ n1788 ;
  assign n2017 = n2009 ^ n2001 ^ n134 ;
  assign n2018 = n2009 ^ n1983 ^ n1220 ;
  assign n2019 = n2009 & n2018 ;
  assign n2020 = n2019 ^ n1896 ^ n1822 ;
  assign n2021 = n2009 ^ n1990 ^ n640 ;
  assign n2022 = n2009 & n2015 ;
  assign n2023 = n2022 ^ n1890 ^ n1772 ;
  assign n2024 = n2009 & n2017 ;
  assign n2025 = n2009 & n2021 ;
  assign n2026 = n2025 ^ n1929 ^ n1824 ;
  assign n2027 = n2009 ^ n1982 ^ n1318 ;
  assign n2028 = n2024 ^ n1900 ^ n1771 ;
  assign n2029 = n2009 & n2027 ;
  assign n2030 = n2029 ^ n1904 ^ n1809 ;
  assign n2031 = n2009 ^ n1993 ^ n458 ;
  assign n2032 = n2008 & n2009 ;
  assign n2033 = n2032 ^ n2009 ^ n1976 ;
  assign n2034 = n2009 & n2031 ;
  assign n2035 = ( x99 & n1880 ) | ( x99 & n2009 ) | ( n1880 & n2009 ) ;
  assign n2036 = ( ~n1880 & n1967 ) | ( ~n1880 & n2035 ) | ( n1967 & n2035 ) ;
  assign n2037 = ~n2035 & n2036 ;
  assign n2038 = n2034 ^ n1919 ^ n1782 ;
  assign n2039 = n1994 ^ n399 ^ 1'b0 ;
  assign n2040 = n1998 ^ n217 ^ 1'b0 ;
  assign n2041 = n1988 ^ n785 ^ 1'b0 ;
  assign n2042 = n2000 ^ n144 ^ 1'b0 ;
  assign n2043 = n2009 ^ n1981 ^ n1416 ;
  assign n2044 = n2009 & n2043 ;
  assign n2045 = n2044 ^ n1951 ^ n1851 ;
  assign n2046 = n2009 & n2041 ;
  assign n2047 = n1947 | n2003 ;
  assign n2048 = n2009 & n2039 ;
  assign n2049 = n1992 ^ n514 ^ 1'b0 ;
  assign n2050 = n2009 & n2049 ;
  assign n2051 = n2009 ^ n1987 ^ n859 ;
  assign n2052 = n2050 ^ n2009 ^ n1961 ;
  assign n2053 = ( x95 & x96 ) | ( x95 & ~n1947 ) | ( x96 & ~n1947 ) ;
  assign n2054 = n2009 ^ n1985 ^ n1034 ;
  assign n2055 = ( x97 & ~n1947 ) | ( x97 & n2053 ) | ( ~n1947 & n2053 ) ;
  assign n2056 = ( ~n1966 & n2047 ) | ( ~n1966 & n2055 ) | ( n2047 & n2055 ) ;
  assign n2057 = ~n2047 & n2056 ;
  assign n2058 = ( n1910 & ~n1947 ) | ( n1910 & n1966 ) | ( ~n1947 & n1966 ) ;
  assign n2059 = n1996 ^ n302 ^ 1'b0 ;
  assign n2060 = ( n2002 & n2003 ) | ( n2002 & ~n2009 ) | ( n2003 & ~n2009 ) ;
  assign n2061 = n2009 & n2059 ;
  assign n2062 = n2061 ^ n2009 ^ n1944 ;
  assign n2063 = ~n1910 & n2002 ;
  assign n2064 = ~n2007 & n2058 ;
  assign n2065 = n2009 & n2051 ;
  assign n2066 = ( n1885 & ~n1947 ) | ( n1885 & n1966 ) | ( ~n1947 & n1966 ) ;
  assign n2067 = n2009 & n2042 ;
  assign n2068 = n1986 ^ n941 ^ 1'b0 ;
  assign n2069 = n2009 ^ n1999 ^ n179 ;
  assign n2070 = n2046 ^ n2009 ^ n1953 ;
  assign n2071 = n2009 & n2069 ;
  assign n2072 = n1980 ^ n1534 ^ 1'b0 ;
  assign n2073 = n2009 & n2072 ;
  assign n2074 = n2009 & n2054 ;
  assign n2075 = n2009 & n2068 ;
  assign n2076 = n2075 ^ n2009 ^ n1920 ;
  assign n2077 = n2009 ^ n1989 ^ n716 ;
  assign n2078 = n2009 ^ n1978 ^ n1652 ;
  assign n2079 = ( n136 & n1910 ) | ( n136 & n2002 ) | ( n1910 & n2002 ) ;
  assign n2080 = n2009 ^ n1991 ^ n572 ;
  assign n2081 = n2009 & n2080 ;
  assign n2082 = n2009 & n2077 ;
  assign n2083 = ( ~n1910 & n2002 ) | ( ~n1910 & n2009 ) | ( n2002 & n2009 ) ;
  assign n2084 = ~n2060 & n2079 ;
  assign n2085 = n2009 & n2040 ;
  assign n2086 = n2074 ^ n1898 ^ n1798 ;
  assign n2087 = ~n1969 & n2009 ;
  assign n2088 = n2007 & ~n2087 ;
  assign n2089 = n2085 ^ n2009 ^ n1960 ;
  assign n2090 = n2073 ^ n2009 ^ n1892 ;
  assign n2091 = n2081 ^ n1913 ^ n1826 ;
  assign n2092 = ( n2028 & ~n2063 ) | ( n2028 & n2083 ) | ( ~n2063 & n2083 ) ;
  assign n2093 = n2082 ^ n1907 ^ n1823 ;
  assign n2094 = n2067 ^ n2009 ^ n1964 ;
  assign n2095 = n2071 ^ n1957 ^ n1789 ;
  assign n2096 = ( n2066 & n2087 ) | ( n2066 & ~n2088 ) | ( n2087 & ~n2088 ) ;
  assign n2097 = n2048 ^ n2009 ^ n1938 ;
  assign n2098 = n2065 ^ n1924 ^ n1779 ;
  assign n2099 = ( ~x99 & n1885 ) | ( ~x99 & n2009 ) | ( n1885 & n2009 ) ;
  assign n2100 = n2096 ^ x101 ^ 1'b0 ;
  assign n2101 = n2009 & n2078 ;
  assign n2102 = n2101 ^ n1955 ^ x103 ;
  assign n2103 = x97 | x98 ;
  assign n2104 = ( x99 & n1885 ) | ( x99 & ~n2103 ) | ( n1885 & ~n2103 ) ;
  assign n2105 = ~x99 & n2009 ;
  assign n2106 = n2105 ^ x100 ^ 1'b0 ;
  assign n2107 = n2037 | n2106 ;
  assign n2108 = n2099 & n2104 ;
  assign n2109 = n2107 & ~n2108 ;
  assign n2110 = ( ~n1766 & n2100 ) | ( ~n1766 & n2109 ) | ( n2100 & n2109 ) ;
  assign n2111 = ( ~n1652 & n2033 ) | ( ~n1652 & n2110 ) | ( n2033 & n2110 ) ;
  assign n2112 = ( ~n1534 & n2102 ) | ( ~n1534 & n2111 ) | ( n2102 & n2111 ) ;
  assign n2113 = ( ~n1416 & n2090 ) | ( ~n1416 & n2112 ) | ( n2090 & n2112 ) ;
  assign n2114 = ( ~n1318 & n2045 ) | ( ~n1318 & n2113 ) | ( n2045 & n2113 ) ;
  assign n2115 = ( ~n1220 & n2030 ) | ( ~n1220 & n2114 ) | ( n2030 & n2114 ) ;
  assign n2116 = ( ~n1118 & n2020 ) | ( ~n1118 & n2115 ) | ( n2020 & n2115 ) ;
  assign n2117 = ( ~n1034 & n2016 ) | ( ~n1034 & n2116 ) | ( n2016 & n2116 ) ;
  assign n2118 = ( ~n941 & n2086 ) | ( ~n941 & n2117 ) | ( n2086 & n2117 ) ;
  assign n2119 = ( ~n859 & n2076 ) | ( ~n859 & n2118 ) | ( n2076 & n2118 ) ;
  assign n2120 = ( ~n785 & n2098 ) | ( ~n785 & n2119 ) | ( n2098 & n2119 ) ;
  assign n2121 = ( ~n716 & n2070 ) | ( ~n716 & n2120 ) | ( n2070 & n2120 ) ;
  assign n2122 = ( ~n640 & n2093 ) | ( ~n640 & n2121 ) | ( n2093 & n2121 ) ;
  assign n2123 = ( ~n572 & n2026 ) | ( ~n572 & n2122 ) | ( n2026 & n2122 ) ;
  assign n2124 = ( ~n514 & n2091 ) | ( ~n514 & n2123 ) | ( n2091 & n2123 ) ;
  assign n2125 = ( ~n458 & n2052 ) | ( ~n458 & n2124 ) | ( n2052 & n2124 ) ;
  assign n2126 = ( ~n399 & n2038 ) | ( ~n399 & n2125 ) | ( n2038 & n2125 ) ;
  assign n2127 = ( ~n345 & n2097 ) | ( ~n345 & n2126 ) | ( n2097 & n2126 ) ;
  assign n2128 = ( ~n302 & n2023 ) | ( ~n302 & n2127 ) | ( n2023 & n2127 ) ;
  assign n2129 = ( ~n261 & n2062 ) | ( ~n261 & n2128 ) | ( n2062 & n2128 ) ;
  assign n2130 = ( ~n217 & n2014 ) | ( ~n217 & n2129 ) | ( n2014 & n2129 ) ;
  assign n2131 = ( ~n179 & n2089 ) | ( ~n179 & n2130 ) | ( n2089 & n2130 ) ;
  assign n2132 = ( ~n144 & n2095 ) | ( ~n144 & n2131 ) | ( n2095 & n2131 ) ;
  assign n2133 = ( ~n134 & n2094 ) | ( ~n134 & n2132 ) | ( n2094 & n2132 ) ;
  assign n2134 = ( ~x30 & n2092 ) | ( ~x30 & n2133 ) | ( n2092 & n2133 ) ;
  assign n2135 = ~n136 & n2134 ;
  assign n2136 = n2028 & n2133 ;
  assign n2137 = n2135 | n2136 ;
  assign n2138 = n2084 | n2137 ;
  assign n2139 = n2064 | n2138 ;
  assign n2140 = n2139 ^ n2114 ^ n1220 ;
  assign n2141 = ( n2037 & ~n2108 ) | ( n2037 & n2139 ) | ( ~n2108 & n2139 ) ;
  assign n2142 = ~n2037 & n2141 ;
  assign n2143 = ~n2103 & n2139 ;
  assign n2144 = n2139 ^ n2119 ^ n785 ;
  assign n2145 = n2139 & n2144 ;
  assign n2146 = n2139 ^ n2122 ^ n572 ;
  assign n2147 = n2145 ^ n2065 ^ n1931 ;
  assign n2148 = n2139 ^ n2113 ^ n1318 ;
  assign n2149 = ( x97 & n2005 ) | ( x97 & n2139 ) | ( n2005 & n2139 ) ;
  assign n2150 = ( n2064 & n2084 ) | ( n2064 & ~n2143 ) | ( n2084 & ~n2143 ) ;
  assign n2151 = n2139 & n2148 ;
  assign n2152 = n2139 & n2140 ;
  assign n2153 = ( ~n2005 & n2057 ) | ( ~n2005 & n2149 ) | ( n2057 & n2149 ) ;
  assign n2154 = ~n2149 & n2153 ;
  assign n2155 = n2151 ^ n2044 ^ n1956 ;
  assign n2156 = n2152 ^ n2029 ^ n1911 ;
  assign n2157 = n2139 & n2146 ;
  assign n2158 = n2157 ^ n2025 ^ n1935 ;
  assign n2159 = n2139 ^ n2123 ^ n514 ;
  assign n2160 = n2139 & n2159 ;
  assign n2161 = n2160 ^ n2081 ^ n1914 ;
  assign n2162 = n2128 ^ n261 ^ 1'b0 ;
  assign n2163 = n2139 & n2162 ;
  assign n2164 = n2163 ^ n2139 ^ n2062 ;
  assign n2165 = n2139 ^ n2129 ^ n217 ;
  assign n2166 = n2139 & n2165 ;
  assign n2167 = n2166 ^ n2013 ^ n1962 ;
  assign n2168 = n2132 ^ n134 ^ 1'b0 ;
  assign n2169 = n2139 & n2168 ;
  assign n2170 = n2169 ^ n2139 ^ n2094 ;
  assign n2171 = n2009 & ~n2137 ;
  assign n2172 = n2143 | n2171 ;
  assign n2173 = ( n2143 & ~n2150 ) | ( n2143 & n2172 ) | ( ~n2150 & n2172 ) ;
  assign n2174 = n2142 ^ n2105 ^ x100 ;
  assign n2175 = n2139 ^ n2109 ^ n1766 ;
  assign n2176 = n2139 & n2175 ;
  assign n2177 = n2176 ^ n2096 ^ x101 ;
  assign n2178 = n2110 ^ n1652 ^ 1'b0 ;
  assign n2179 = n2139 & n2178 ;
  assign n2180 = n2179 ^ n2139 ^ n2033 ;
  assign n2181 = n2139 ^ n2111 ^ n1534 ;
  assign n2182 = n2139 & n2181 ;
  assign n2183 = n2182 ^ n2101 ^ n1979 ;
  assign n2184 = n2112 ^ n1416 ^ 1'b0 ;
  assign n2185 = n2139 & n2184 ;
  assign n2186 = n2185 ^ n2139 ^ n2090 ;
  assign n2187 = n2139 ^ n2115 ^ n1118 ;
  assign n2188 = n2139 & n2187 ;
  assign n2189 = n2188 ^ n2019 ^ n1897 ;
  assign n2190 = n2139 ^ n2116 ^ n1034 ;
  assign n2191 = n2139 & n2190 ;
  assign n2192 = n2139 ^ n2117 ^ n941 ;
  assign n2193 = n2139 & n2192 ;
  assign n2194 = n2193 ^ n2074 ^ n1899 ;
  assign n2195 = n2118 ^ n859 ^ 1'b0 ;
  assign n2196 = n2139 & n2195 ;
  assign n2197 = n2196 ^ n2139 ^ n2076 ;
  assign n2198 = n2120 ^ n716 ^ 1'b0 ;
  assign n2199 = n2139 & n2198 ;
  assign n2200 = n2199 ^ n2139 ^ n2070 ;
  assign n2201 = n2139 ^ n2121 ^ n640 ;
  assign n2202 = n2139 & n2201 ;
  assign n2203 = n2202 ^ n2082 ^ n1908 ;
  assign n2204 = n2124 ^ n458 ^ 1'b0 ;
  assign n2205 = n2139 & n2204 ;
  assign n2206 = n2205 ^ n2139 ^ n2052 ;
  assign n2207 = n2139 ^ n2125 ^ n399 ;
  assign n2208 = n2139 & n2207 ;
  assign n2209 = n2191 ^ n2011 ^ n1893 ;
  assign n2210 = n2208 ^ n2034 ^ n1963 ;
  assign n2211 = n2126 ^ n345 ^ 1'b0 ;
  assign n2212 = n2139 & n2211 ;
  assign n2213 = n2212 ^ n2139 ^ n2097 ;
  assign n2214 = n2139 ^ n2127 ^ n302 ;
  assign n2215 = n2139 & n2214 ;
  assign n2216 = n2215 ^ n2022 ^ n1906 ;
  assign n2217 = n2130 ^ n179 ^ 1'b0 ;
  assign n2218 = n2139 & n2217 ;
  assign n2219 = n2218 ^ n2139 ^ n2089 ;
  assign n2220 = n2139 ^ n2131 ^ n144 ;
  assign n2221 = n2139 & n2220 ;
  assign n2222 = n2221 ^ n2071 ^ n1968 ;
  assign n2223 = ( n136 & n2028 ) | ( n136 & n2133 ) | ( n2028 & n2133 ) ;
  assign n2224 = ( n2133 & n2136 ) | ( n2133 & ~n2139 ) | ( n2136 & ~n2139 ) ;
  assign n2225 = n2223 & ~n2224 ;
  assign n2226 = ( ~x97 & n2009 ) | ( ~x97 & n2139 ) | ( n2009 & n2139 ) ;
  assign n2227 = ~x97 & n2139 ;
  assign n2228 = n2227 ^ x98 ^ 1'b0 ;
  assign n2229 = n2154 | n2228 ;
  assign n2230 = ( n2028 & ~n2133 ) | ( n2028 & n2139 ) | ( ~n2133 & n2139 ) ;
  assign n2231 = n2173 ^ x99 ^ 1'b0 ;
  assign n2232 = n2028 & ~n2133 ;
  assign n2233 = x95 | x96 ;
  assign n2234 = ( x97 & n2009 ) | ( x97 & ~n2233 ) | ( n2009 & ~n2233 ) ;
  assign n2235 = n2226 & n2234 ;
  assign n2236 = n2229 & ~n2235 ;
  assign n2237 = ( ~n1885 & n2231 ) | ( ~n1885 & n2236 ) | ( n2231 & n2236 ) ;
  assign n2238 = ( ~n1766 & n2174 ) | ( ~n1766 & n2237 ) | ( n2174 & n2237 ) ;
  assign n2239 = ( ~n1652 & n2177 ) | ( ~n1652 & n2238 ) | ( n2177 & n2238 ) ;
  assign n2240 = ( ~n1534 & n2180 ) | ( ~n1534 & n2239 ) | ( n2180 & n2239 ) ;
  assign n2241 = ( ~n1416 & n2183 ) | ( ~n1416 & n2240 ) | ( n2183 & n2240 ) ;
  assign n2242 = ( ~n1318 & n2186 ) | ( ~n1318 & n2241 ) | ( n2186 & n2241 ) ;
  assign n2243 = ( ~n1220 & n2155 ) | ( ~n1220 & n2242 ) | ( n2155 & n2242 ) ;
  assign n2244 = ( ~n1118 & n2156 ) | ( ~n1118 & n2243 ) | ( n2156 & n2243 ) ;
  assign n2245 = ( ~n1034 & n2189 ) | ( ~n1034 & n2244 ) | ( n2189 & n2244 ) ;
  assign n2246 = ( ~n941 & n2209 ) | ( ~n941 & n2245 ) | ( n2209 & n2245 ) ;
  assign n2247 = ( ~n859 & n2194 ) | ( ~n859 & n2246 ) | ( n2194 & n2246 ) ;
  assign n2248 = ( ~n785 & n2197 ) | ( ~n785 & n2247 ) | ( n2197 & n2247 ) ;
  assign n2249 = ( ~n716 & n2147 ) | ( ~n716 & n2248 ) | ( n2147 & n2248 ) ;
  assign n2250 = ( ~n640 & n2200 ) | ( ~n640 & n2249 ) | ( n2200 & n2249 ) ;
  assign n2251 = ( ~n572 & n2203 ) | ( ~n572 & n2250 ) | ( n2203 & n2250 ) ;
  assign n2252 = ( ~n514 & n2158 ) | ( ~n514 & n2251 ) | ( n2158 & n2251 ) ;
  assign n2253 = ( ~n458 & n2161 ) | ( ~n458 & n2252 ) | ( n2161 & n2252 ) ;
  assign n2254 = ( ~n399 & n2206 ) | ( ~n399 & n2253 ) | ( n2206 & n2253 ) ;
  assign n2255 = ( ~n345 & n2210 ) | ( ~n345 & n2254 ) | ( n2210 & n2254 ) ;
  assign n2256 = ( ~n302 & n2213 ) | ( ~n302 & n2255 ) | ( n2213 & n2255 ) ;
  assign n2257 = ( ~n261 & n2216 ) | ( ~n261 & n2256 ) | ( n2216 & n2256 ) ;
  assign n2258 = ( ~n217 & n2164 ) | ( ~n217 & n2257 ) | ( n2164 & n2257 ) ;
  assign n2259 = ( ~n179 & n2167 ) | ( ~n179 & n2258 ) | ( n2167 & n2258 ) ;
  assign n2260 = ( ~n144 & n2219 ) | ( ~n144 & n2259 ) | ( n2219 & n2259 ) ;
  assign n2261 = ( ~n134 & n2222 ) | ( ~n134 & n2260 ) | ( n2222 & n2260 ) ;
  assign n2262 = n2170 & n2261 ;
  assign n2263 = ( n2028 & ~n2139 ) | ( n2028 & n2262 ) | ( ~n2139 & n2262 ) ;
  assign n2264 = ( n2170 & n2230 ) | ( n2170 & ~n2232 ) | ( n2230 & ~n2232 ) ;
  assign n2265 = ( ~x30 & n2261 ) | ( ~x30 & n2264 ) | ( n2261 & n2264 ) ;
  assign n2266 = ~n136 & n2265 ;
  assign n2267 = n2262 | n2266 ;
  assign n2268 = ( n2225 & ~n2263 ) | ( n2225 & n2267 ) | ( ~n2263 & n2267 ) ;
  assign n2269 = n2263 | n2268 ;
  assign n2270 = n2269 ^ n2238 ^ n1652 ;
  assign n2271 = n2269 ^ n2250 ^ n572 ;
  assign n2272 = n2269 & n2271 ;
  assign n2273 = n2272 ^ n2202 ^ n2093 ;
  assign n2274 = n2269 ^ n2244 ^ n1034 ;
  assign n2275 = n2269 & n2274 ;
  assign n2276 = n2275 ^ n2188 ^ n2020 ;
  assign n2277 = n2269 & n2270 ;
  assign n2278 = n2277 ^ n2176 ^ n2100 ;
  assign n2279 = n2269 ^ n2242 ^ n1220 ;
  assign n2280 = n2269 & n2279 ;
  assign n2281 = n2280 ^ n2151 ^ n2045 ;
  assign n2282 = n2269 ^ n2245 ^ n941 ;
  assign n2283 = n2269 & n2282 ;
  assign n2284 = n2283 ^ n2191 ^ n2016 ;
  assign n2285 = n2269 ^ n2248 ^ n716 ;
  assign n2286 = n2269 & n2285 ;
  assign n2287 = n2286 ^ n2145 ^ n2098 ;
  assign n2288 = n2269 ^ n2251 ^ n514 ;
  assign n2289 = n2269 & n2288 ;
  assign n2290 = n2289 ^ n2157 ^ n2026 ;
  assign n2291 = ( n2154 & ~n2235 ) | ( n2154 & n2269 ) | ( ~n2235 & n2269 ) ;
  assign n2292 = ~n2154 & n2291 ;
  assign n2293 = n2269 ^ n2260 ^ n134 ;
  assign n2294 = n2269 & n2293 ;
  assign n2295 = n2294 ^ n2221 ^ n2095 ;
  assign n2296 = ~n2233 & n2269 ;
  assign n2297 = n2269 ^ n2236 ^ n1885 ;
  assign n2298 = n2259 ^ n144 ^ 1'b0 ;
  assign n2299 = n2269 & n2298 ;
  assign n2300 = n2225 & ~n2296 ;
  assign n2301 = n2299 ^ n2269 ^ n2219 ;
  assign n2302 = ( n2139 & ~n2267 ) | ( n2139 & n2296 ) | ( ~n2267 & n2296 ) ;
  assign n2303 = n2249 ^ n640 ^ 1'b0 ;
  assign n2304 = n2247 ^ n785 ^ 1'b0 ;
  assign n2305 = n2269 & n2304 ;
  assign n2306 = n2269 ^ n2246 ^ n859 ;
  assign n2307 = n2269 ^ n2240 ^ n1416 ;
  assign n2308 = n2269 & n2306 ;
  assign n2309 = n2269 ^ n2252 ^ n458 ;
  assign n2310 = n2269 & n2307 ;
  assign n2311 = n2269 & n2309 ;
  assign n2312 = n2269 & n2297 ;
  assign n2313 = n2255 ^ n302 ^ 1'b0 ;
  assign n2314 = n2241 ^ n1318 ^ 1'b0 ;
  assign n2315 = n2269 & n2314 ;
  assign n2316 = n2253 ^ n399 ^ 1'b0 ;
  assign n2317 = n2269 ^ n2258 ^ n179 ;
  assign n2318 = ( n2261 & n2262 ) | ( n2261 & ~n2269 ) | ( n2262 & ~n2269 ) ;
  assign n2319 = n2269 ^ n2237 ^ n1766 ;
  assign n2320 = n2269 & n2303 ;
  assign n2321 = n2269 & n2316 ;
  assign n2322 = n2239 ^ n1534 ^ 1'b0 ;
  assign n2323 = n2269 & n2322 ;
  assign n2324 = n2308 ^ n2193 ^ n2086 ;
  assign n2325 = n2310 ^ n2182 ^ n2102 ;
  assign n2326 = n2311 ^ n2160 ^ n2091 ;
  assign n2327 = n2269 ^ n2256 ^ n261 ;
  assign n2328 = ( n2296 & ~n2300 ) | ( n2296 & n2302 ) | ( ~n2300 & n2302 ) ;
  assign n2329 = n2323 ^ n2269 ^ n2180 ;
  assign n2330 = n2292 ^ n2227 ^ x98 ;
  assign n2331 = n2257 ^ n217 ^ 1'b0 ;
  assign n2332 = n2269 & n2319 ;
  assign n2333 = n2321 ^ n2269 ^ n2206 ;
  assign n2334 = n2269 & n2331 ;
  assign n2335 = n2312 ^ n2173 ^ x99 ;
  assign n2336 = n2305 ^ n2269 ^ n2197 ;
  assign n2337 = n2269 & n2313 ;
  assign n2338 = n2269 & n2317 ;
  assign n2339 = n2269 ^ n2254 ^ n345 ;
  assign n2340 = n2338 ^ n2166 ^ n2014 ;
  assign n2341 = n2320 ^ n2269 ^ n2200 ;
  assign n2342 = n2269 & n2327 ;
  assign n2343 = n2342 ^ n2215 ^ n2023 ;
  assign n2344 = n2315 ^ n2269 ^ n2186 ;
  assign n2345 = n2332 ^ n2142 ^ n2106 ;
  assign n2346 = ( n136 & n2170 ) | ( n136 & n2261 ) | ( n2170 & n2261 ) ;
  assign n2347 = n2269 ^ n2243 ^ n1118 ;
  assign n2348 = n2269 & n2347 ;
  assign n2349 = n2269 & n2339 ;
  assign n2350 = n2349 ^ n2208 ^ n2038 ;
  assign n2351 = n2337 ^ n2269 ^ n2213 ;
  assign n2352 = n2348 ^ n2152 ^ n2030 ;
  assign n2353 = ~n2318 & n2346 ;
  assign n2354 = n2334 ^ n2269 ^ n2164 ;
  assign n2355 = x92 | x93 ;
  assign n2356 = ( x95 & ~n2137 ) | ( x95 & n2355 ) | ( ~n2137 & n2355 ) ;
  assign n2357 = ( ~x95 & n2139 ) | ( ~x95 & n2269 ) | ( n2139 & n2269 ) ;
  assign n2358 = ( x95 & n2139 ) | ( x95 & ~n2355 ) | ( n2139 & ~n2355 ) ;
  assign n2359 = ( n136 & n2170 ) | ( n136 & ~n2261 ) | ( n2170 & ~n2261 ) ;
  assign n2360 = ( n2170 & ~n2261 ) | ( n2170 & n2269 ) | ( ~n2261 & n2269 ) ;
  assign n2361 = x95 & n2269 ;
  assign n2362 = ( ~n2139 & n2356 ) | ( ~n2139 & n2361 ) | ( n2356 & n2361 ) ;
  assign n2363 = ~n2361 & n2362 ;
  assign n2364 = n2357 & n2358 ;
  assign n2365 = n2361 ^ n2269 ^ x96 ;
  assign n2366 = n2363 | n2365 ;
  assign n2367 = ( n2295 & ~n2359 ) | ( n2295 & n2360 ) | ( ~n2359 & n2360 ) ;
  assign n2368 = n2363 | n2364 ;
  assign n2369 = n2170 & ~n2269 ;
  assign n2370 = n2328 ^ x97 ^ 1'b0 ;
  assign n2371 = ~n2364 & n2366 ;
  assign n2372 = ( ~n2009 & n2370 ) | ( ~n2009 & n2371 ) | ( n2370 & n2371 ) ;
  assign n2373 = ( ~n1885 & n2330 ) | ( ~n1885 & n2372 ) | ( n2330 & n2372 ) ;
  assign n2374 = ( ~n1766 & n2335 ) | ( ~n1766 & n2373 ) | ( n2335 & n2373 ) ;
  assign n2375 = ( ~n1652 & n2345 ) | ( ~n1652 & n2374 ) | ( n2345 & n2374 ) ;
  assign n2376 = ( ~n1534 & n2278 ) | ( ~n1534 & n2375 ) | ( n2278 & n2375 ) ;
  assign n2377 = ( ~n1416 & n2329 ) | ( ~n1416 & n2376 ) | ( n2329 & n2376 ) ;
  assign n2378 = ( ~n1318 & n2325 ) | ( ~n1318 & n2377 ) | ( n2325 & n2377 ) ;
  assign n2379 = ( ~n1220 & n2344 ) | ( ~n1220 & n2378 ) | ( n2344 & n2378 ) ;
  assign n2380 = ( ~n1118 & n2281 ) | ( ~n1118 & n2379 ) | ( n2281 & n2379 ) ;
  assign n2381 = ( ~n1034 & n2352 ) | ( ~n1034 & n2380 ) | ( n2352 & n2380 ) ;
  assign n2382 = ( ~n941 & n2276 ) | ( ~n941 & n2381 ) | ( n2276 & n2381 ) ;
  assign n2383 = ( ~n859 & n2284 ) | ( ~n859 & n2382 ) | ( n2284 & n2382 ) ;
  assign n2384 = ( ~n785 & n2324 ) | ( ~n785 & n2383 ) | ( n2324 & n2383 ) ;
  assign n2385 = ( ~n716 & n2336 ) | ( ~n716 & n2384 ) | ( n2336 & n2384 ) ;
  assign n2386 = ( ~n640 & n2287 ) | ( ~n640 & n2385 ) | ( n2287 & n2385 ) ;
  assign n2387 = ( ~n572 & n2341 ) | ( ~n572 & n2386 ) | ( n2341 & n2386 ) ;
  assign n2388 = ( ~n514 & n2273 ) | ( ~n514 & n2387 ) | ( n2273 & n2387 ) ;
  assign n2389 = ( ~n458 & n2290 ) | ( ~n458 & n2388 ) | ( n2290 & n2388 ) ;
  assign n2390 = ( ~n399 & n2326 ) | ( ~n399 & n2389 ) | ( n2326 & n2389 ) ;
  assign n2391 = n2390 ^ n345 ^ 1'b0 ;
  assign n2392 = ( ~n345 & n2333 ) | ( ~n345 & n2390 ) | ( n2333 & n2390 ) ;
  assign n2393 = ( ~n302 & n2350 ) | ( ~n302 & n2392 ) | ( n2350 & n2392 ) ;
  assign n2394 = ( ~n261 & n2351 ) | ( ~n261 & n2393 ) | ( n2351 & n2393 ) ;
  assign n2395 = ( ~n217 & n2343 ) | ( ~n217 & n2394 ) | ( n2343 & n2394 ) ;
  assign n2396 = ( ~n179 & n2354 ) | ( ~n179 & n2395 ) | ( n2354 & n2395 ) ;
  assign n2397 = ( ~n144 & n2340 ) | ( ~n144 & n2396 ) | ( n2340 & n2396 ) ;
  assign n2398 = ( ~n134 & n2301 ) | ( ~n134 & n2397 ) | ( n2301 & n2397 ) ;
  assign n2399 = n2295 & n2398 ;
  assign n2400 = ~n136 & n2398 ;
  assign n2401 = ( ~n136 & n2367 ) | ( ~n136 & n2400 ) | ( n2367 & n2400 ) ;
  assign n2402 = n2353 | n2401 ;
  assign n2403 = n2399 | n2402 ;
  assign n2404 = n2369 | n2403 ;
  assign n2405 = n2404 ^ n2380 ^ n1034 ;
  assign n2406 = n2404 & n2405 ;
  assign n2407 = n2376 ^ n1416 ^ 1'b0 ;
  assign n2408 = n2404 & n2407 ;
  assign n2409 = n2408 ^ n2404 ^ n2329 ;
  assign n2410 = n2368 & n2404 ;
  assign n2411 = n2410 ^ n2404 ^ n2365 ;
  assign n2412 = n2404 ^ n2377 ^ n1318 ;
  assign n2413 = n2404 & n2412 ;
  assign n2414 = n2404 ^ n2389 ^ n399 ;
  assign n2415 = n2404 ^ n2373 ^ n1766 ;
  assign n2416 = n2404 & n2415 ;
  assign n2417 = n2404 & n2414 ;
  assign n2418 = n2413 ^ n2310 ^ n2183 ;
  assign n2419 = n2416 ^ n2312 ^ n2231 ;
  assign n2420 = n2417 ^ n2311 ^ n2161 ;
  assign n2421 = n2404 ^ n2381 ^ n941 ;
  assign n2422 = n2404 & n2421 ;
  assign n2423 = n2422 ^ n2275 ^ n2189 ;
  assign n2424 = n2391 & n2404 ;
  assign n2425 = n2406 ^ n2348 ^ n2156 ;
  assign n2426 = n2404 ^ n2372 ^ n1885 ;
  assign n2427 = n2404 & n2426 ;
  assign n2428 = n2404 ^ n2382 ^ n859 ;
  assign n2429 = n2427 ^ n2292 ^ n2228 ;
  assign n2430 = n2424 ^ n2404 ^ n2333 ;
  assign n2431 = n2404 & n2428 ;
  assign n2432 = n2431 ^ n2283 ^ n2209 ;
  assign n2433 = n2404 ^ n2375 ^ n1534 ;
  assign n2434 = ~n2355 & n2404 ;
  assign n2435 = n2378 ^ n1220 ^ 1'b0 ;
  assign n2436 = n2395 ^ n179 ^ 1'b0 ;
  assign n2437 = n2393 ^ n261 ^ 1'b0 ;
  assign n2438 = n2404 & n2435 ;
  assign n2439 = n2438 ^ n2404 ^ n2344 ;
  assign n2440 = ( n2295 & n2353 ) | ( n2295 & ~n2369 ) | ( n2353 & ~n2369 ) ;
  assign n2441 = n2404 & n2437 ;
  assign n2442 = n2353 | n2369 ;
  assign n2443 = n2386 ^ n572 ^ 1'b0 ;
  assign n2444 = n2397 ^ n134 ^ 1'b0 ;
  assign n2445 = n2404 & n2444 ;
  assign n2446 = n2404 & n2443 ;
  assign n2447 = n2446 ^ n2404 ^ n2341 ;
  assign n2448 = ( x88 & x89 ) | ( x88 & ~n2369 ) | ( x89 & ~n2369 ) ;
  assign n2449 = n2404 ^ n2374 ^ n1652 ;
  assign n2450 = n2404 ^ n2379 ^ n1118 ;
  assign n2451 = n2404 & n2450 ;
  assign n2452 = n2404 ^ n2394 ^ n217 ;
  assign n2453 = ( x90 & ~n2369 ) | ( x90 & n2448 ) | ( ~n2369 & n2448 ) ;
  assign n2454 = n2269 & ~n2403 ;
  assign n2455 = n2451 ^ n2280 ^ n2155 ;
  assign n2456 = n2404 ^ n2383 ^ n785 ;
  assign n2457 = n2404 & n2456 ;
  assign n2458 = ( n2398 & n2399 ) | ( n2398 & ~n2404 ) | ( n2399 & ~n2404 ) ;
  assign n2459 = n2445 ^ n2404 ^ n2301 ;
  assign n2460 = n2404 ^ n2385 ^ n640 ;
  assign n2461 = n2404 & n2452 ;
  assign n2462 = n2457 ^ n2308 ^ n2194 ;
  assign n2463 = ( n136 & n2295 ) | ( n136 & n2398 ) | ( n2295 & n2398 ) ;
  assign n2464 = ~n2458 & n2463 ;
  assign n2465 = ( n2295 & ~n2398 ) | ( n2295 & n2404 ) | ( ~n2398 & n2404 ) ;
  assign n2466 = n2461 ^ n2342 ^ n2216 ;
  assign n2467 = n2384 ^ n716 ^ 1'b0 ;
  assign n2468 = ( ~n2399 & n2442 ) | ( ~n2399 & n2453 ) | ( n2442 & n2453 ) ;
  assign n2469 = ~n2442 & n2468 ;
  assign n2470 = n2404 ^ n2396 ^ n144 ;
  assign n2471 = n2295 & ~n2398 ;
  assign n2472 = ~n2403 & n2440 ;
  assign n2473 = ( n2459 & n2465 ) | ( n2459 & ~n2471 ) | ( n2465 & ~n2471 ) ;
  assign n2474 = n2434 | n2454 ;
  assign n2475 = n2404 & n2470 ;
  assign n2476 = n2404 & n2436 ;
  assign n2477 = n2476 ^ n2404 ^ n2354 ;
  assign n2478 = n2404 & n2449 ;
  assign n2479 = n2404 & n2467 ;
  assign n2480 = n2479 ^ n2404 ^ n2336 ;
  assign n2481 = n2404 & n2433 ;
  assign n2482 = n2404 ^ n2388 ^ n458 ;
  assign n2483 = n2481 ^ n2277 ^ n2177 ;
  assign n2484 = n2404 & n2482 ;
  assign n2485 = n2484 ^ n2289 ^ n2158 ;
  assign n2486 = n2478 ^ n2332 ^ n2174 ;
  assign n2487 = n2404 & n2460 ;
  assign n2488 = n2487 ^ n2286 ^ n2147 ;
  assign n2489 = n2475 ^ n2338 ^ n2167 ;
  assign n2490 = n2404 ^ n2371 ^ n2009 ;
  assign n2491 = n2404 & n2490 ;
  assign n2492 = n2404 ^ n2387 ^ n514 ;
  assign n2493 = n2404 ^ n2392 ^ n302 ;
  assign n2494 = n2404 & n2493 ;
  assign n2495 = n2404 & n2492 ;
  assign n2496 = n2491 ^ n2328 ^ x97 ;
  assign n2497 = n2494 ^ n2349 ^ n2210 ;
  assign n2498 = n2441 ^ n2404 ^ n2351 ;
  assign n2499 = n2495 ^ n2272 ^ n2203 ;
  assign n2500 = x92 & n2404 ;
  assign n2501 = x90 | x91 ;
  assign n2502 = n2500 ^ n2404 ^ x93 ;
  assign n2503 = ( x92 & ~n2267 ) | ( x92 & n2501 ) | ( ~n2267 & n2501 ) ;
  assign n2504 = ( ~n2269 & n2500 ) | ( ~n2269 & n2503 ) | ( n2500 & n2503 ) ;
  assign n2505 = x92 | n2501 ;
  assign n2506 = ~n2500 & n2504 ;
  assign n2507 = ( n2269 & n2500 ) | ( n2269 & ~n2505 ) | ( n2500 & ~n2505 ) ;
  assign n2508 = n2502 | n2506 ;
  assign n2509 = ~n2507 & n2508 ;
  assign n2510 = n2506 | n2507 ;
  assign n2511 = n2474 ^ x95 ^ 1'b0 ;
  assign n2512 = ( ~n2139 & n2509 ) | ( ~n2139 & n2511 ) | ( n2509 & n2511 ) ;
  assign n2513 = ( ~n2009 & n2411 ) | ( ~n2009 & n2512 ) | ( n2411 & n2512 ) ;
  assign n2514 = ( ~n1885 & n2496 ) | ( ~n1885 & n2513 ) | ( n2496 & n2513 ) ;
  assign n2515 = ( ~n1766 & n2429 ) | ( ~n1766 & n2514 ) | ( n2429 & n2514 ) ;
  assign n2516 = ( ~n1652 & n2419 ) | ( ~n1652 & n2515 ) | ( n2419 & n2515 ) ;
  assign n2517 = ( ~n1534 & n2486 ) | ( ~n1534 & n2516 ) | ( n2486 & n2516 ) ;
  assign n2518 = ( ~n1416 & n2483 ) | ( ~n1416 & n2517 ) | ( n2483 & n2517 ) ;
  assign n2519 = ( ~n1318 & n2409 ) | ( ~n1318 & n2518 ) | ( n2409 & n2518 ) ;
  assign n2520 = ( ~n1220 & n2418 ) | ( ~n1220 & n2519 ) | ( n2418 & n2519 ) ;
  assign n2521 = ( ~n1118 & n2439 ) | ( ~n1118 & n2520 ) | ( n2439 & n2520 ) ;
  assign n2522 = ( ~n1034 & n2455 ) | ( ~n1034 & n2521 ) | ( n2455 & n2521 ) ;
  assign n2523 = ( ~n941 & n2425 ) | ( ~n941 & n2522 ) | ( n2425 & n2522 ) ;
  assign n2524 = ( ~n859 & n2423 ) | ( ~n859 & n2523 ) | ( n2423 & n2523 ) ;
  assign n2525 = ( ~n785 & n2432 ) | ( ~n785 & n2524 ) | ( n2432 & n2524 ) ;
  assign n2526 = ( ~n716 & n2462 ) | ( ~n716 & n2525 ) | ( n2462 & n2525 ) ;
  assign n2527 = ( ~n640 & n2480 ) | ( ~n640 & n2526 ) | ( n2480 & n2526 ) ;
  assign n2528 = ( ~n572 & n2488 ) | ( ~n572 & n2527 ) | ( n2488 & n2527 ) ;
  assign n2529 = ( ~n514 & n2447 ) | ( ~n514 & n2528 ) | ( n2447 & n2528 ) ;
  assign n2530 = ( ~n458 & n2499 ) | ( ~n458 & n2529 ) | ( n2499 & n2529 ) ;
  assign n2531 = ( ~n399 & n2485 ) | ( ~n399 & n2530 ) | ( n2485 & n2530 ) ;
  assign n2532 = ( ~n345 & n2420 ) | ( ~n345 & n2531 ) | ( n2420 & n2531 ) ;
  assign n2533 = ( ~n302 & n2430 ) | ( ~n302 & n2532 ) | ( n2430 & n2532 ) ;
  assign n2534 = ( ~n261 & n2497 ) | ( ~n261 & n2533 ) | ( n2497 & n2533 ) ;
  assign n2535 = ( ~n217 & n2498 ) | ( ~n217 & n2534 ) | ( n2498 & n2534 ) ;
  assign n2536 = ( ~n179 & n2466 ) | ( ~n179 & n2535 ) | ( n2466 & n2535 ) ;
  assign n2537 = ( ~n144 & n2477 ) | ( ~n144 & n2536 ) | ( n2477 & n2536 ) ;
  assign n2538 = ( ~n134 & n2489 ) | ( ~n134 & n2537 ) | ( n2489 & n2537 ) ;
  assign n2539 = n2459 & n2538 ;
  assign n2540 = ( ~x30 & n2473 ) | ( ~x30 & n2538 ) | ( n2473 & n2538 ) ;
  assign n2541 = ~n136 & n2540 ;
  assign n2542 = n2464 | n2539 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = n2472 | n2543 ;
  assign n2545 = n2544 ^ n2537 ^ n134 ;
  assign n2546 = n2544 ^ n2514 ^ n1766 ;
  assign n2547 = n2544 ^ n2516 ^ n1534 ;
  assign n2548 = n2544 & n2545 ;
  assign n2549 = n2510 & n2544 ;
  assign n2550 = n2549 ^ n2544 ^ n2502 ;
  assign n2551 = n2544 & n2546 ;
  assign n2552 = n2551 ^ n2427 ^ n2330 ;
  assign n2553 = ( x90 & n2401 ) | ( x90 & n2544 ) | ( n2401 & n2544 ) ;
  assign n2554 = ( ~n2401 & n2469 ) | ( ~n2401 & n2553 ) | ( n2469 & n2553 ) ;
  assign n2555 = ~n2553 & n2554 ;
  assign n2556 = n2544 ^ n2515 ^ n1652 ;
  assign n2557 = n2544 & n2556 ;
  assign n2558 = n2544 ^ n2531 ^ n345 ;
  assign n2559 = n2544 & n2558 ;
  assign n2560 = n2544 ^ n2525 ^ n716 ;
  assign n2561 = n2544 & n2560 ;
  assign n2562 = n2557 ^ n2416 ^ n2335 ;
  assign n2563 = n2561 ^ n2457 ^ n2324 ;
  assign n2564 = n2559 ^ n2417 ^ n2326 ;
  assign n2565 = n2544 ^ n2527 ^ n572 ;
  assign n2566 = n2534 ^ n217 ^ 1'b0 ;
  assign n2567 = n2544 ^ n2529 ^ n458 ;
  assign n2568 = n2544 & n2565 ;
  assign n2569 = n2544 & n2567 ;
  assign n2570 = n2568 ^ n2487 ^ n2287 ;
  assign n2571 = n2569 ^ n2495 ^ n2273 ;
  assign n2572 = n2544 & n2566 ;
  assign n2573 = n2544 ^ n2530 ^ n399 ;
  assign n2574 = n2572 ^ n2544 ^ n2498 ;
  assign n2575 = n2544 & n2573 ;
  assign n2576 = n2544 & n2547 ;
  assign n2577 = n2575 ^ n2484 ^ n2290 ;
  assign n2578 = n2548 ^ n2475 ^ n2340 ;
  assign n2579 = n2576 ^ n2478 ^ n2345 ;
  assign n2580 = n2518 ^ n1318 ^ 1'b0 ;
  assign n2581 = n2544 & n2580 ;
  assign n2582 = n2581 ^ n2544 ^ n2409 ;
  assign n2583 = ( n2404 & n2464 ) | ( n2404 & ~n2472 ) | ( n2464 & ~n2472 ) ;
  assign n2584 = n2544 ^ n2513 ^ n1885 ;
  assign n2585 = ~n2501 & n2544 ;
  assign n2586 = n2532 ^ n302 ^ 1'b0 ;
  assign n2587 = n2544 & n2586 ;
  assign n2588 = n2587 ^ n2544 ^ n2430 ;
  assign n2589 = n2544 ^ n2521 ^ n1034 ;
  assign n2590 = n2543 & ~n2585 ;
  assign n2591 = n2526 ^ n640 ^ 1'b0 ;
  assign n2592 = n2520 ^ n1118 ^ 1'b0 ;
  assign n2593 = n2512 ^ n2009 ^ 1'b0 ;
  assign n2594 = n2544 & n2589 ;
  assign n2595 = n2594 ^ n2451 ^ n2281 ;
  assign n2596 = n2544 & n2591 ;
  assign n2597 = n2544 ^ n2524 ^ n785 ;
  assign n2598 = ( n2459 & n2464 ) | ( n2459 & ~n2472 ) | ( n2464 & ~n2472 ) ;
  assign n2599 = n2528 ^ n514 ^ 1'b0 ;
  assign n2600 = n2544 & n2599 ;
  assign n2601 = n2600 ^ n2544 ^ n2447 ;
  assign n2602 = n2544 ^ n2533 ^ n261 ;
  assign n2603 = ( n136 & n2459 ) | ( n136 & n2538 ) | ( n2459 & n2538 ) ;
  assign n2604 = n2544 ^ n2519 ^ n1220 ;
  assign n2605 = ~n2543 & n2598 ;
  assign n2606 = ( ~n2459 & n2538 ) | ( ~n2459 & n2544 ) | ( n2538 & n2544 ) ;
  assign n2607 = n2596 ^ n2544 ^ n2480 ;
  assign n2608 = ~n2459 & n2538 ;
  assign n2609 = n2544 ^ n2522 ^ n941 ;
  assign n2610 = n2544 ^ n2535 ^ n179 ;
  assign n2611 = n2544 & n2593 ;
  assign n2612 = n2544 & n2592 ;
  assign n2613 = ( n2538 & n2539 ) | ( n2538 & ~n2544 ) | ( n2539 & ~n2544 ) ;
  assign n2614 = ( x86 & x87 ) | ( x86 & ~n2472 ) | ( x87 & ~n2472 ) ;
  assign n2615 = n2603 & ~n2613 ;
  assign n2616 = n2472 | n2539 ;
  assign n2617 = ( x88 & ~n2472 ) | ( x88 & n2614 ) | ( ~n2472 & n2614 ) ;
  assign n2618 = n2536 ^ n144 ^ 1'b0 ;
  assign n2619 = n2544 & n2597 ;
  assign n2620 = n2619 ^ n2431 ^ n2284 ;
  assign n2621 = n2544 ^ n2523 ^ n859 ;
  assign n2622 = n2544 & n2621 ;
  assign n2623 = ( ~n2464 & n2616 ) | ( ~n2464 & n2617 ) | ( n2616 & n2617 ) ;
  assign n2624 = ~n2616 & n2623 ;
  assign n2625 = n2622 ^ n2422 ^ n2276 ;
  assign n2626 = n2544 & n2610 ;
  assign n2627 = ( n2578 & n2606 ) | ( n2578 & ~n2608 ) | ( n2606 & ~n2608 ) ;
  assign n2628 = n2544 & n2609 ;
  assign n2629 = ( n2583 & n2585 ) | ( n2583 & ~n2590 ) | ( n2585 & ~n2590 ) ;
  assign n2630 = n2626 ^ n2461 ^ n2343 ;
  assign n2631 = n2628 ^ n2406 ^ n2352 ;
  assign n2632 = n2612 ^ n2544 ^ n2439 ;
  assign n2633 = n2544 ^ n2517 ^ n1416 ;
  assign n2634 = n2544 & n2633 ;
  assign n2635 = n2634 ^ n2481 ^ n2278 ;
  assign n2636 = n2544 & n2584 ;
  assign n2637 = n2636 ^ n2491 ^ n2370 ;
  assign n2638 = n2544 & n2602 ;
  assign n2639 = n2638 ^ n2494 ^ n2350 ;
  assign n2640 = n2544 & n2604 ;
  assign n2641 = n2640 ^ n2413 ^ n2325 ;
  assign n2642 = n2544 & n2618 ;
  assign n2643 = n2642 ^ n2544 ^ n2477 ;
  assign n2644 = n2629 ^ x92 ^ 1'b0 ;
  assign n2645 = x88 | x89 ;
  assign n2646 = ( x90 & n2404 ) | ( x90 & ~n2645 ) | ( n2404 & ~n2645 ) ;
  assign n2647 = ( ~x90 & n2404 ) | ( ~x90 & n2544 ) | ( n2404 & n2544 ) ;
  assign n2648 = n2646 & n2647 ;
  assign n2649 = ~x90 & n2544 ;
  assign n2650 = n2649 ^ x91 ^ 1'b0 ;
  assign n2651 = n2555 | n2650 ;
  assign n2652 = ~n2648 & n2651 ;
  assign n2653 = ( ~n2269 & n2644 ) | ( ~n2269 & n2652 ) | ( n2644 & n2652 ) ;
  assign n2654 = ( ~n2139 & n2550 ) | ( ~n2139 & n2653 ) | ( n2550 & n2653 ) ;
  assign n2655 = n2544 ^ n2509 ^ n2139 ;
  assign n2656 = n2544 & n2655 ;
  assign n2657 = n2656 ^ n2474 ^ x95 ;
  assign n2658 = ( ~n2009 & n2654 ) | ( ~n2009 & n2657 ) | ( n2654 & n2657 ) ;
  assign n2659 = n2611 ^ n2544 ^ n2411 ;
  assign n2660 = ( ~n1885 & n2658 ) | ( ~n1885 & n2659 ) | ( n2658 & n2659 ) ;
  assign n2661 = ( ~n1766 & n2637 ) | ( ~n1766 & n2660 ) | ( n2637 & n2660 ) ;
  assign n2662 = ( ~n1652 & n2552 ) | ( ~n1652 & n2661 ) | ( n2552 & n2661 ) ;
  assign n2663 = ( ~n1534 & n2562 ) | ( ~n1534 & n2662 ) | ( n2562 & n2662 ) ;
  assign n2664 = ( ~n1416 & n2579 ) | ( ~n1416 & n2663 ) | ( n2579 & n2663 ) ;
  assign n2665 = ( ~n1318 & n2635 ) | ( ~n1318 & n2664 ) | ( n2635 & n2664 ) ;
  assign n2666 = ( ~n1220 & n2582 ) | ( ~n1220 & n2665 ) | ( n2582 & n2665 ) ;
  assign n2667 = ( ~n1118 & n2641 ) | ( ~n1118 & n2666 ) | ( n2641 & n2666 ) ;
  assign n2668 = ( ~n1034 & n2632 ) | ( ~n1034 & n2667 ) | ( n2632 & n2667 ) ;
  assign n2669 = ( ~n941 & n2595 ) | ( ~n941 & n2668 ) | ( n2595 & n2668 ) ;
  assign n2670 = ( ~n859 & n2631 ) | ( ~n859 & n2669 ) | ( n2631 & n2669 ) ;
  assign n2671 = ( ~n785 & n2625 ) | ( ~n785 & n2670 ) | ( n2625 & n2670 ) ;
  assign n2672 = ( ~n716 & n2620 ) | ( ~n716 & n2671 ) | ( n2620 & n2671 ) ;
  assign n2673 = ( ~n640 & n2563 ) | ( ~n640 & n2672 ) | ( n2563 & n2672 ) ;
  assign n2674 = ( ~n572 & n2607 ) | ( ~n572 & n2673 ) | ( n2607 & n2673 ) ;
  assign n2675 = ( ~n514 & n2570 ) | ( ~n514 & n2674 ) | ( n2570 & n2674 ) ;
  assign n2676 = ( ~n458 & n2601 ) | ( ~n458 & n2675 ) | ( n2601 & n2675 ) ;
  assign n2677 = ( ~n399 & n2571 ) | ( ~n399 & n2676 ) | ( n2571 & n2676 ) ;
  assign n2678 = ( ~n345 & n2577 ) | ( ~n345 & n2677 ) | ( n2577 & n2677 ) ;
  assign n2679 = ( ~n302 & n2564 ) | ( ~n302 & n2678 ) | ( n2564 & n2678 ) ;
  assign n2680 = ( ~n261 & n2588 ) | ( ~n261 & n2679 ) | ( n2588 & n2679 ) ;
  assign n2681 = ( ~n217 & n2639 ) | ( ~n217 & n2680 ) | ( n2639 & n2680 ) ;
  assign n2682 = ( ~n179 & n2574 ) | ( ~n179 & n2681 ) | ( n2574 & n2681 ) ;
  assign n2683 = ( ~n144 & n2630 ) | ( ~n144 & n2682 ) | ( n2630 & n2682 ) ;
  assign n2684 = ( ~n134 & n2643 ) | ( ~n134 & n2683 ) | ( n2643 & n2683 ) ;
  assign n2685 = n2578 & n2684 ;
  assign n2686 = ( ~x30 & n2627 ) | ( ~x30 & n2684 ) | ( n2627 & n2684 ) ;
  assign n2687 = ~n136 & n2686 ;
  assign n2688 = n2685 | n2687 ;
  assign n2689 = n2615 | n2688 ;
  assign n2690 = n2605 | n2689 ;
  assign n2691 = ~n2645 & n2690 ;
  assign n2692 = ( n2605 & n2615 ) | ( n2605 & ~n2691 ) | ( n2615 & ~n2691 ) ;
  assign n2693 = n2544 & ~n2688 ;
  assign n2694 = n2691 | n2693 ;
  assign n2695 = ( n2691 & ~n2692 ) | ( n2691 & n2694 ) | ( ~n2692 & n2694 ) ;
  assign n2696 = ( n2555 & ~n2648 ) | ( n2555 & n2690 ) | ( ~n2648 & n2690 ) ;
  assign n2697 = ~n2555 & n2696 ;
  assign n2698 = n2690 ^ n2661 ^ n1652 ;
  assign n2699 = n2690 & n2698 ;
  assign n2700 = n2699 ^ n2551 ^ n2429 ;
  assign n2701 = n2690 ^ n2664 ^ n1318 ;
  assign n2702 = n2690 & n2701 ;
  assign n2703 = n2702 ^ n2634 ^ n2483 ;
  assign n2704 = n2690 ^ n2668 ^ n941 ;
  assign n2705 = n2690 & n2704 ;
  assign n2706 = n2705 ^ n2594 ^ n2455 ;
  assign n2707 = n2690 ^ n2670 ^ n785 ;
  assign n2708 = n2690 & n2707 ;
  assign n2709 = n2708 ^ n2622 ^ n2423 ;
  assign n2710 = n2690 ^ n2671 ^ n716 ;
  assign n2711 = n2690 & n2710 ;
  assign n2712 = n2711 ^ n2619 ^ n2432 ;
  assign n2713 = n2690 ^ n2674 ^ n514 ;
  assign n2714 = n2690 & n2713 ;
  assign n2715 = n2714 ^ n2568 ^ n2488 ;
  assign n2716 = n2690 ^ n2660 ^ n1766 ;
  assign n2717 = n2690 & n2716 ;
  assign n2718 = n2690 ^ n2654 ^ n2009 ;
  assign n2719 = n2717 ^ n2636 ^ n2496 ;
  assign n2720 = ( x88 & n2541 ) | ( x88 & n2690 ) | ( n2541 & n2690 ) ;
  assign n2721 = ( ~n2541 & n2624 ) | ( ~n2541 & n2720 ) | ( n2624 & n2720 ) ;
  assign n2722 = n2658 ^ n1885 ^ 1'b0 ;
  assign n2723 = n2690 ^ n2680 ^ n217 ;
  assign n2724 = n2681 ^ n179 ^ 1'b0 ;
  assign n2725 = n2690 ^ n2669 ^ n859 ;
  assign n2726 = n2690 ^ n2662 ^ n1534 ;
  assign n2727 = n2653 ^ n2139 ^ 1'b0 ;
  assign n2728 = n2690 ^ n2663 ^ n1416 ;
  assign n2729 = n2673 ^ n572 ^ 1'b0 ;
  assign n2730 = n2690 ^ n2666 ^ n1118 ;
  assign n2731 = n2690 & n2727 ;
  assign n2732 = n2731 ^ n2690 ^ n2550 ;
  assign n2733 = n2683 ^ n134 ^ 1'b0 ;
  assign n2734 = n2675 ^ n458 ^ 1'b0 ;
  assign n2735 = n2679 ^ n261 ^ 1'b0 ;
  assign n2736 = n2690 ^ n2682 ^ n144 ;
  assign n2737 = n2690 ^ n2678 ^ n302 ;
  assign n2738 = n2690 ^ n2677 ^ n345 ;
  assign n2739 = n2690 ^ n2672 ^ n640 ;
  assign n2740 = n2690 ^ n2676 ^ n399 ;
  assign n2741 = n2690 & n2726 ;
  assign n2742 = n2741 ^ n2557 ^ n2419 ;
  assign n2743 = n2690 & n2728 ;
  assign n2744 = n2690 & n2735 ;
  assign n2745 = n2743 ^ n2576 ^ n2486 ;
  assign n2746 = n2690 & n2737 ;
  assign n2747 = n2746 ^ n2559 ^ n2420 ;
  assign n2748 = n2690 & n2723 ;
  assign n2749 = n2748 ^ n2638 ^ n2497 ;
  assign n2750 = n2690 & n2736 ;
  assign n2751 = n2750 ^ n2626 ^ n2466 ;
  assign n2752 = n2690 & n2724 ;
  assign n2753 = n2690 & n2738 ;
  assign n2754 = n2753 ^ n2575 ^ n2485 ;
  assign n2755 = n2690 & n2740 ;
  assign n2756 = n2690 & n2718 ;
  assign n2757 = n2755 ^ n2569 ^ n2499 ;
  assign n2758 = n2756 ^ n2656 ^ n2511 ;
  assign n2759 = ~n2720 & n2721 ;
  assign n2760 = n2690 & n2733 ;
  assign n2761 = n2690 & n2729 ;
  assign n2762 = n2667 ^ n1034 ^ 1'b0 ;
  assign n2763 = n2690 & n2762 ;
  assign n2764 = n2763 ^ n2690 ^ n2632 ;
  assign n2765 = n2690 & n2734 ;
  assign n2766 = n2765 ^ n2690 ^ n2601 ;
  assign n2767 = n2690 & n2722 ;
  assign n2768 = n2767 ^ n2690 ^ n2659 ;
  assign n2769 = n2744 ^ n2690 ^ n2588 ;
  assign n2770 = n2690 & n2730 ;
  assign n2771 = n2770 ^ n2640 ^ n2418 ;
  assign n2772 = n2752 ^ n2690 ^ n2574 ;
  assign n2773 = n2760 ^ n2690 ^ n2643 ;
  assign n2774 = n2690 & n2739 ;
  assign n2775 = n2690 & n2725 ;
  assign n2776 = n2775 ^ n2628 ^ n2425 ;
  assign n2777 = n2774 ^ n2561 ^ n2462 ;
  assign n2778 = ~x88 & n2690 ;
  assign n2779 = ( n2684 & n2685 ) | ( n2684 & ~n2690 ) | ( n2685 & ~n2690 ) ;
  assign n2780 = n2269 & n2652 ;
  assign n2781 = ( n136 & n2578 ) | ( n136 & n2684 ) | ( n2578 & n2684 ) ;
  assign n2782 = n2778 ^ x89 ^ 1'b0 ;
  assign n2783 = n2759 | n2782 ;
  assign n2784 = ( ~n2269 & n2690 ) | ( ~n2269 & n2780 ) | ( n2690 & n2780 ) ;
  assign n2785 = n2665 ^ n1220 ^ 1'b0 ;
  assign n2786 = ( ~n2652 & n2780 ) | ( ~n2652 & n2784 ) | ( n2780 & n2784 ) ;
  assign n2787 = n2578 & ~n2684 ;
  assign n2788 = n2690 & n2785 ;
  assign n2789 = ~n2779 & n2781 ;
  assign n2790 = n2788 ^ n2690 ^ n2582 ;
  assign n2791 = n2761 ^ n2690 ^ n2607 ;
  assign n2792 = x86 | x87 ;
  assign n2793 = n2695 ^ x90 ^ 1'b0 ;
  assign n2794 = ( ~x88 & n2544 ) | ( ~x88 & n2690 ) | ( n2544 & n2690 ) ;
  assign n2795 = n2697 ^ n2649 ^ x91 ;
  assign n2796 = ( n2578 & ~n2690 ) | ( n2578 & n2789 ) | ( ~n2690 & n2789 ) ;
  assign n2797 = n2786 ^ n2629 ^ x92 ;
  assign n2798 = ( x88 & n2544 ) | ( x88 & ~n2792 ) | ( n2544 & ~n2792 ) ;
  assign n2799 = n2794 & n2798 ;
  assign n2800 = n2783 & ~n2799 ;
  assign n2801 = ( ~n2404 & n2793 ) | ( ~n2404 & n2800 ) | ( n2793 & n2800 ) ;
  assign n2802 = ( ~n2269 & n2795 ) | ( ~n2269 & n2801 ) | ( n2795 & n2801 ) ;
  assign n2803 = ( ~n2139 & n2797 ) | ( ~n2139 & n2802 ) | ( n2797 & n2802 ) ;
  assign n2804 = ( ~n2009 & n2732 ) | ( ~n2009 & n2803 ) | ( n2732 & n2803 ) ;
  assign n2805 = ( ~n1885 & n2758 ) | ( ~n1885 & n2804 ) | ( n2758 & n2804 ) ;
  assign n2806 = ( ~n1766 & n2768 ) | ( ~n1766 & n2805 ) | ( n2768 & n2805 ) ;
  assign n2807 = ( ~n1652 & n2719 ) | ( ~n1652 & n2806 ) | ( n2719 & n2806 ) ;
  assign n2808 = ( ~n1534 & n2700 ) | ( ~n1534 & n2807 ) | ( n2700 & n2807 ) ;
  assign n2809 = ( ~n1416 & n2742 ) | ( ~n1416 & n2808 ) | ( n2742 & n2808 ) ;
  assign n2810 = ( ~n1318 & n2745 ) | ( ~n1318 & n2809 ) | ( n2745 & n2809 ) ;
  assign n2811 = ( ~n1220 & n2703 ) | ( ~n1220 & n2810 ) | ( n2703 & n2810 ) ;
  assign n2812 = ( ~n1118 & n2790 ) | ( ~n1118 & n2811 ) | ( n2790 & n2811 ) ;
  assign n2813 = ( ~n1034 & n2771 ) | ( ~n1034 & n2812 ) | ( n2771 & n2812 ) ;
  assign n2814 = ( ~n941 & n2764 ) | ( ~n941 & n2813 ) | ( n2764 & n2813 ) ;
  assign n2815 = ( n2578 & ~n2684 ) | ( n2578 & n2690 ) | ( ~n2684 & n2690 ) ;
  assign n2816 = ( n2773 & ~n2787 ) | ( n2773 & n2815 ) | ( ~n2787 & n2815 ) ;
  assign n2817 = ( ~n859 & n2706 ) | ( ~n859 & n2814 ) | ( n2706 & n2814 ) ;
  assign n2818 = ( ~n785 & n2776 ) | ( ~n785 & n2817 ) | ( n2776 & n2817 ) ;
  assign n2819 = ( ~n716 & n2709 ) | ( ~n716 & n2818 ) | ( n2709 & n2818 ) ;
  assign n2820 = ( ~n640 & n2712 ) | ( ~n640 & n2819 ) | ( n2712 & n2819 ) ;
  assign n2821 = ( ~n572 & n2777 ) | ( ~n572 & n2820 ) | ( n2777 & n2820 ) ;
  assign n2822 = ( ~n514 & n2791 ) | ( ~n514 & n2821 ) | ( n2791 & n2821 ) ;
  assign n2823 = ( ~n458 & n2715 ) | ( ~n458 & n2822 ) | ( n2715 & n2822 ) ;
  assign n2824 = ( ~n399 & n2766 ) | ( ~n399 & n2823 ) | ( n2766 & n2823 ) ;
  assign n2825 = n2823 ^ n399 ^ 1'b0 ;
  assign n2826 = ( ~n345 & n2757 ) | ( ~n345 & n2824 ) | ( n2757 & n2824 ) ;
  assign n2827 = n2821 ^ n514 ^ 1'b0 ;
  assign n2828 = ( ~n302 & n2754 ) | ( ~n302 & n2826 ) | ( n2754 & n2826 ) ;
  assign n2829 = ( ~n261 & n2747 ) | ( ~n261 & n2828 ) | ( n2747 & n2828 ) ;
  assign n2830 = ( ~n217 & n2769 ) | ( ~n217 & n2829 ) | ( n2769 & n2829 ) ;
  assign n2831 = ( ~n179 & n2749 ) | ( ~n179 & n2830 ) | ( n2749 & n2830 ) ;
  assign n2832 = ( ~n144 & n2772 ) | ( ~n144 & n2831 ) | ( n2772 & n2831 ) ;
  assign n2833 = ( ~n134 & n2751 ) | ( ~n134 & n2832 ) | ( n2751 & n2832 ) ;
  assign n2834 = ( ~x30 & n2816 ) | ( ~x30 & n2833 ) | ( n2816 & n2833 ) ;
  assign n2835 = ~n136 & n2834 ;
  assign n2836 = ~n2773 & n2833 ;
  assign n2837 = ( n2833 & n2835 ) | ( n2833 & ~n2836 ) | ( n2835 & ~n2836 ) ;
  assign n2838 = n2789 | n2837 ;
  assign n2839 = n2796 | n2838 ;
  assign n2840 = n2839 ^ n2832 ^ n134 ;
  assign n2841 = n2839 & n2840 ;
  assign n2842 = n2841 ^ n2750 ^ n2630 ;
  assign n2843 = ~n2792 & n2839 ;
  assign n2844 = n2690 & ~n2838 ;
  assign n2845 = n2843 | n2844 ;
  assign n2846 = ( n2759 & ~n2799 ) | ( n2759 & n2839 ) | ( ~n2799 & n2839 ) ;
  assign n2847 = ~n2759 & n2846 ;
  assign n2848 = n2839 ^ n2801 ^ n2269 ;
  assign n2849 = n2839 ^ n2808 ^ n1416 ;
  assign n2850 = n2839 & n2849 ;
  assign n2851 = n2850 ^ n2741 ^ n2562 ;
  assign n2852 = n2839 ^ n2809 ^ n1318 ;
  assign n2853 = n2839 & n2852 ;
  assign n2854 = n2853 ^ n2743 ^ n2579 ;
  assign n2855 = n2839 ^ n2812 ^ n1034 ;
  assign n2856 = n2839 & n2855 ;
  assign n2857 = n2856 ^ n2770 ^ n2641 ;
  assign n2858 = n2839 ^ n2814 ^ n859 ;
  assign n2859 = n2839 & n2858 ;
  assign n2860 = n2839 & n2848 ;
  assign n2861 = n2860 ^ n2697 ^ n2650 ;
  assign n2862 = n2859 ^ n2705 ^ n2595 ;
  assign n2863 = n2839 ^ n2820 ^ n572 ;
  assign n2864 = n2839 & n2863 ;
  assign n2865 = n2864 ^ n2774 ^ n2563 ;
  assign n2866 = n2827 & n2839 ;
  assign n2867 = n2866 ^ n2839 ^ n2791 ;
  assign n2868 = n2839 ^ n2822 ^ n458 ;
  assign n2869 = n2839 & n2868 ;
  assign n2870 = n2869 ^ n2714 ^ n2570 ;
  assign n2871 = n2825 & n2839 ;
  assign n2872 = n2871 ^ n2839 ^ n2766 ;
  assign n2873 = n2839 ^ n2824 ^ n345 ;
  assign n2874 = n2839 & n2873 ;
  assign n2875 = n2874 ^ n2755 ^ n2571 ;
  assign n2876 = n2839 ^ n2826 ^ n302 ;
  assign n2877 = n2839 & n2876 ;
  assign n2878 = n2877 ^ n2753 ^ n2577 ;
  assign n2879 = n2839 ^ n2828 ^ n261 ;
  assign n2880 = n2839 & n2879 ;
  assign n2881 = n2880 ^ n2746 ^ n2564 ;
  assign n2882 = n2829 ^ n217 ^ 1'b0 ;
  assign n2883 = n2839 & n2882 ;
  assign n2884 = n2883 ^ n2839 ^ n2769 ;
  assign n2885 = n2831 ^ n144 ^ 1'b0 ;
  assign n2886 = n2839 & n2885 ;
  assign n2887 = n2886 ^ n2839 ^ n2772 ;
  assign n2888 = n2847 ^ n2778 ^ x89 ;
  assign n2889 = n2839 ^ n2800 ^ n2404 ;
  assign n2890 = n2839 & n2889 ;
  assign n2891 = n2890 ^ n2695 ^ x90 ;
  assign n2892 = n2839 ^ n2802 ^ n2139 ;
  assign n2893 = n2839 & n2892 ;
  assign n2894 = n2893 ^ n2786 ^ n2644 ;
  assign n2895 = n2803 ^ n2009 ^ 1'b0 ;
  assign n2896 = n2839 & n2895 ;
  assign n2897 = n2896 ^ n2839 ^ n2732 ;
  assign n2898 = n2839 ^ n2804 ^ n1885 ;
  assign n2899 = n2839 & n2898 ;
  assign n2900 = n2899 ^ n2756 ^ n2657 ;
  assign n2901 = n2839 ^ n2806 ^ n1652 ;
  assign n2902 = n2839 & n2901 ;
  assign n2903 = n2902 ^ n2717 ^ n2637 ;
  assign n2904 = n2839 ^ n2807 ^ n1534 ;
  assign n2905 = n2839 & n2904 ;
  assign n2906 = n2905 ^ n2699 ^ n2552 ;
  assign n2907 = n2839 ^ n2810 ^ n1220 ;
  assign n2908 = n2839 & n2907 ;
  assign n2909 = n2805 ^ n1766 ^ 1'b0 ;
  assign n2910 = n2839 & n2909 ;
  assign n2911 = n2910 ^ n2839 ^ n2768 ;
  assign n2912 = n2908 ^ n2702 ^ n2635 ;
  assign n2913 = n2811 ^ n1118 ^ 1'b0 ;
  assign n2914 = n2839 & n2913 ;
  assign n2915 = n2914 ^ n2839 ^ n2790 ;
  assign n2916 = n2813 ^ n941 ^ 1'b0 ;
  assign n2917 = n2839 & n2916 ;
  assign n2918 = n2917 ^ n2839 ^ n2764 ;
  assign n2919 = n2839 ^ n2817 ^ n785 ;
  assign n2920 = n2839 & n2919 ;
  assign n2921 = n2920 ^ n2775 ^ n2631 ;
  assign n2922 = n2839 ^ n2818 ^ n716 ;
  assign n2923 = n2839 & n2922 ;
  assign n2924 = n2923 ^ n2708 ^ n2625 ;
  assign n2925 = n2839 ^ n2819 ^ n640 ;
  assign n2926 = n2839 & n2925 ;
  assign n2927 = n2926 ^ n2711 ^ n2620 ;
  assign n2928 = n2839 ^ n2830 ^ n179 ;
  assign n2929 = n2839 & n2928 ;
  assign n2930 = n2929 ^ n2748 ^ n2639 ;
  assign n2931 = x84 | x85 ;
  assign n2932 = ( x86 & ~n2688 ) | ( x86 & n2931 ) | ( ~n2688 & n2931 ) ;
  assign n2933 = x86 & n2839 ;
  assign n2934 = ( ~n2690 & n2932 ) | ( ~n2690 & n2933 ) | ( n2932 & n2933 ) ;
  assign n2935 = ~n2933 & n2934 ;
  assign n2936 = n2845 ^ x88 ^ 1'b0 ;
  assign n2937 = x86 | n2931 ;
  assign n2938 = ( n2690 & n2933 ) | ( n2690 & ~n2937 ) | ( n2933 & ~n2937 ) ;
  assign n2939 = n2933 ^ n2839 ^ x87 ;
  assign n2940 = n2935 | n2939 ;
  assign n2941 = ~n2938 & n2940 ;
  assign n2942 = ( ~n2544 & n2936 ) | ( ~n2544 & n2941 ) | ( n2936 & n2941 ) ;
  assign n2943 = ( ~n2404 & n2888 ) | ( ~n2404 & n2942 ) | ( n2888 & n2942 ) ;
  assign n2944 = ( ~n2269 & n2891 ) | ( ~n2269 & n2943 ) | ( n2891 & n2943 ) ;
  assign n2945 = ( ~n2139 & n2861 ) | ( ~n2139 & n2944 ) | ( n2861 & n2944 ) ;
  assign n2946 = ( ~n2009 & n2894 ) | ( ~n2009 & n2945 ) | ( n2894 & n2945 ) ;
  assign n2947 = ( ~n1885 & n2897 ) | ( ~n1885 & n2946 ) | ( n2897 & n2946 ) ;
  assign n2948 = ( ~n1766 & n2900 ) | ( ~n1766 & n2947 ) | ( n2900 & n2947 ) ;
  assign n2949 = ( ~n1652 & n2911 ) | ( ~n1652 & n2948 ) | ( n2911 & n2948 ) ;
  assign n2950 = ( ~n1534 & n2903 ) | ( ~n1534 & n2949 ) | ( n2903 & n2949 ) ;
  assign n2951 = ( ~n1416 & n2906 ) | ( ~n1416 & n2950 ) | ( n2906 & n2950 ) ;
  assign n2952 = ( n2773 & n2833 ) | ( n2773 & ~n2839 ) | ( n2833 & ~n2839 ) ;
  assign n2953 = ( ~n1318 & n2851 ) | ( ~n1318 & n2951 ) | ( n2851 & n2951 ) ;
  assign n2954 = ( ~n1220 & n2854 ) | ( ~n1220 & n2953 ) | ( n2854 & n2953 ) ;
  assign n2955 = ( ~n1118 & n2912 ) | ( ~n1118 & n2954 ) | ( n2912 & n2954 ) ;
  assign n2956 = ( ~n1034 & n2915 ) | ( ~n1034 & n2955 ) | ( n2915 & n2955 ) ;
  assign n2957 = ( ~n941 & n2857 ) | ( ~n941 & n2956 ) | ( n2857 & n2956 ) ;
  assign n2958 = ( ~n859 & n2918 ) | ( ~n859 & n2957 ) | ( n2918 & n2957 ) ;
  assign n2959 = n2833 ^ n2773 ^ 1'b0 ;
  assign n2960 = n2833 & n2952 ;
  assign n2961 = n2935 | n2938 ;
  assign n2962 = ( ~n785 & n2862 ) | ( ~n785 & n2958 ) | ( n2862 & n2958 ) ;
  assign n2963 = ( n136 & n2773 ) | ( n136 & n2833 ) | ( n2773 & n2833 ) ;
  assign n2964 = n2773 & ~n2839 ;
  assign n2965 = ( n2773 & ~n2833 ) | ( n2773 & n2839 ) | ( ~n2833 & n2839 ) ;
  assign n2966 = ( ~n716 & n2921 ) | ( ~n716 & n2962 ) | ( n2921 & n2962 ) ;
  assign n2967 = ( ~n640 & n2924 ) | ( ~n640 & n2966 ) | ( n2924 & n2966 ) ;
  assign n2968 = ( ~n2960 & n2963 ) | ( ~n2960 & n2964 ) | ( n2963 & n2964 ) ;
  assign n2969 = n2948 ^ n1652 ^ 1'b0 ;
  assign n2970 = ( ~n572 & n2927 ) | ( ~n572 & n2967 ) | ( n2927 & n2967 ) ;
  assign n2971 = ( n2833 & ~n2959 ) | ( n2833 & n2965 ) | ( ~n2959 & n2965 ) ;
  assign n2972 = ( ~n514 & n2865 ) | ( ~n514 & n2970 ) | ( n2865 & n2970 ) ;
  assign n2973 = ( x79 & x80 ) | ( x79 & ~n2964 ) | ( x80 & ~n2964 ) ;
  assign n2974 = ( x81 & ~n2964 ) | ( x81 & n2973 ) | ( ~n2964 & n2973 ) ;
  assign n2975 = ( ~n458 & n2867 ) | ( ~n458 & n2972 ) | ( n2867 & n2972 ) ;
  assign n2976 = n2946 ^ n1885 ^ 1'b0 ;
  assign n2977 = n2972 ^ n458 ^ 1'b0 ;
  assign n2978 = n2955 ^ n1034 ^ 1'b0 ;
  assign n2979 = ( n2835 & ~n2968 ) | ( n2835 & n2971 ) | ( ~n2968 & n2971 ) ;
  assign n2980 = ( ~n399 & n2870 ) | ( ~n399 & n2975 ) | ( n2870 & n2975 ) ;
  assign n2981 = ( ~n345 & n2872 ) | ( ~n345 & n2980 ) | ( n2872 & n2980 ) ;
  assign n2982 = ( ~n302 & n2875 ) | ( ~n302 & n2981 ) | ( n2875 & n2981 ) ;
  assign n2983 = ( ~n261 & n2878 ) | ( ~n261 & n2982 ) | ( n2878 & n2982 ) ;
  assign n2984 = ( ~n217 & n2881 ) | ( ~n217 & n2983 ) | ( n2881 & n2983 ) ;
  assign n2985 = ( ~n179 & n2884 ) | ( ~n179 & n2984 ) | ( n2884 & n2984 ) ;
  assign n2986 = ( ~n144 & n2930 ) | ( ~n144 & n2985 ) | ( n2930 & n2985 ) ;
  assign n2987 = ( ~n134 & n2887 ) | ( ~n134 & n2986 ) | ( n2887 & n2986 ) ;
  assign n2988 = ( ~n136 & n2842 ) | ( ~n136 & n2987 ) | ( n2842 & n2987 ) ;
  assign n2989 = n2842 & n2987 ;
  assign n2990 = ( n2968 & n2974 ) | ( n2968 & ~n2989 ) | ( n2974 & ~n2989 ) ;
  assign n2991 = n2971 | n2988 ;
  assign n2992 = ~n136 & n2991 ;
  assign n2993 = ~n2968 & n2990 ;
  assign n2994 = n2989 | n2992 ;
  assign n2995 = n2968 | n2994 ;
  assign n2996 = n2995 ^ n2944 ^ n2139 ;
  assign n2997 = n2995 ^ n2966 ^ n640 ;
  assign n2998 = n2961 & n2995 ;
  assign n2999 = n2977 & n2995 ;
  assign n3000 = n2976 & n2995 ;
  assign n3001 = n2995 & n2997 ;
  assign n3002 = n2995 ^ n2956 ^ n941 ;
  assign n3003 = n2998 ^ n2995 ^ n2939 ;
  assign n3004 = n2995 ^ n2985 ^ n144 ;
  assign n3005 = n2995 ^ n2975 ^ n399 ;
  assign n3006 = n2995 & n3002 ;
  assign n3007 = n2969 & n2995 ;
  assign n3008 = n2995 ^ n2945 ^ n2009 ;
  assign n3009 = n2995 & n3008 ;
  assign n3010 = ~n2931 & n2995 ;
  assign n3011 = n2994 & ~n3010 ;
  assign n3012 = ( n2979 & n3010 ) | ( n2979 & ~n3011 ) | ( n3010 & ~n3011 ) ;
  assign n3013 = n2995 & n3005 ;
  assign n3014 = n2995 ^ n2970 ^ n514 ;
  assign n3015 = n2995 & n3014 ;
  assign n3016 = n2995 ^ n2958 ^ n785 ;
  assign n3017 = n2995 & n3016 ;
  assign n3018 = n2978 & n2995 ;
  assign n3019 = n2995 ^ n2983 ^ n217 ;
  assign n3020 = n2995 & n3004 ;
  assign n3021 = n2995 & n3019 ;
  assign n3022 = n2995 & n2996 ;
  assign n3023 = n2995 ^ n2981 ^ n302 ;
  assign n3024 = n2995 & n3023 ;
  assign n3025 = n3020 ^ n2929 ^ n2749 ;
  assign n3026 = n3024 ^ n2874 ^ n2757 ;
  assign n3027 = n2999 ^ n2995 ^ n2867 ;
  assign n3028 = n2995 ^ n2954 ^ n1118 ;
  assign n3029 = n2995 & n3028 ;
  assign n3030 = n3000 ^ n2995 ^ n2897 ;
  assign n3031 = n3018 ^ n2995 ^ n2915 ;
  assign n3032 = n3001 ^ n2923 ^ n2709 ;
  assign n3033 = n3022 ^ n2860 ^ n2795 ;
  assign n3034 = n3013 ^ n2869 ^ n2715 ;
  assign n3035 = n3029 ^ n2908 ^ n2703 ;
  assign n3036 = n3015 ^ n2864 ^ n2777 ;
  assign n3037 = n3007 ^ n2995 ^ n2911 ;
  assign n3038 = n3006 ^ n2856 ^ n2771 ;
  assign n3039 = n3009 ^ n2893 ^ n2797 ;
  assign n3040 = n3017 ^ n2859 ^ n2706 ;
  assign n3041 = n3021 ^ n2880 ^ n2747 ;
  assign n3042 = n2995 ^ n2982 ^ n261 ;
  assign n3043 = n2995 ^ n2950 ^ n1416 ;
  assign n3044 = n2995 & n3042 ;
  assign n3045 = n2995 ^ n2951 ^ n1318 ;
  assign n3046 = n2986 ^ n134 ^ 1'b0 ;
  assign n3047 = n2995 ^ n2962 ^ n716 ;
  assign n3048 = n2995 ^ n2953 ^ n1220 ;
  assign n3049 = n2980 ^ n345 ^ 1'b0 ;
  assign n3050 = n3044 ^ n2877 ^ n2754 ;
  assign n3051 = ( ~n2842 & n2989 ) | ( ~n2842 & n2995 ) | ( n2989 & n2995 ) ;
  assign n3052 = n2995 & n3049 ;
  assign n3053 = ( ~n2987 & n2989 ) | ( ~n2987 & n3051 ) | ( n2989 & n3051 ) ;
  assign n3054 = ( n2987 & n2988 ) | ( n2987 & n2995 ) | ( n2988 & n2995 ) ;
  assign n3055 = n2842 & ~n3054 ;
  assign n3056 = n3055 ^ n3054 ^ n2988 ;
  assign n3057 = n2995 ^ n2943 ^ n2269 ;
  assign n3058 = n2995 & n3048 ;
  assign n3059 = n2995 ^ n2947 ^ n1766 ;
  assign n3060 = n2957 ^ n859 ^ 1'b0 ;
  assign n3061 = n2995 & n3060 ;
  assign n3062 = n3061 ^ n2995 ^ n2918 ;
  assign n3063 = n2842 & ~n2995 ;
  assign n3064 = n3058 ^ n2853 ^ n2745 ;
  assign n3065 = n2995 & n3043 ;
  assign n3066 = n2995 ^ n2942 ^ n2404 ;
  assign n3067 = n3065 ^ n2905 ^ n2700 ;
  assign n3068 = n2995 & n3046 ;
  assign n3069 = n3052 ^ n2995 ^ n2872 ;
  assign n3070 = n2995 & n3045 ;
  assign n3071 = n2995 ^ n2949 ^ n1534 ;
  assign n3072 = n2995 & n3071 ;
  assign n3073 = n3070 ^ n2850 ^ n2742 ;
  assign n3074 = n2995 ^ n2967 ^ n572 ;
  assign n3075 = n3072 ^ n2902 ^ n2719 ;
  assign n3076 = n2995 & n3047 ;
  assign n3077 = n3076 ^ n2920 ^ n2776 ;
  assign n3078 = n2995 & n3074 ;
  assign n3079 = n2984 ^ n179 ^ 1'b0 ;
  assign n3080 = n3078 ^ n2926 ^ n2712 ;
  assign n3081 = n2995 & n3079 ;
  assign n3082 = n2995 & n3059 ;
  assign n3083 = n2995 & n3057 ;
  assign n3084 = n3083 ^ n2890 ^ n2793 ;
  assign n3085 = n3081 ^ n2995 ^ n2884 ;
  assign n3086 = n2995 ^ n2941 ^ n2544 ;
  assign n3087 = n3068 ^ n2995 ^ n2887 ;
  assign n3088 = n3082 ^ n2899 ^ n2758 ;
  assign n3089 = n2995 & n3066 ;
  assign n3090 = n3089 ^ n2847 ^ n2782 ;
  assign n3091 = n3012 ^ x86 ^ 1'b0 ;
  assign n3092 = x84 & n2995 ;
  assign n3093 = x81 | x82 ;
  assign n3094 = x84 | n3093 ;
  assign n3095 = ( n2839 & n3092 ) | ( n2839 & ~n3094 ) | ( n3092 & ~n3094 ) ;
  assign n3096 = n3092 ^ n2995 ^ x85 ;
  assign n3097 = ( x84 & ~n2837 ) | ( x84 & n3093 ) | ( ~n2837 & n3093 ) ;
  assign n3098 = ( ~n2839 & n3092 ) | ( ~n2839 & n3097 ) | ( n3092 & n3097 ) ;
  assign n3099 = ~n3092 & n3098 ;
  assign n3100 = n3096 | n3099 ;
  assign n3101 = ~n3095 & n3100 ;
  assign n3102 = ( ~n2690 & n3091 ) | ( ~n2690 & n3101 ) | ( n3091 & n3101 ) ;
  assign n3103 = ( ~n2544 & n3003 ) | ( ~n2544 & n3102 ) | ( n3003 & n3102 ) ;
  assign n3104 = n2995 & n3086 ;
  assign n3105 = n3104 ^ n2845 ^ x88 ;
  assign n3106 = ( ~n2404 & n3103 ) | ( ~n2404 & n3105 ) | ( n3103 & n3105 ) ;
  assign n3107 = ( ~n2269 & n3090 ) | ( ~n2269 & n3106 ) | ( n3090 & n3106 ) ;
  assign n3108 = ( ~n2139 & n3084 ) | ( ~n2139 & n3107 ) | ( n3084 & n3107 ) ;
  assign n3109 = ( ~n2009 & n3033 ) | ( ~n2009 & n3108 ) | ( n3033 & n3108 ) ;
  assign n3110 = ( ~n1885 & n3039 ) | ( ~n1885 & n3109 ) | ( n3039 & n3109 ) ;
  assign n3111 = ( ~n1766 & n3030 ) | ( ~n1766 & n3110 ) | ( n3030 & n3110 ) ;
  assign n3112 = ( ~n1652 & n3088 ) | ( ~n1652 & n3111 ) | ( n3088 & n3111 ) ;
  assign n3113 = ( ~n1534 & n3037 ) | ( ~n1534 & n3112 ) | ( n3037 & n3112 ) ;
  assign n3114 = ( ~n1416 & n3075 ) | ( ~n1416 & n3113 ) | ( n3075 & n3113 ) ;
  assign n3115 = ( ~n1318 & n3067 ) | ( ~n1318 & n3114 ) | ( n3067 & n3114 ) ;
  assign n3116 = ( ~n1220 & n3073 ) | ( ~n1220 & n3115 ) | ( n3073 & n3115 ) ;
  assign n3117 = ( ~n1118 & n3064 ) | ( ~n1118 & n3116 ) | ( n3064 & n3116 ) ;
  assign n3118 = ( ~n1034 & n3035 ) | ( ~n1034 & n3117 ) | ( n3035 & n3117 ) ;
  assign n3119 = ( ~n941 & n3031 ) | ( ~n941 & n3118 ) | ( n3031 & n3118 ) ;
  assign n3120 = ( ~n859 & n3038 ) | ( ~n859 & n3119 ) | ( n3038 & n3119 ) ;
  assign n3121 = ( ~n785 & n3062 ) | ( ~n785 & n3120 ) | ( n3062 & n3120 ) ;
  assign n3122 = ( ~n716 & n3040 ) | ( ~n716 & n3121 ) | ( n3040 & n3121 ) ;
  assign n3123 = ( ~n640 & n3077 ) | ( ~n640 & n3122 ) | ( n3077 & n3122 ) ;
  assign n3124 = ( ~n572 & n3032 ) | ( ~n572 & n3123 ) | ( n3032 & n3123 ) ;
  assign n3125 = ( ~n514 & n3080 ) | ( ~n514 & n3124 ) | ( n3080 & n3124 ) ;
  assign n3126 = ( ~n458 & n3036 ) | ( ~n458 & n3125 ) | ( n3036 & n3125 ) ;
  assign n3127 = ( ~n399 & n3027 ) | ( ~n399 & n3126 ) | ( n3027 & n3126 ) ;
  assign n3128 = ( ~n345 & n3034 ) | ( ~n345 & n3127 ) | ( n3034 & n3127 ) ;
  assign n3129 = ( ~n302 & n3069 ) | ( ~n302 & n3128 ) | ( n3069 & n3128 ) ;
  assign n3130 = ( ~n261 & n3026 ) | ( ~n261 & n3129 ) | ( n3026 & n3129 ) ;
  assign n3131 = ( ~n217 & n3050 ) | ( ~n217 & n3130 ) | ( n3050 & n3130 ) ;
  assign n3132 = ( ~n179 & n3041 ) | ( ~n179 & n3131 ) | ( n3041 & n3131 ) ;
  assign n3133 = ( ~n144 & n3085 ) | ( ~n144 & n3132 ) | ( n3085 & n3132 ) ;
  assign n3134 = ( ~n134 & n3025 ) | ( ~n134 & n3133 ) | ( n3025 & n3133 ) ;
  assign n3135 = n3087 | n3134 ;
  assign n3136 = ( ~x30 & n3053 ) | ( ~x30 & n3135 ) | ( n3053 & n3135 ) ;
  assign n3137 = ~n136 & n3136 ;
  assign n3138 = n3063 | n3137 ;
  assign n3139 = n3087 & n3134 ;
  assign n3140 = n3138 | n3139 ;
  assign n3141 = n3056 | n3140 ;
  assign n3142 = n3141 ^ n3121 ^ n716 ;
  assign n3143 = n3141 & n3142 ;
  assign n3144 = n3143 ^ n3017 ^ n2862 ;
  assign n3145 = ( x81 & n2992 ) | ( x81 & n3141 ) | ( n2992 & n3141 ) ;
  assign n3146 = n3141 ^ n3103 ^ n2404 ;
  assign n3147 = ( ~n2992 & n2993 ) | ( ~n2992 & n3145 ) | ( n2993 & n3145 ) ;
  assign n3148 = n3141 ^ n3122 ^ n640 ;
  assign n3149 = n3099 & n3141 ;
  assign n3150 = n3141 ^ n3123 ^ n572 ;
  assign n3151 = n3141 ^ n3116 ^ n1118 ;
  assign n3152 = n3141 ^ n3130 ^ n217 ;
  assign n3153 = n3141 ^ n3131 ^ n179 ;
  assign n3154 = n3141 & n3148 ;
  assign n3155 = n3141 ^ n3125 ^ n458 ;
  assign n3156 = n3154 ^ n3076 ^ n2921 ;
  assign n3157 = n3141 ^ n3129 ^ n261 ;
  assign n3158 = n3141 ^ n3111 ^ n1652 ;
  assign n3159 = n3141 & n3150 ;
  assign n3160 = n3159 ^ n3001 ^ n2924 ;
  assign n3161 = n3141 & n3155 ;
  assign n3162 = n3161 ^ n3015 ^ n2865 ;
  assign n3163 = n3141 & n3152 ;
  assign n3164 = n3163 ^ n3044 ^ n2878 ;
  assign n3165 = n3141 & n3146 ;
  assign n3166 = n3165 ^ n3104 ^ n2936 ;
  assign n3167 = n3141 & n3153 ;
  assign n3168 = n3167 ^ n3021 ^ n2881 ;
  assign n3169 = n3141 ^ n3133 ^ n134 ;
  assign n3170 = n3141 & n3157 ;
  assign n3171 = n3170 ^ n3024 ^ n2875 ;
  assign n3172 = n3141 & n3151 ;
  assign n3173 = n3172 ^ n3058 ^ n2854 ;
  assign n3174 = n3141 & n3158 ;
  assign n3175 = n3174 ^ n3082 ^ n2900 ;
  assign n3176 = n3141 & n3169 ;
  assign n3177 = n3176 ^ n3020 ^ n2930 ;
  assign n3178 = ( n3095 & n3141 ) | ( n3095 & ~n3149 ) | ( n3141 & ~n3149 ) ;
  assign n3179 = ~n3145 & n3147 ;
  assign n3180 = n3178 ^ n3096 ^ n3095 ;
  assign n3181 = n3141 ^ n3108 ^ n2009 ;
  assign n3182 = n3132 ^ n144 ^ 1'b0 ;
  assign n3183 = n3128 ^ n302 ^ 1'b0 ;
  assign n3184 = ( ~n3135 & n3139 ) | ( ~n3135 & n3141 ) | ( n3139 & n3141 ) ;
  assign n3185 = n3141 & n3183 ;
  assign n3186 = n3185 ^ n3141 ^ n3069 ;
  assign n3187 = n3141 & n3181 ;
  assign n3188 = n3141 & n3182 ;
  assign n3189 = n3112 ^ n1534 ^ 1'b0 ;
  assign n3190 = ( n136 & n3134 ) | ( n136 & n3139 ) | ( n3134 & n3139 ) ;
  assign n3191 = n3141 ^ n3119 ^ n859 ;
  assign n3192 = n3141 ^ n3113 ^ n1416 ;
  assign n3193 = n3120 ^ n785 ^ 1'b0 ;
  assign n3194 = ( n136 & n3087 ) | ( n136 & n3134 ) | ( n3087 & n3134 ) ;
  assign n3195 = ( ~n3056 & n3063 ) | ( ~n3056 & n3087 ) | ( n3063 & n3087 ) ;
  assign n3196 = n3141 ^ n3127 ^ n345 ;
  assign n3197 = n3188 ^ n3141 ^ n3085 ;
  assign n3198 = n3093 & n3141 ;
  assign n3199 = n3141 ^ n3124 ^ n514 ;
  assign n3200 = n3141 ^ n3107 ^ n2139 ;
  assign n3201 = ( n2995 & n3063 ) | ( n2995 & ~n3141 ) | ( n3063 & ~n3141 ) ;
  assign n3202 = n3141 & n3193 ;
  assign n3203 = n3102 ^ n2544 ^ 1'b0 ;
  assign n3204 = n3141 ^ n3101 ^ n2690 ;
  assign n3205 = n3141 & n3189 ;
  assign n3206 = n3141 ^ n3114 ^ n1318 ;
  assign n3207 = n3126 ^ n399 ^ 1'b0 ;
  assign n3208 = n3141 & n3207 ;
  assign n3209 = n3141 ^ n3117 ^ n1034 ;
  assign n3210 = n3187 ^ n3022 ^ n2861 ;
  assign n3211 = ( x77 & x78 ) | ( x77 & ~n3056 ) | ( x78 & ~n3056 ) ;
  assign n3212 = n3118 ^ n941 ^ 1'b0 ;
  assign n3213 = n3141 & n3206 ;
  assign n3214 = n3202 ^ n3141 ^ n3062 ;
  assign n3215 = n3141 & n3200 ;
  assign n3216 = n3141 & n3209 ;
  assign n3217 = n3141 ^ n3106 ^ n2269 ;
  assign n3218 = n3141 & n3192 ;
  assign n3219 = n3213 ^ n3065 ^ n2906 ;
  assign n3220 = n3141 & n3217 ;
  assign n3221 = ( x79 & ~n3056 ) | ( x79 & n3211 ) | ( ~n3056 & n3211 ) ;
  assign n3222 = n3056 | n3063 ;
  assign n3223 = n3110 ^ n1766 ^ 1'b0 ;
  assign n3224 = n3218 ^ n3072 ^ n2903 ;
  assign n3225 = ( ~n3139 & n3221 ) | ( ~n3139 & n3222 ) | ( n3221 & n3222 ) ;
  assign n3226 = n3141 ^ n3115 ^ n1220 ;
  assign n3227 = n3141 & n3226 ;
  assign n3228 = n3215 ^ n3083 ^ n2891 ;
  assign n3229 = n3208 ^ n3141 ^ n3027 ;
  assign n3230 = n3141 & n3212 ;
  assign n3231 = n3141 ^ n3109 ^ n1885 ;
  assign n3232 = ( n3139 & ~n3141 ) | ( n3139 & n3190 ) | ( ~n3141 & n3190 ) ;
  assign n3233 = n3141 & n3203 ;
  assign n3234 = n3233 ^ n3141 ^ n3003 ;
  assign n3235 = n3141 & n3191 ;
  assign n3236 = ~n3140 & n3195 ;
  assign n3237 = n3141 & n3204 ;
  assign n3238 = n3237 ^ n3012 ^ x86 ;
  assign n3239 = n3205 ^ n3141 ^ n3037 ;
  assign n3240 = n3141 & n3199 ;
  assign n3241 = n3141 & n3223 ;
  assign n3242 = n3241 ^ n3141 ^ n3030 ;
  assign n3243 = n3141 & n3231 ;
  assign n3244 = n3243 ^ n3009 ^ n2894 ;
  assign n3245 = ( ~n136 & n3139 ) | ( ~n136 & n3184 ) | ( n3139 & n3184 ) ;
  assign n3246 = ( n3141 & ~n3198 ) | ( n3141 & n3201 ) | ( ~n3198 & n3201 ) ;
  assign n3247 = n3227 ^ n3070 ^ n2851 ;
  assign n3248 = n3232 ^ n3194 ^ 1'b0 ;
  assign n3249 = n3240 ^ n3078 ^ n2927 ;
  assign n3250 = n3141 & n3196 ;
  assign n3251 = n3236 | n3248 ;
  assign n3252 = n3235 ^ n3006 ^ n2857 ;
  assign n3253 = n3250 ^ n3013 ^ n2870 ;
  assign n3254 = n3216 ^ n3029 ^ n2912 ;
  assign n3255 = n3230 ^ n3141 ^ n3031 ;
  assign n3256 = ~n3222 & n3225 ;
  assign n3257 = n3220 ^ n3089 ^ n2888 ;
  assign n3258 = n3246 ^ x84 ^ 1'b0 ;
  assign n3259 = x79 | x80 ;
  assign n3260 = ( x81 & n2995 ) | ( x81 & ~n3259 ) | ( n2995 & ~n3259 ) ;
  assign n3261 = ( ~x81 & n2995 ) | ( ~x81 & n3141 ) | ( n2995 & n3141 ) ;
  assign n3262 = n3260 & n3261 ;
  assign n3263 = ~x81 & n3141 ;
  assign n3264 = n3263 ^ x82 ^ 1'b0 ;
  assign n3265 = n3179 | n3264 ;
  assign n3266 = ~n3262 & n3265 ;
  assign n3267 = ( ~n2839 & n3258 ) | ( ~n2839 & n3266 ) | ( n3258 & n3266 ) ;
  assign n3268 = ( ~n2690 & n3180 ) | ( ~n2690 & n3267 ) | ( n3180 & n3267 ) ;
  assign n3269 = ( ~n2544 & n3238 ) | ( ~n2544 & n3268 ) | ( n3238 & n3268 ) ;
  assign n3270 = ( ~n2404 & n3234 ) | ( ~n2404 & n3269 ) | ( n3234 & n3269 ) ;
  assign n3271 = ( ~n2269 & n3166 ) | ( ~n2269 & n3270 ) | ( n3166 & n3270 ) ;
  assign n3272 = ( ~n2139 & n3257 ) | ( ~n2139 & n3271 ) | ( n3257 & n3271 ) ;
  assign n3273 = ( ~n2009 & n3228 ) | ( ~n2009 & n3272 ) | ( n3228 & n3272 ) ;
  assign n3274 = ( ~n1885 & n3210 ) | ( ~n1885 & n3273 ) | ( n3210 & n3273 ) ;
  assign n3275 = ( ~n1766 & n3244 ) | ( ~n1766 & n3274 ) | ( n3244 & n3274 ) ;
  assign n3276 = ( ~n1652 & n3242 ) | ( ~n1652 & n3275 ) | ( n3242 & n3275 ) ;
  assign n3277 = ( ~n1534 & n3175 ) | ( ~n1534 & n3276 ) | ( n3175 & n3276 ) ;
  assign n3278 = ( ~n1416 & n3239 ) | ( ~n1416 & n3277 ) | ( n3239 & n3277 ) ;
  assign n3279 = ( ~n1318 & n3224 ) | ( ~n1318 & n3278 ) | ( n3224 & n3278 ) ;
  assign n3280 = ( ~n1220 & n3219 ) | ( ~n1220 & n3279 ) | ( n3219 & n3279 ) ;
  assign n3281 = ( ~n1118 & n3247 ) | ( ~n1118 & n3280 ) | ( n3247 & n3280 ) ;
  assign n3282 = ( ~n1034 & n3173 ) | ( ~n1034 & n3281 ) | ( n3173 & n3281 ) ;
  assign n3283 = ( ~n941 & n3254 ) | ( ~n941 & n3282 ) | ( n3254 & n3282 ) ;
  assign n3284 = ( ~n859 & n3255 ) | ( ~n859 & n3283 ) | ( n3255 & n3283 ) ;
  assign n3285 = ( ~n785 & n3252 ) | ( ~n785 & n3284 ) | ( n3252 & n3284 ) ;
  assign n3286 = ( ~n716 & n3214 ) | ( ~n716 & n3285 ) | ( n3214 & n3285 ) ;
  assign n3287 = ( ~n640 & n3144 ) | ( ~n640 & n3286 ) | ( n3144 & n3286 ) ;
  assign n3288 = ( ~n572 & n3156 ) | ( ~n572 & n3287 ) | ( n3156 & n3287 ) ;
  assign n3289 = ( ~n514 & n3160 ) | ( ~n514 & n3288 ) | ( n3160 & n3288 ) ;
  assign n3290 = ( ~n458 & n3249 ) | ( ~n458 & n3289 ) | ( n3249 & n3289 ) ;
  assign n3291 = ( ~n399 & n3162 ) | ( ~n399 & n3290 ) | ( n3162 & n3290 ) ;
  assign n3292 = ( ~n345 & n3229 ) | ( ~n345 & n3291 ) | ( n3229 & n3291 ) ;
  assign n3293 = ( ~n302 & n3253 ) | ( ~n302 & n3292 ) | ( n3253 & n3292 ) ;
  assign n3294 = ( ~n261 & n3186 ) | ( ~n261 & n3293 ) | ( n3186 & n3293 ) ;
  assign n3295 = ( ~n217 & n3171 ) | ( ~n217 & n3294 ) | ( n3171 & n3294 ) ;
  assign n3296 = ( ~n179 & n3164 ) | ( ~n179 & n3295 ) | ( n3164 & n3295 ) ;
  assign n3297 = ( ~n144 & n3168 ) | ( ~n144 & n3296 ) | ( n3168 & n3296 ) ;
  assign n3298 = ( ~n134 & n3197 ) | ( ~n134 & n3297 ) | ( n3197 & n3297 ) ;
  assign n3299 = ( ~n136 & n3177 ) | ( ~n136 & n3298 ) | ( n3177 & n3298 ) ;
  assign n3300 = n136 & ~n3299 ;
  assign n3301 = ( n3245 & n3299 ) | ( n3245 & ~n3300 ) | ( n3299 & ~n3300 ) ;
  assign n3302 = n3251 | n3301 ;
  assign n3303 = ( n3179 & ~n3262 ) | ( n3179 & n3302 ) | ( ~n3262 & n3302 ) ;
  assign n3304 = ~n3179 & n3303 ;
  assign n3305 = n3302 ^ n3273 ^ n1885 ;
  assign n3306 = n3302 & n3305 ;
  assign n3307 = n3306 ^ n3187 ^ n3033 ;
  assign n3308 = n3302 ^ n3274 ^ n1766 ;
  assign n3309 = n3302 & n3308 ;
  assign n3310 = n3309 ^ n3243 ^ n3039 ;
  assign n3311 = n3302 ^ n3276 ^ n1534 ;
  assign n3312 = n3302 & n3311 ;
  assign n3313 = n3312 ^ n3174 ^ n3088 ;
  assign n3314 = n3302 ^ n3278 ^ n1318 ;
  assign n3315 = n3302 & n3314 ;
  assign n3316 = n3315 ^ n3218 ^ n3075 ;
  assign n3317 = n3302 ^ n3279 ^ n1220 ;
  assign n3318 = n3302 & n3317 ;
  assign n3319 = n3318 ^ n3213 ^ n3067 ;
  assign n3320 = n3302 ^ n3280 ^ n1118 ;
  assign n3321 = n3302 & n3320 ;
  assign n3322 = n3321 ^ n3227 ^ n3073 ;
  assign n3323 = n3302 ^ n3284 ^ n785 ;
  assign n3324 = n3302 & n3323 ;
  assign n3325 = n3324 ^ n3235 ^ n3038 ;
  assign n3326 = n3302 ^ n3288 ^ n514 ;
  assign n3327 = n3302 & n3326 ;
  assign n3328 = n3327 ^ n3159 ^ n3032 ;
  assign n3329 = n3302 ^ n3290 ^ n399 ;
  assign n3330 = n3302 & n3329 ;
  assign n3331 = n3330 ^ n3161 ^ n3036 ;
  assign n3332 = n3302 ^ n3294 ^ n217 ;
  assign n3333 = n3302 & n3332 ;
  assign n3334 = n3333 ^ n3170 ^ n3026 ;
  assign n3335 = n3302 ^ n3295 ^ n179 ;
  assign n3336 = n3302 & n3335 ;
  assign n3337 = n3336 ^ n3163 ^ n3050 ;
  assign n3338 = n3302 ^ n3296 ^ n144 ;
  assign n3339 = n3302 & n3338 ;
  assign n3340 = n3339 ^ n3167 ^ n3041 ;
  assign n3341 = n3297 ^ n134 ^ 1'b0 ;
  assign n3342 = n3302 & n3341 ;
  assign n3343 = n3342 ^ n3302 ^ n3197 ;
  assign n3344 = n3302 ^ n3268 ^ n2544 ;
  assign n3345 = n3302 & n3344 ;
  assign n3346 = n3345 ^ n3237 ^ n3091 ;
  assign n3347 = ( n3137 & n3141 ) | ( n3137 & ~n3251 ) | ( n3141 & ~n3251 ) ;
  assign n3348 = ~n3259 & n3302 ;
  assign n3349 = n3301 & ~n3348 ;
  assign n3350 = ( n3347 & n3348 ) | ( n3347 & ~n3349 ) | ( n3348 & ~n3349 ) ;
  assign n3351 = ( x79 & n3137 ) | ( x79 & n3302 ) | ( n3137 & n3302 ) ;
  assign n3352 = ( ~n3137 & n3256 ) | ( ~n3137 & n3351 ) | ( n3256 & n3351 ) ;
  assign n3353 = n3304 ^ n3263 ^ x82 ;
  assign n3354 = n3302 ^ n3266 ^ n2839 ;
  assign n3355 = n3302 & n3354 ;
  assign n3356 = n3355 ^ n3246 ^ x84 ;
  assign n3357 = n3267 ^ n2690 ^ 1'b0 ;
  assign n3358 = n3302 & n3357 ;
  assign n3359 = n3358 ^ n3302 ^ n3180 ;
  assign n3360 = n3269 ^ n2404 ^ 1'b0 ;
  assign n3361 = n3302 & n3360 ;
  assign n3362 = n3361 ^ n3302 ^ n3234 ;
  assign n3363 = n3302 ^ n3270 ^ n2269 ;
  assign n3364 = n3302 & n3363 ;
  assign n3365 = n3364 ^ n3165 ^ n3105 ;
  assign n3366 = n3302 ^ n3271 ^ n2139 ;
  assign n3367 = n3302 & n3366 ;
  assign n3368 = n3367 ^ n3220 ^ n3090 ;
  assign n3369 = n3302 ^ n3272 ^ n2009 ;
  assign n3370 = n3302 & n3369 ;
  assign n3371 = n3370 ^ n3215 ^ n3084 ;
  assign n3372 = n3275 ^ n1652 ^ 1'b0 ;
  assign n3373 = n3302 & n3372 ;
  assign n3374 = n3373 ^ n3302 ^ n3242 ;
  assign n3375 = n3277 ^ n1416 ^ 1'b0 ;
  assign n3376 = n3302 & n3375 ;
  assign n3377 = n3376 ^ n3302 ^ n3239 ;
  assign n3378 = n3302 ^ n3281 ^ n1034 ;
  assign n3379 = n3302 & n3378 ;
  assign n3380 = n3379 ^ n3172 ^ n3064 ;
  assign n3381 = n3302 ^ n3282 ^ n941 ;
  assign n3382 = n3302 & n3381 ;
  assign n3383 = n3382 ^ n3216 ^ n3035 ;
  assign n3384 = ~n3351 & n3352 ;
  assign n3385 = n3283 ^ n859 ^ 1'b0 ;
  assign n3386 = n3302 & n3385 ;
  assign n3387 = n3386 ^ n3302 ^ n3255 ;
  assign n3388 = n3285 ^ n716 ^ 1'b0 ;
  assign n3389 = n3302 & n3388 ;
  assign n3390 = n3389 ^ n3302 ^ n3214 ;
  assign n3391 = n3302 ^ n3286 ^ n640 ;
  assign n3392 = n3302 & n3391 ;
  assign n3393 = n3392 ^ n3143 ^ n3040 ;
  assign n3394 = n3302 ^ n3287 ^ n572 ;
  assign n3395 = n3302 & n3394 ;
  assign n3396 = n3395 ^ n3154 ^ n3077 ;
  assign n3397 = n3302 ^ n3289 ^ n458 ;
  assign n3398 = n3302 & n3397 ;
  assign n3399 = n3398 ^ n3240 ^ n3080 ;
  assign n3400 = n3291 ^ n345 ^ 1'b0 ;
  assign n3401 = n3302 & n3400 ;
  assign n3402 = n3401 ^ n3302 ^ n3229 ;
  assign n3403 = n3302 ^ n3292 ^ n302 ;
  assign n3404 = n3302 & n3403 ;
  assign n3405 = n3404 ^ n3250 ^ n3034 ;
  assign n3406 = n3293 ^ n261 ^ 1'b0 ;
  assign n3407 = n3302 & n3406 ;
  assign n3408 = n3407 ^ n3302 ^ n3186 ;
  assign n3409 = x77 | x78 ;
  assign n3410 = ( x79 & n3141 ) | ( x79 & ~n3409 ) | ( n3141 & ~n3409 ) ;
  assign n3411 = n3350 ^ x81 ^ 1'b0 ;
  assign n3412 = ( ~x79 & n3141 ) | ( ~x79 & n3302 ) | ( n3141 & n3302 ) ;
  assign n3413 = ~x79 & n3302 ;
  assign n3414 = n3410 & n3412 ;
  assign n3415 = ( ~n3177 & n3298 ) | ( ~n3177 & n3302 ) | ( n3298 & n3302 ) ;
  assign n3416 = ~n3177 & n3298 ;
  assign n3417 = n3413 ^ x80 ^ 1'b0 ;
  assign n3418 = n3384 | n3417 ;
  assign n3419 = ~n3414 & n3418 ;
  assign n3420 = ( ~n2995 & n3411 ) | ( ~n2995 & n3419 ) | ( n3411 & n3419 ) ;
  assign n3421 = ( ~n2839 & n3353 ) | ( ~n2839 & n3420 ) | ( n3353 & n3420 ) ;
  assign n3422 = ( ~n2690 & n3356 ) | ( ~n2690 & n3421 ) | ( n3356 & n3421 ) ;
  assign n3423 = ( ~n2544 & n3359 ) | ( ~n2544 & n3422 ) | ( n3359 & n3422 ) ;
  assign n3424 = ( ~n2404 & n3346 ) | ( ~n2404 & n3423 ) | ( n3346 & n3423 ) ;
  assign n3425 = ( ~n2269 & n3362 ) | ( ~n2269 & n3424 ) | ( n3362 & n3424 ) ;
  assign n3426 = ( ~n2139 & n3365 ) | ( ~n2139 & n3425 ) | ( n3365 & n3425 ) ;
  assign n3427 = ( ~n2009 & n3368 ) | ( ~n2009 & n3426 ) | ( n3368 & n3426 ) ;
  assign n3428 = ( ~n1885 & n3371 ) | ( ~n1885 & n3427 ) | ( n3371 & n3427 ) ;
  assign n3429 = ( ~n1766 & n3307 ) | ( ~n1766 & n3428 ) | ( n3307 & n3428 ) ;
  assign n3430 = ( ~n1652 & n3310 ) | ( ~n1652 & n3429 ) | ( n3310 & n3429 ) ;
  assign n3431 = ( n136 & n3177 ) | ( n136 & n3298 ) | ( n3177 & n3298 ) ;
  assign n3432 = ( n3177 & n3298 ) | ( n3177 & ~n3302 ) | ( n3298 & ~n3302 ) ;
  assign n3433 = ~n3298 & n3431 ;
  assign n3434 = ( ~n1534 & n3374 ) | ( ~n1534 & n3430 ) | ( n3374 & n3430 ) ;
  assign n3435 = ( ~n1416 & n3313 ) | ( ~n1416 & n3434 ) | ( n3313 & n3434 ) ;
  assign n3436 = ( ~n1318 & n3377 ) | ( ~n1318 & n3435 ) | ( n3377 & n3435 ) ;
  assign n3437 = ( ~n1220 & n3316 ) | ( ~n1220 & n3436 ) | ( n3316 & n3436 ) ;
  assign n3438 = ( ~n1118 & n3319 ) | ( ~n1118 & n3437 ) | ( n3319 & n3437 ) ;
  assign n3439 = ( ~n1034 & n3322 ) | ( ~n1034 & n3438 ) | ( n3322 & n3438 ) ;
  assign n3440 = ( ~n941 & n3380 ) | ( ~n941 & n3439 ) | ( n3380 & n3439 ) ;
  assign n3441 = ( ~n859 & n3383 ) | ( ~n859 & n3440 ) | ( n3383 & n3440 ) ;
  assign n3442 = ( ~n785 & n3387 ) | ( ~n785 & n3441 ) | ( n3387 & n3441 ) ;
  assign n3443 = ( ~n716 & n3325 ) | ( ~n716 & n3442 ) | ( n3325 & n3442 ) ;
  assign n3444 = ( ~n640 & n3390 ) | ( ~n640 & n3443 ) | ( n3390 & n3443 ) ;
  assign n3445 = ( n3343 & n3415 ) | ( n3343 & ~n3416 ) | ( n3415 & ~n3416 ) ;
  assign n3446 = ( ~n572 & n3393 ) | ( ~n572 & n3444 ) | ( n3393 & n3444 ) ;
  assign n3447 = ( n3431 & ~n3432 ) | ( n3431 & n3433 ) | ( ~n3432 & n3433 ) ;
  assign n3448 = ( ~n514 & n3396 ) | ( ~n514 & n3446 ) | ( n3396 & n3446 ) ;
  assign n3449 = ( ~n458 & n3328 ) | ( ~n458 & n3448 ) | ( n3328 & n3448 ) ;
  assign n3450 = ( ~n399 & n3399 ) | ( ~n399 & n3449 ) | ( n3399 & n3449 ) ;
  assign n3451 = ( ~n345 & n3331 ) | ( ~n345 & n3450 ) | ( n3331 & n3450 ) ;
  assign n3452 = ( ~n302 & n3402 ) | ( ~n302 & n3451 ) | ( n3402 & n3451 ) ;
  assign n3453 = ( ~n261 & n3405 ) | ( ~n261 & n3452 ) | ( n3405 & n3452 ) ;
  assign n3454 = ( ~n217 & n3408 ) | ( ~n217 & n3453 ) | ( n3408 & n3453 ) ;
  assign n3455 = ( ~n179 & n3334 ) | ( ~n179 & n3454 ) | ( n3334 & n3454 ) ;
  assign n3456 = ( ~n144 & n3337 ) | ( ~n144 & n3455 ) | ( n3337 & n3455 ) ;
  assign n3457 = ( ~n134 & n3340 ) | ( ~n134 & n3456 ) | ( n3340 & n3456 ) ;
  assign n3458 = n3343 & n3457 ;
  assign n3459 = ( n3177 & ~n3302 ) | ( n3177 & n3458 ) | ( ~n3302 & n3458 ) ;
  assign n3460 = ( ~x30 & n3445 ) | ( ~x30 & n3457 ) | ( n3445 & n3457 ) ;
  assign n3461 = ~n136 & n3460 ;
  assign n3462 = n3458 | n3461 ;
  assign n3463 = ( n3447 & ~n3459 ) | ( n3447 & n3462 ) | ( ~n3459 & n3462 ) ;
  assign n3464 = n3459 | n3463 ;
  assign n3465 = ( n3384 & ~n3414 ) | ( n3384 & n3464 ) | ( ~n3414 & n3464 ) ;
  assign n3466 = ~n3384 & n3465 ;
  assign n3467 = n3464 ^ n3421 ^ n2690 ;
  assign n3468 = n3464 & n3467 ;
  assign n3469 = n3468 ^ n3355 ^ n3258 ;
  assign n3470 = n3464 ^ n3425 ^ n2139 ;
  assign n3471 = n3464 & n3470 ;
  assign n3472 = n3464 ^ n3426 ^ n2009 ;
  assign n3473 = n3464 & n3472 ;
  assign n3474 = n3473 ^ n3367 ^ n3257 ;
  assign n3475 = n3464 ^ n3434 ^ n1416 ;
  assign n3476 = n3464 & n3475 ;
  assign n3477 = n3476 ^ n3312 ^ n3175 ;
  assign n3478 = n3464 ^ n3436 ^ n1220 ;
  assign n3479 = n3464 & n3478 ;
  assign n3480 = n3479 ^ n3315 ^ n3224 ;
  assign n3481 = n3464 ^ n3440 ^ n859 ;
  assign n3482 = n3464 & n3481 ;
  assign n3483 = n3482 ^ n3382 ^ n3254 ;
  assign n3484 = n3464 ^ n3442 ^ n716 ;
  assign n3485 = n3464 & n3484 ;
  assign n3486 = n3485 ^ n3324 ^ n3252 ;
  assign n3487 = n3464 ^ n3444 ^ n572 ;
  assign n3488 = n3464 & n3487 ;
  assign n3489 = n3488 ^ n3392 ^ n3144 ;
  assign n3490 = n3471 ^ n3364 ^ n3166 ;
  assign n3491 = n3464 ^ n3446 ^ n514 ;
  assign n3492 = n3464 & n3491 ;
  assign n3493 = n3492 ^ n3395 ^ n3156 ;
  assign n3494 = n3464 ^ n3449 ^ n399 ;
  assign n3495 = n3464 & n3494 ;
  assign n3496 = n3495 ^ n3398 ^ n3249 ;
  assign n3497 = n3464 ^ n3456 ^ n134 ;
  assign n3498 = n3464 & n3497 ;
  assign n3499 = n3498 ^ n3339 ^ n3168 ;
  assign n3500 = n3464 ^ n3452 ^ n261 ;
  assign n3501 = n3464 ^ n3454 ^ n179 ;
  assign n3502 = n3464 ^ n3455 ^ n144 ;
  assign n3503 = n3464 ^ n3450 ^ n345 ;
  assign n3504 = n3464 ^ n3429 ^ n1652 ;
  assign n3505 = n3435 ^ n1318 ^ 1'b0 ;
  assign n3506 = n3464 ^ n3448 ^ n458 ;
  assign n3507 = n3464 ^ n3439 ^ n941 ;
  assign n3508 = n3424 ^ n2269 ^ 1'b0 ;
  assign n3509 = n3464 ^ n3428 ^ n1766 ;
  assign n3510 = n3464 & n3509 ;
  assign n3511 = n3464 & n3500 ;
  assign n3512 = n3511 ^ n3404 ^ n3253 ;
  assign n3513 = n2995 & n3419 ;
  assign n3514 = n3451 ^ n302 ^ 1'b0 ;
  assign n3515 = n3464 & n3514 ;
  assign n3516 = n3515 ^ n3464 ^ n3402 ;
  assign n3517 = n3443 ^ n640 ^ 1'b0 ;
  assign n3518 = ( ~n2995 & n3464 ) | ( ~n2995 & n3513 ) | ( n3464 & n3513 ) ;
  assign n3519 = n3464 & n3505 ;
  assign n3520 = ( ~n3419 & n3513 ) | ( ~n3419 & n3518 ) | ( n3513 & n3518 ) ;
  assign n3521 = ~n3409 & n3464 ;
  assign n3522 = n3464 & n3507 ;
  assign n3523 = n3522 ^ n3379 ^ n3173 ;
  assign n3524 = n3441 ^ n785 ^ 1'b0 ;
  assign n3525 = n3464 & n3502 ;
  assign n3526 = n3430 ^ n1534 ^ 1'b0 ;
  assign n3527 = n3519 ^ n3464 ^ n3377 ;
  assign n3528 = n3520 ^ n3350 ^ x81 ;
  assign n3529 = n3525 ^ n3336 ^ n3164 ;
  assign n3530 = n3464 & n3504 ;
  assign n3531 = n3530 ^ n3309 ^ n3244 ;
  assign n3532 = ( n3302 & ~n3462 ) | ( n3302 & n3521 ) | ( ~n3462 & n3521 ) ;
  assign n3533 = n3422 ^ n2544 ^ 1'b0 ;
  assign n3534 = n3453 ^ n217 ^ 1'b0 ;
  assign n3535 = ( n136 & n3343 ) | ( n136 & n3457 ) | ( n3343 & n3457 ) ;
  assign n3536 = n3464 & n3517 ;
  assign n3537 = ( n3457 & n3458 ) | ( n3457 & ~n3464 ) | ( n3458 & ~n3464 ) ;
  assign n3538 = n3464 & n3533 ;
  assign n3539 = n3464 ^ n3420 ^ n2839 ;
  assign n3540 = n3464 & n3534 ;
  assign n3541 = n3464 ^ n3437 ^ n1118 ;
  assign n3542 = n3538 ^ n3464 ^ n3359 ;
  assign n3543 = n3464 & n3526 ;
  assign n3544 = n3464 & n3503 ;
  assign n3545 = n3544 ^ n3330 ^ n3162 ;
  assign n3546 = n3464 & n3524 ;
  assign n3547 = n3447 & ~n3521 ;
  assign n3548 = n3543 ^ n3464 ^ n3374 ;
  assign n3549 = n3464 & n3506 ;
  assign n3550 = n3464 ^ n3438 ^ n1034 ;
  assign n3551 = n3549 ^ n3327 ^ n3160 ;
  assign n3552 = n3464 & n3550 ;
  assign n3553 = n3464 ^ n3423 ^ n2404 ;
  assign n3554 = n3464 & n3539 ;
  assign n3555 = n3510 ^ n3306 ^ n3210 ;
  assign n3556 = n3552 ^ n3321 ^ n3247 ;
  assign n3557 = n3464 & n3553 ;
  assign n3558 = n3557 ^ n3345 ^ n3238 ;
  assign n3559 = n3466 ^ n3413 ^ x80 ;
  assign n3560 = n3464 ^ n3427 ^ n1885 ;
  assign n3561 = n3554 ^ n3304 ^ n3264 ;
  assign n3562 = n3464 & n3560 ;
  assign n3563 = n3562 ^ n3370 ^ n3228 ;
  assign n3564 = n3535 & ~n3537 ;
  assign n3565 = n3464 & n3541 ;
  assign n3566 = n3565 ^ n3318 ^ n3219 ;
  assign n3567 = n3540 ^ n3464 ^ n3408 ;
  assign n3568 = n3546 ^ n3464 ^ n3387 ;
  assign n3569 = n3464 & n3508 ;
  assign n3570 = n3464 & n3501 ;
  assign n3571 = ( n3521 & n3532 ) | ( n3521 & ~n3547 ) | ( n3532 & ~n3547 ) ;
  assign n3572 = n3570 ^ n3333 ^ n3171 ;
  assign n3573 = n3536 ^ n3464 ^ n3390 ;
  assign n3574 = n3569 ^ n3464 ^ n3362 ;
  assign n3575 = n3343 & ~n3464 ;
  assign n3576 = x75 | x76 ;
  assign n3577 = ( ~x77 & n3302 ) | ( ~x77 & n3464 ) | ( n3302 & n3464 ) ;
  assign n3578 = n3571 ^ x79 ^ 1'b0 ;
  assign n3579 = ( x77 & ~n3301 ) | ( x77 & n3576 ) | ( ~n3301 & n3576 ) ;
  assign n3580 = ( x77 & n3302 ) | ( x77 & ~n3576 ) | ( n3302 & ~n3576 ) ;
  assign n3581 = n3577 & n3580 ;
  assign n3582 = n3343 & ~n3457 ;
  assign n3583 = x77 & n3464 ;
  assign n3584 = ( ~n3302 & n3579 ) | ( ~n3302 & n3583 ) | ( n3579 & n3583 ) ;
  assign n3585 = n3583 ^ n3464 ^ x78 ;
  assign n3586 = ~n3583 & n3584 ;
  assign n3587 = n3585 | n3586 ;
  assign n3588 = ~n3581 & n3587 ;
  assign n3589 = ( ~n3141 & n3578 ) | ( ~n3141 & n3588 ) | ( n3578 & n3588 ) ;
  assign n3590 = ( ~n2995 & n3559 ) | ( ~n2995 & n3589 ) | ( n3559 & n3589 ) ;
  assign n3591 = ( ~n2839 & n3528 ) | ( ~n2839 & n3590 ) | ( n3528 & n3590 ) ;
  assign n3592 = ( ~n2690 & n3561 ) | ( ~n2690 & n3591 ) | ( n3561 & n3591 ) ;
  assign n3593 = ( ~n2544 & n3469 ) | ( ~n2544 & n3592 ) | ( n3469 & n3592 ) ;
  assign n3594 = ( ~n2404 & n3542 ) | ( ~n2404 & n3593 ) | ( n3542 & n3593 ) ;
  assign n3595 = ( ~n2269 & n3558 ) | ( ~n2269 & n3594 ) | ( n3558 & n3594 ) ;
  assign n3596 = ( ~n2139 & n3574 ) | ( ~n2139 & n3595 ) | ( n3574 & n3595 ) ;
  assign n3597 = ( ~n2009 & n3490 ) | ( ~n2009 & n3596 ) | ( n3490 & n3596 ) ;
  assign n3598 = ( ~n1885 & n3474 ) | ( ~n1885 & n3597 ) | ( n3474 & n3597 ) ;
  assign n3599 = ( ~n1766 & n3563 ) | ( ~n1766 & n3598 ) | ( n3563 & n3598 ) ;
  assign n3600 = ( ~n1652 & n3555 ) | ( ~n1652 & n3599 ) | ( n3555 & n3599 ) ;
  assign n3601 = ( ~n1534 & n3531 ) | ( ~n1534 & n3600 ) | ( n3531 & n3600 ) ;
  assign n3602 = ( ~n1416 & n3548 ) | ( ~n1416 & n3601 ) | ( n3548 & n3601 ) ;
  assign n3603 = ( n3343 & ~n3457 ) | ( n3343 & n3464 ) | ( ~n3457 & n3464 ) ;
  assign n3604 = ( ~n1318 & n3477 ) | ( ~n1318 & n3602 ) | ( n3477 & n3602 ) ;
  assign n3605 = ( ~n1220 & n3527 ) | ( ~n1220 & n3604 ) | ( n3527 & n3604 ) ;
  assign n3606 = ( ~n1118 & n3480 ) | ( ~n1118 & n3605 ) | ( n3480 & n3605 ) ;
  assign n3607 = ( ~n1034 & n3566 ) | ( ~n1034 & n3606 ) | ( n3566 & n3606 ) ;
  assign n3608 = ( ~n941 & n3556 ) | ( ~n941 & n3607 ) | ( n3556 & n3607 ) ;
  assign n3609 = ( ~n859 & n3523 ) | ( ~n859 & n3608 ) | ( n3523 & n3608 ) ;
  assign n3610 = ( ~n785 & n3483 ) | ( ~n785 & n3609 ) | ( n3483 & n3609 ) ;
  assign n3611 = ( ~n716 & n3568 ) | ( ~n716 & n3610 ) | ( n3568 & n3610 ) ;
  assign n3612 = ( ~n640 & n3486 ) | ( ~n640 & n3611 ) | ( n3486 & n3611 ) ;
  assign n3613 = n3581 | n3586 ;
  assign n3614 = ( ~n572 & n3573 ) | ( ~n572 & n3612 ) | ( n3573 & n3612 ) ;
  assign n3615 = ( ~n514 & n3489 ) | ( ~n514 & n3614 ) | ( n3489 & n3614 ) ;
  assign n3616 = ( n3499 & ~n3582 ) | ( n3499 & n3603 ) | ( ~n3582 & n3603 ) ;
  assign n3617 = ( ~n458 & n3493 ) | ( ~n458 & n3615 ) | ( n3493 & n3615 ) ;
  assign n3618 = ( ~n399 & n3551 ) | ( ~n399 & n3617 ) | ( n3551 & n3617 ) ;
  assign n3619 = ( ~n345 & n3496 ) | ( ~n345 & n3618 ) | ( n3496 & n3618 ) ;
  assign n3620 = ( ~n302 & n3545 ) | ( ~n302 & n3619 ) | ( n3545 & n3619 ) ;
  assign n3621 = ( ~n261 & n3516 ) | ( ~n261 & n3620 ) | ( n3516 & n3620 ) ;
  assign n3622 = ( ~n217 & n3512 ) | ( ~n217 & n3621 ) | ( n3512 & n3621 ) ;
  assign n3623 = ( ~n179 & n3567 ) | ( ~n179 & n3622 ) | ( n3567 & n3622 ) ;
  assign n3624 = ( ~n144 & n3572 ) | ( ~n144 & n3623 ) | ( n3572 & n3623 ) ;
  assign n3625 = ( ~n134 & n3529 ) | ( ~n134 & n3624 ) | ( n3529 & n3624 ) ;
  assign n3626 = ( ~x30 & n3616 ) | ( ~x30 & n3625 ) | ( n3616 & n3625 ) ;
  assign n3627 = ~n136 & n3626 ;
  assign n3628 = n3499 & n3625 ;
  assign n3629 = n3564 | n3628 ;
  assign n3630 = n3627 | n3629 ;
  assign n3631 = n3575 | n3630 ;
  assign n3632 = n3613 & n3631 ;
  assign n3633 = n3632 ^ n3631 ^ n3585 ;
  assign n3634 = n3631 ^ n3591 ^ n2690 ;
  assign n3635 = n3631 & n3634 ;
  assign n3636 = n3635 ^ n3554 ^ n3353 ;
  assign n3637 = n3631 ^ n3592 ^ n2544 ;
  assign n3638 = n3631 & n3637 ;
  assign n3639 = n3638 ^ n3468 ^ n3356 ;
  assign n3640 = n3631 ^ n3594 ^ n2269 ;
  assign n3641 = n3631 ^ n3596 ^ n2009 ;
  assign n3642 = n3631 & n3641 ;
  assign n3643 = n3642 ^ n3471 ^ n3365 ;
  assign n3644 = n3631 ^ n3608 ^ n859 ;
  assign n3645 = n3631 & n3644 ;
  assign n3646 = n3645 ^ n3522 ^ n3380 ;
  assign n3647 = n3631 & n3640 ;
  assign n3648 = n3647 ^ n3557 ^ n3346 ;
  assign n3649 = n3631 ^ n3609 ^ n785 ;
  assign n3650 = n3631 & n3649 ;
  assign n3651 = n3650 ^ n3482 ^ n3383 ;
  assign n3652 = n3631 ^ n3611 ^ n640 ;
  assign n3653 = n3631 & n3652 ;
  assign n3654 = n3653 ^ n3485 ^ n3325 ;
  assign n3655 = n3631 ^ n3614 ^ n514 ;
  assign n3656 = n3631 & n3655 ;
  assign n3657 = n3656 ^ n3488 ^ n3393 ;
  assign n3658 = n3631 ^ n3615 ^ n458 ;
  assign n3659 = n3631 & n3658 ;
  assign n3660 = n3659 ^ n3492 ^ n3396 ;
  assign n3661 = n3631 ^ n3618 ^ n345 ;
  assign n3662 = n3631 & n3661 ;
  assign n3663 = n3662 ^ n3495 ^ n3399 ;
  assign n3664 = n3631 ^ n3619 ^ n302 ;
  assign n3665 = n3631 & n3664 ;
  assign n3666 = n3665 ^ n3544 ^ n3331 ;
  assign n3667 = n3631 ^ n3624 ^ n134 ;
  assign n3668 = n3631 & n3667 ;
  assign n3669 = n3668 ^ n3525 ^ n3337 ;
  assign n3670 = n3610 ^ n716 ^ 1'b0 ;
  assign n3671 = n3631 & n3670 ;
  assign n3672 = n3671 ^ n3631 ^ n3568 ;
  assign n3673 = ( x70 & x71 ) | ( x70 & ~n3575 ) | ( x71 & ~n3575 ) ;
  assign n3674 = ( x73 & ~n3575 ) | ( x73 & n3673 ) | ( ~n3575 & n3673 ) ;
  assign n3675 = n3631 ^ n3605 ^ n1118 ;
  assign n3676 = n3631 ^ n3607 ^ n941 ;
  assign n3677 = n3631 & n3675 ;
  assign n3678 = n3677 ^ n3479 ^ n3316 ;
  assign n3679 = n3604 ^ n1220 ^ 1'b0 ;
  assign n3680 = n3575 | n3628 ;
  assign n3681 = ( ~n3564 & n3674 ) | ( ~n3564 & n3680 ) | ( n3674 & n3680 ) ;
  assign n3682 = n3631 ^ n3597 ^ n1885 ;
  assign n3683 = ~n3680 & n3681 ;
  assign n3684 = n3631 & n3676 ;
  assign n3685 = n3631 ^ n3623 ^ n144 ;
  assign n3686 = n3631 & n3685 ;
  assign n3687 = n3686 ^ n3570 ^ n3334 ;
  assign n3688 = n3595 ^ n2139 ^ 1'b0 ;
  assign n3689 = n3631 & n3688 ;
  assign n3690 = n3689 ^ n3631 ^ n3574 ;
  assign n3691 = n3631 ^ n3602 ^ n1318 ;
  assign n3692 = n3631 ^ n3590 ^ n2839 ;
  assign n3693 = n3631 ^ n3617 ^ n399 ;
  assign n3694 = ( ~n3499 & n3625 ) | ( ~n3499 & n3631 ) | ( n3625 & n3631 ) ;
  assign n3695 = ~n3499 & n3625 ;
  assign n3696 = ( n3669 & n3694 ) | ( n3669 & ~n3695 ) | ( n3694 & ~n3695 ) ;
  assign n3697 = n3631 & n3691 ;
  assign n3698 = n3697 ^ n3476 ^ n3313 ;
  assign n3699 = n3631 ^ n3606 ^ n1034 ;
  assign n3700 = n3612 ^ n572 ^ 1'b0 ;
  assign n3701 = n3622 ^ n179 ^ 1'b0 ;
  assign n3702 = n3631 & n3692 ;
  assign n3703 = n3631 & n3682 ;
  assign n3704 = n3703 ^ n3473 ^ n3368 ;
  assign n3705 = n3631 & n3700 ;
  assign n3706 = n3702 ^ n3520 ^ n3411 ;
  assign n3707 = n3631 ^ n3599 ^ n1652 ;
  assign n3708 = n3631 & n3699 ;
  assign n3709 = ( n3499 & n3564 ) | ( n3499 & ~n3575 ) | ( n3564 & ~n3575 ) ;
  assign n3710 = n3631 & n3707 ;
  assign n3711 = n3620 ^ n261 ^ 1'b0 ;
  assign n3712 = n3601 ^ n1416 ^ 1'b0 ;
  assign n3713 = n3631 & n3712 ;
  assign n3714 = n3631 ^ n3621 ^ n217 ;
  assign n3715 = n3710 ^ n3510 ^ n3307 ;
  assign n3716 = n3684 ^ n3552 ^ n3322 ;
  assign n3717 = n3631 & n3693 ;
  assign n3718 = n3631 & n3714 ;
  assign n3719 = n3705 ^ n3631 ^ n3573 ;
  assign n3720 = n3717 ^ n3549 ^ n3328 ;
  assign n3721 = n3631 & n3711 ;
  assign n3722 = n3721 ^ n3631 ^ n3516 ;
  assign n3723 = n3464 & ~n3630 ;
  assign n3724 = n3708 ^ n3565 ^ n3319 ;
  assign n3725 = n3713 ^ n3631 ^ n3548 ;
  assign n3726 = ~n3576 & n3631 ;
  assign n3727 = n3723 | n3726 ;
  assign n3728 = ~n3630 & n3709 ;
  assign n3729 = n3631 ^ n3598 ^ n1766 ;
  assign n3730 = n3593 ^ n2404 ^ 1'b0 ;
  assign n3731 = n3631 & n3730 ;
  assign n3732 = ( n3625 & n3628 ) | ( n3625 & ~n3631 ) | ( n3628 & ~n3631 ) ;
  assign n3733 = n3631 & n3679 ;
  assign n3734 = n3733 ^ n3631 ^ n3527 ;
  assign n3735 = n3631 ^ n3600 ^ n1534 ;
  assign n3736 = n3718 ^ n3511 ^ n3405 ;
  assign n3737 = n3631 & n3735 ;
  assign n3738 = n3731 ^ n3631 ^ n3542 ;
  assign n3739 = ( n136 & n3499 ) | ( n136 & n3625 ) | ( n3499 & n3625 ) ;
  assign n3740 = n3631 & n3729 ;
  assign n3741 = n3740 ^ n3562 ^ n3371 ;
  assign n3742 = n3631 & n3701 ;
  assign n3743 = ~n3732 & n3739 ;
  assign n3744 = n3742 ^ n3631 ^ n3567 ;
  assign n3745 = n3631 ^ n3589 ^ n2995 ;
  assign n3746 = n3631 & n3745 ;
  assign n3747 = n3746 ^ n3466 ^ n3417 ;
  assign n3748 = n3737 ^ n3530 ^ n3310 ;
  assign n3749 = n3727 ^ x77 ^ 1'b0 ;
  assign n3750 = x75 & n3631 ;
  assign n3751 = x73 | x74 ;
  assign n3752 = x75 | n3751 ;
  assign n3753 = n3750 ^ n3631 ^ x76 ;
  assign n3754 = ( x75 & ~n3462 ) | ( x75 & n3751 ) | ( ~n3462 & n3751 ) ;
  assign n3755 = ( ~n3464 & n3750 ) | ( ~n3464 & n3754 ) | ( n3750 & n3754 ) ;
  assign n3756 = ~n3750 & n3755 ;
  assign n3757 = ( n3464 & n3750 ) | ( n3464 & ~n3752 ) | ( n3750 & ~n3752 ) ;
  assign n3758 = n3753 | n3756 ;
  assign n3759 = ~n3757 & n3758 ;
  assign n3760 = ( ~n3302 & n3749 ) | ( ~n3302 & n3759 ) | ( n3749 & n3759 ) ;
  assign n3761 = ( ~n3141 & n3633 ) | ( ~n3141 & n3760 ) | ( n3633 & n3760 ) ;
  assign n3762 = n3631 ^ n3588 ^ n3141 ;
  assign n3763 = n3631 & n3762 ;
  assign n3764 = n3763 ^ n3571 ^ x79 ;
  assign n3765 = ( ~n2995 & n3761 ) | ( ~n2995 & n3764 ) | ( n3761 & n3764 ) ;
  assign n3766 = ( ~n2839 & n3747 ) | ( ~n2839 & n3765 ) | ( n3747 & n3765 ) ;
  assign n3767 = ( ~n2690 & n3706 ) | ( ~n2690 & n3766 ) | ( n3706 & n3766 ) ;
  assign n3768 = ( ~n2544 & n3636 ) | ( ~n2544 & n3767 ) | ( n3636 & n3767 ) ;
  assign n3769 = ( ~n2404 & n3639 ) | ( ~n2404 & n3768 ) | ( n3639 & n3768 ) ;
  assign n3770 = ( ~n2269 & n3738 ) | ( ~n2269 & n3769 ) | ( n3738 & n3769 ) ;
  assign n3771 = ( ~n2139 & n3648 ) | ( ~n2139 & n3770 ) | ( n3648 & n3770 ) ;
  assign n3772 = ( ~n2009 & n3690 ) | ( ~n2009 & n3771 ) | ( n3690 & n3771 ) ;
  assign n3773 = ( ~n1885 & n3643 ) | ( ~n1885 & n3772 ) | ( n3643 & n3772 ) ;
  assign n3774 = ( ~n1766 & n3704 ) | ( ~n1766 & n3773 ) | ( n3704 & n3773 ) ;
  assign n3775 = ( ~n1652 & n3741 ) | ( ~n1652 & n3774 ) | ( n3741 & n3774 ) ;
  assign n3776 = ( ~n1534 & n3715 ) | ( ~n1534 & n3775 ) | ( n3715 & n3775 ) ;
  assign n3777 = ( ~n1416 & n3748 ) | ( ~n1416 & n3776 ) | ( n3748 & n3776 ) ;
  assign n3778 = ( ~n1318 & n3725 ) | ( ~n1318 & n3777 ) | ( n3725 & n3777 ) ;
  assign n3779 = ( ~n1220 & n3698 ) | ( ~n1220 & n3778 ) | ( n3698 & n3778 ) ;
  assign n3780 = ( ~n1118 & n3734 ) | ( ~n1118 & n3779 ) | ( n3734 & n3779 ) ;
  assign n3781 = ( ~n1034 & n3678 ) | ( ~n1034 & n3780 ) | ( n3678 & n3780 ) ;
  assign n3782 = ( ~n941 & n3724 ) | ( ~n941 & n3781 ) | ( n3724 & n3781 ) ;
  assign n3783 = ( ~n859 & n3716 ) | ( ~n859 & n3782 ) | ( n3716 & n3782 ) ;
  assign n3784 = ( ~n785 & n3646 ) | ( ~n785 & n3783 ) | ( n3646 & n3783 ) ;
  assign n3785 = ( ~n716 & n3651 ) | ( ~n716 & n3784 ) | ( n3651 & n3784 ) ;
  assign n3786 = n3756 | n3757 ;
  assign n3787 = ( ~n640 & n3672 ) | ( ~n640 & n3785 ) | ( n3672 & n3785 ) ;
  assign n3788 = ( ~n572 & n3654 ) | ( ~n572 & n3787 ) | ( n3654 & n3787 ) ;
  assign n3789 = ( ~n514 & n3719 ) | ( ~n514 & n3788 ) | ( n3719 & n3788 ) ;
  assign n3790 = ( ~n458 & n3657 ) | ( ~n458 & n3789 ) | ( n3657 & n3789 ) ;
  assign n3791 = ( ~n399 & n3660 ) | ( ~n399 & n3790 ) | ( n3660 & n3790 ) ;
  assign n3792 = ( ~n345 & n3720 ) | ( ~n345 & n3791 ) | ( n3720 & n3791 ) ;
  assign n3793 = ( ~n302 & n3663 ) | ( ~n302 & n3792 ) | ( n3663 & n3792 ) ;
  assign n3794 = ( ~n261 & n3666 ) | ( ~n261 & n3793 ) | ( n3666 & n3793 ) ;
  assign n3795 = ( ~n217 & n3722 ) | ( ~n217 & n3794 ) | ( n3722 & n3794 ) ;
  assign n3796 = ( ~n179 & n3736 ) | ( ~n179 & n3795 ) | ( n3736 & n3795 ) ;
  assign n3797 = ( ~n144 & n3744 ) | ( ~n144 & n3796 ) | ( n3744 & n3796 ) ;
  assign n3798 = ( ~n134 & n3687 ) | ( ~n134 & n3797 ) | ( n3687 & n3797 ) ;
  assign n3799 = ( ~x30 & n3696 ) | ( ~x30 & n3798 ) | ( n3696 & n3798 ) ;
  assign n3800 = ~n136 & n3799 ;
  assign n3801 = n3669 & n3798 ;
  assign n3802 = n3728 | n3801 ;
  assign n3803 = n3800 | n3802 ;
  assign n3804 = n3743 | n3803 ;
  assign n3805 = n3804 ^ n3797 ^ n134 ;
  assign n3806 = n3804 & n3805 ;
  assign n3807 = n3806 ^ n3686 ^ n3572 ;
  assign n3808 = n3804 ^ n3761 ^ n2995 ;
  assign n3809 = n3804 & n3808 ;
  assign n3810 = n3809 ^ n3763 ^ n3578 ;
  assign n3811 = n3786 & n3804 ;
  assign n3812 = n3811 ^ n3804 ^ n3753 ;
  assign n3813 = n3804 ^ n3775 ^ n1534 ;
  assign n3814 = n3804 & n3813 ;
  assign n3815 = n3814 ^ n3710 ^ n3555 ;
  assign n3816 = n3804 ^ n3780 ^ n1034 ;
  assign n3817 = n3804 & n3816 ;
  assign n3818 = n3817 ^ n3677 ^ n3480 ;
  assign n3819 = n3804 ^ n3783 ^ n785 ;
  assign n3820 = n3804 & n3819 ;
  assign n3821 = n3820 ^ n3645 ^ n3523 ;
  assign n3822 = n3804 ^ n3784 ^ n716 ;
  assign n3823 = n3804 & n3822 ;
  assign n3824 = n3823 ^ n3650 ^ n3483 ;
  assign n3825 = n3804 ^ n3787 ^ n572 ;
  assign n3826 = n3804 & n3825 ;
  assign n3827 = n3826 ^ n3653 ^ n3486 ;
  assign n3828 = n3804 ^ n3789 ^ n458 ;
  assign n3829 = n3804 & n3828 ;
  assign n3830 = n3829 ^ n3656 ^ n3489 ;
  assign n3831 = n3804 ^ n3790 ^ n399 ;
  assign n3832 = n3804 & n3831 ;
  assign n3833 = n3832 ^ n3659 ^ n3493 ;
  assign n3834 = n3804 ^ n3791 ^ n345 ;
  assign n3835 = n3804 & n3834 ;
  assign n3836 = n3835 ^ n3717 ^ n3551 ;
  assign n3837 = n3804 ^ n3772 ^ n1885 ;
  assign n3838 = n3769 ^ n2269 ^ 1'b0 ;
  assign n3839 = n3804 ^ n3766 ^ n2690 ;
  assign n3840 = n3804 ^ n3770 ^ n2139 ;
  assign n3841 = n3804 & n3840 ;
  assign n3842 = n3804 & n3838 ;
  assign n3843 = n3804 ^ n3768 ^ n2404 ;
  assign n3844 = n3804 & n3843 ;
  assign n3845 = n3779 ^ n1118 ^ 1'b0 ;
  assign n3846 = n3771 ^ n2009 ^ 1'b0 ;
  assign n3847 = n3804 & n3846 ;
  assign n3848 = n3777 ^ n1318 ^ 1'b0 ;
  assign n3849 = n3760 ^ n3141 ^ 1'b0 ;
  assign n3850 = n3804 & n3848 ;
  assign n3851 = n3804 ^ n3765 ^ n2839 ;
  assign n3852 = n3804 ^ n3767 ^ n2544 ;
  assign n3853 = n3804 ^ n3792 ^ n302 ;
  assign n3854 = n3796 ^ n144 ^ 1'b0 ;
  assign n3855 = n3804 & n3854 ;
  assign n3856 = n3804 & n3837 ;
  assign n3857 = n3804 ^ n3773 ^ n1766 ;
  assign n3858 = n3804 ^ n3793 ^ n261 ;
  assign n3859 = n3804 & n3858 ;
  assign n3860 = n3804 ^ n3795 ^ n179 ;
  assign n3861 = n3804 & n3860 ;
  assign n3862 = n3788 ^ n514 ^ 1'b0 ;
  assign n3863 = n3804 & n3853 ;
  assign n3864 = n3804 & n3839 ;
  assign n3865 = n3804 ^ n3774 ^ n1652 ;
  assign n3866 = n3804 & n3865 ;
  assign n3867 = n3863 ^ n3662 ^ n3496 ;
  assign n3868 = ( x73 & n3627 ) | ( x73 & n3804 ) | ( n3627 & n3804 ) ;
  assign n3869 = n3804 ^ n3782 ^ n859 ;
  assign n3870 = n3804 & n3869 ;
  assign n3871 = n3785 ^ n640 ^ 1'b0 ;
  assign n3872 = n3804 & n3871 ;
  assign n3873 = ( ~n3627 & n3683 ) | ( ~n3627 & n3868 ) | ( n3683 & n3868 ) ;
  assign n3874 = n3794 ^ n217 ^ 1'b0 ;
  assign n3875 = n3804 ^ n3776 ^ n1416 ;
  assign n3876 = n3864 ^ n3702 ^ n3528 ;
  assign n3877 = n3804 ^ n3778 ^ n1220 ;
  assign n3878 = n3804 & n3852 ;
  assign n3879 = n3842 ^ n3804 ^ n3738 ;
  assign n3880 = n3859 ^ n3665 ^ n3545 ;
  assign n3881 = n3861 ^ n3718 ^ n3512 ;
  assign n3882 = n3855 ^ n3804 ^ n3744 ;
  assign n3883 = n3804 & n3862 ;
  assign n3884 = n3804 & n3857 ;
  assign n3885 = n3841 ^ n3647 ^ n3558 ;
  assign n3886 = n3804 & n3851 ;
  assign n3887 = n3886 ^ n3746 ^ n3559 ;
  assign n3888 = n3804 ^ n3781 ^ n941 ;
  assign n3889 = n3804 & n3888 ;
  assign n3890 = n3889 ^ n3708 ^ n3566 ;
  assign n3891 = n3883 ^ n3804 ^ n3719 ;
  assign n3892 = n3804 & n3874 ;
  assign n3893 = n3870 ^ n3684 ^ n3556 ;
  assign n3894 = n3892 ^ n3804 ^ n3722 ;
  assign n3895 = n3804 & n3877 ;
  assign n3896 = ~n3868 & n3873 ;
  assign n3897 = n3804 & n3849 ;
  assign n3898 = n3897 ^ n3804 ^ n3633 ;
  assign n3899 = n3878 ^ n3635 ^ n3561 ;
  assign n3900 = n3856 ^ n3642 ^ n3490 ;
  assign n3901 = n3844 ^ n3638 ^ n3469 ;
  assign n3902 = n3847 ^ n3804 ^ n3690 ;
  assign n3903 = n3804 & n3875 ;
  assign n3904 = n3903 ^ n3737 ^ n3531 ;
  assign n3905 = n3804 & n3845 ;
  assign n3906 = n3895 ^ n3697 ^ n3477 ;
  assign n3907 = n3884 ^ n3703 ^ n3474 ;
  assign n3908 = n3905 ^ n3804 ^ n3734 ;
  assign n3909 = n3866 ^ n3740 ^ n3563 ;
  assign n3910 = n3850 ^ n3804 ^ n3725 ;
  assign n3911 = ( n3798 & n3801 ) | ( n3798 & ~n3804 ) | ( n3801 & ~n3804 ) ;
  assign n3912 = ( x68 & x69 ) | ( x68 & ~n3743 ) | ( x69 & ~n3743 ) ;
  assign n3913 = ( ~x73 & n3631 ) | ( ~x73 & n3804 ) | ( n3631 & n3804 ) ;
  assign n3914 = n3743 | n3801 ;
  assign n3915 = ~n3751 & n3804 ;
  assign n3916 = n3803 & ~n3915 ;
  assign n3917 = ~n3669 & n3798 ;
  assign n3918 = x70 | x71 ;
  assign n3919 = ( x73 & n3631 ) | ( x73 & ~n3918 ) | ( n3631 & ~n3918 ) ;
  assign n3920 = n3913 & n3919 ;
  assign n3921 = ~x73 & n3804 ;
  assign n3922 = n3921 ^ x74 ^ 1'b0 ;
  assign n3923 = ( n3631 & n3728 ) | ( n3631 & ~n3743 ) | ( n3728 & ~n3743 ) ;
  assign n3924 = ( n3915 & ~n3916 ) | ( n3915 & n3923 ) | ( ~n3916 & n3923 ) ;
  assign n3925 = n3924 ^ x75 ^ 1'b0 ;
  assign n3926 = n3896 | n3922 ;
  assign n3927 = ~n3920 & n3926 ;
  assign n3928 = ( ~n3464 & n3925 ) | ( ~n3464 & n3927 ) | ( n3925 & n3927 ) ;
  assign n3929 = ( ~n3302 & n3812 ) | ( ~n3302 & n3928 ) | ( n3812 & n3928 ) ;
  assign n3930 = ( ~n3669 & n3798 ) | ( ~n3669 & n3804 ) | ( n3798 & n3804 ) ;
  assign n3931 = n3804 ^ n3759 ^ n3302 ;
  assign n3932 = ( x70 & ~n3743 ) | ( x70 & n3912 ) | ( ~n3743 & n3912 ) ;
  assign n3933 = n3804 & n3931 ;
  assign n3934 = n3933 ^ n3727 ^ x77 ;
  assign n3935 = ( ~n3141 & n3929 ) | ( ~n3141 & n3934 ) | ( n3929 & n3934 ) ;
  assign n3936 = ( ~n2995 & n3898 ) | ( ~n2995 & n3935 ) | ( n3898 & n3935 ) ;
  assign n3937 = ( ~n2839 & n3810 ) | ( ~n2839 & n3936 ) | ( n3810 & n3936 ) ;
  assign n3938 = ( ~n2690 & n3887 ) | ( ~n2690 & n3937 ) | ( n3887 & n3937 ) ;
  assign n3939 = ( ~n2544 & n3876 ) | ( ~n2544 & n3938 ) | ( n3876 & n3938 ) ;
  assign n3940 = ( ~n2404 & n3899 ) | ( ~n2404 & n3939 ) | ( n3899 & n3939 ) ;
  assign n3941 = ( ~n3728 & n3914 ) | ( ~n3728 & n3932 ) | ( n3914 & n3932 ) ;
  assign n3942 = ( ~n2269 & n3901 ) | ( ~n2269 & n3940 ) | ( n3901 & n3940 ) ;
  assign n3943 = ( ~n2139 & n3879 ) | ( ~n2139 & n3942 ) | ( n3879 & n3942 ) ;
  assign n3944 = ( ~n2009 & n3885 ) | ( ~n2009 & n3943 ) | ( n3885 & n3943 ) ;
  assign n3945 = ( ~n1885 & n3902 ) | ( ~n1885 & n3944 ) | ( n3902 & n3944 ) ;
  assign n3946 = ( ~n1766 & n3900 ) | ( ~n1766 & n3945 ) | ( n3900 & n3945 ) ;
  assign n3947 = ( ~n1652 & n3907 ) | ( ~n1652 & n3946 ) | ( n3907 & n3946 ) ;
  assign n3948 = ( ~n1534 & n3909 ) | ( ~n1534 & n3947 ) | ( n3909 & n3947 ) ;
  assign n3949 = ( ~n1416 & n3815 ) | ( ~n1416 & n3948 ) | ( n3815 & n3948 ) ;
  assign n3950 = ( ~n1318 & n3904 ) | ( ~n1318 & n3949 ) | ( n3904 & n3949 ) ;
  assign n3951 = ( ~n1220 & n3910 ) | ( ~n1220 & n3950 ) | ( n3910 & n3950 ) ;
  assign n3952 = n3872 ^ n3804 ^ n3672 ;
  assign n3953 = n3944 ^ n1885 ^ 1'b0 ;
  assign n3954 = ( ~n1118 & n3906 ) | ( ~n1118 & n3951 ) | ( n3906 & n3951 ) ;
  assign n3955 = ( ~n1034 & n3908 ) | ( ~n1034 & n3954 ) | ( n3908 & n3954 ) ;
  assign n3956 = ( ~n941 & n3818 ) | ( ~n941 & n3955 ) | ( n3818 & n3955 ) ;
  assign n3957 = ( n3669 & n3728 ) | ( n3669 & ~n3743 ) | ( n3728 & ~n3743 ) ;
  assign n3958 = ~n3803 & n3957 ;
  assign n3959 = ( ~n859 & n3890 ) | ( ~n859 & n3956 ) | ( n3890 & n3956 ) ;
  assign n3960 = n3950 ^ n1220 ^ 1'b0 ;
  assign n3961 = n3954 ^ n1034 ^ 1'b0 ;
  assign n3962 = ~n3914 & n3941 ;
  assign n3963 = ( n3807 & ~n3917 ) | ( n3807 & n3930 ) | ( ~n3917 & n3930 ) ;
  assign n3964 = ( ~n785 & n3893 ) | ( ~n785 & n3959 ) | ( n3893 & n3959 ) ;
  assign n3965 = ( ~n716 & n3821 ) | ( ~n716 & n3964 ) | ( n3821 & n3964 ) ;
  assign n3966 = n3928 ^ n3302 ^ 1'b0 ;
  assign n3967 = ( n136 & n3669 ) | ( n136 & n3798 ) | ( n3669 & n3798 ) ;
  assign n3968 = ( ~n640 & n3824 ) | ( ~n640 & n3965 ) | ( n3824 & n3965 ) ;
  assign n3969 = ( ~n572 & n3952 ) | ( ~n572 & n3968 ) | ( n3952 & n3968 ) ;
  assign n3970 = ~n3911 & n3967 ;
  assign n3971 = ( ~n514 & n3827 ) | ( ~n514 & n3969 ) | ( n3827 & n3969 ) ;
  assign n3972 = ( ~n458 & n3891 ) | ( ~n458 & n3971 ) | ( n3891 & n3971 ) ;
  assign n3973 = ( ~n399 & n3830 ) | ( ~n399 & n3972 ) | ( n3830 & n3972 ) ;
  assign n3974 = ( ~n345 & n3833 ) | ( ~n345 & n3973 ) | ( n3833 & n3973 ) ;
  assign n3975 = ( ~n302 & n3836 ) | ( ~n302 & n3974 ) | ( n3836 & n3974 ) ;
  assign n3976 = ( ~n261 & n3867 ) | ( ~n261 & n3975 ) | ( n3867 & n3975 ) ;
  assign n3977 = ( ~n217 & n3880 ) | ( ~n217 & n3976 ) | ( n3880 & n3976 ) ;
  assign n3978 = ( ~n179 & n3894 ) | ( ~n179 & n3977 ) | ( n3894 & n3977 ) ;
  assign n3979 = ( ~n144 & n3881 ) | ( ~n144 & n3978 ) | ( n3881 & n3978 ) ;
  assign n3980 = ( ~n134 & n3882 ) | ( ~n134 & n3979 ) | ( n3882 & n3979 ) ;
  assign n3981 = n3807 & n3980 ;
  assign n3982 = ( ~x30 & n3963 ) | ( ~x30 & n3980 ) | ( n3963 & n3980 ) ;
  assign n3983 = ~n136 & n3982 ;
  assign n3984 = n3981 | n3983 ;
  assign n3985 = n3970 | n3984 ;
  assign n3986 = n3958 | n3985 ;
  assign n3987 = ~n3918 & n3986 ;
  assign n3988 = ( n3958 & n3970 ) | ( n3958 & ~n3987 ) | ( n3970 & ~n3987 ) ;
  assign n3989 = ( n3896 & ~n3920 ) | ( n3896 & n3986 ) | ( ~n3920 & n3986 ) ;
  assign n3990 = ~n3896 & n3989 ;
  assign n3991 = n3966 & n3986 ;
  assign n3992 = n3991 ^ n3986 ^ n3812 ;
  assign n3993 = n3986 ^ n3937 ^ n2690 ;
  assign n3994 = n3986 ^ n3939 ^ n2404 ;
  assign n3995 = n3986 & n3994 ;
  assign n3996 = n3995 ^ n3878 ^ n3636 ;
  assign n3997 = n3986 ^ n3940 ^ n2269 ;
  assign n3998 = n3986 & n3997 ;
  assign n3999 = n3998 ^ n3844 ^ n3639 ;
  assign n4000 = n3953 & n3986 ;
  assign n4001 = n4000 ^ n3986 ^ n3902 ;
  assign n4002 = n3986 ^ n3945 ^ n1766 ;
  assign n4003 = n3986 & n4002 ;
  assign n4004 = n4003 ^ n3856 ^ n3643 ;
  assign n4005 = n3986 ^ n3946 ^ n1652 ;
  assign n4006 = n3986 & n4005 ;
  assign n4007 = n4006 ^ n3884 ^ n3704 ;
  assign n4008 = n3986 ^ n3947 ^ n1534 ;
  assign n4009 = n3986 & n4008 ;
  assign n4010 = n4009 ^ n3866 ^ n3741 ;
  assign n4011 = n3986 ^ n3949 ^ n1318 ;
  assign n4012 = n3986 & n4011 ;
  assign n4013 = n4012 ^ n3903 ^ n3748 ;
  assign n4014 = n3960 & n3986 ;
  assign n4015 = n4014 ^ n3986 ^ n3910 ;
  assign n4016 = n3986 ^ n3951 ^ n1118 ;
  assign n4017 = n3986 & n4016 ;
  assign n4018 = n4017 ^ n3895 ^ n3698 ;
  assign n4019 = n3961 & n3986 ;
  assign n4020 = n4019 ^ n3986 ^ n3908 ;
  assign n4021 = n3986 ^ n3964 ^ n716 ;
  assign n4022 = n3986 & n4021 ;
  assign n4023 = n4022 ^ n3820 ^ n3646 ;
  assign n4024 = n3986 ^ n3969 ^ n514 ;
  assign n4025 = n3986 & n4024 ;
  assign n4026 = n4025 ^ n3826 ^ n3654 ;
  assign n4027 = n3971 ^ n458 ^ 1'b0 ;
  assign n4028 = n3986 & n4027 ;
  assign n4029 = n4028 ^ n3986 ^ n3891 ;
  assign n4030 = n3986 ^ n3973 ^ n345 ;
  assign n4031 = n3986 & n4030 ;
  assign n4032 = n4031 ^ n3832 ^ n3660 ;
  assign n4033 = n3986 ^ n3975 ^ n261 ;
  assign n4034 = n3986 & n4033 ;
  assign n4035 = n4034 ^ n3863 ^ n3663 ;
  assign n4036 = n3977 ^ n179 ^ 1'b0 ;
  assign n4037 = n3986 & n4036 ;
  assign n4038 = n4037 ^ n3986 ^ n3894 ;
  assign n4039 = n3986 ^ n3978 ^ n144 ;
  assign n4040 = n3986 & n4039 ;
  assign n4041 = n4040 ^ n3861 ^ n3736 ;
  assign n4042 = n3979 ^ n134 ^ 1'b0 ;
  assign n4043 = n3986 & n4042 ;
  assign n4044 = n4043 ^ n3986 ^ n3882 ;
  assign n4045 = n3986 ^ n3948 ^ n1416 ;
  assign n4046 = n3986 & n4045 ;
  assign n4047 = n3986 ^ n3938 ^ n2544 ;
  assign n4048 = n4046 ^ n3814 ^ n3715 ;
  assign n4049 = ( n136 & n3807 ) | ( n136 & n3980 ) | ( n3807 & n3980 ) ;
  assign n4050 = n3986 ^ n3955 ^ n941 ;
  assign n4051 = n3986 ^ n3976 ^ n217 ;
  assign n4052 = n3986 & n3993 ;
  assign n4053 = n4052 ^ n3886 ^ n3747 ;
  assign n4054 = n3804 & ~n3984 ;
  assign n4055 = n3987 | n4054 ;
  assign n4056 = n3986 ^ n3974 ^ n302 ;
  assign n4057 = n3986 ^ n3929 ^ n3141 ;
  assign n4058 = n3942 ^ n2139 ^ 1'b0 ;
  assign n4059 = n3986 ^ n3936 ^ n2839 ;
  assign n4060 = n3968 ^ n572 ^ 1'b0 ;
  assign n4061 = n3986 ^ n3972 ^ n399 ;
  assign n4062 = n3935 ^ n2995 ^ 1'b0 ;
  assign n4063 = n3986 ^ n3943 ^ n2009 ;
  assign n4064 = ( n3980 & n3981 ) | ( n3980 & ~n3986 ) | ( n3981 & ~n3986 ) ;
  assign n4065 = n3986 ^ n3965 ^ n640 ;
  assign n4066 = n3986 ^ n3959 ^ n785 ;
  assign n4067 = n3986 & n4047 ;
  assign n4068 = n4067 ^ n3864 ^ n3706 ;
  assign n4069 = n3990 ^ n3921 ^ x74 ;
  assign n4070 = n3986 ^ n3956 ^ n859 ;
  assign n4071 = n3986 & n4070 ;
  assign n4072 = n3986 & n4058 ;
  assign n4073 = n4071 ^ n3889 ^ n3724 ;
  assign n4074 = ( n3987 & ~n3988 ) | ( n3987 & n4055 ) | ( ~n3988 & n4055 ) ;
  assign n4075 = n3986 & n4065 ;
  assign n4076 = n3986 & n4061 ;
  assign n4077 = n4075 ^ n3823 ^ n3651 ;
  assign n4078 = n4076 ^ n3829 ^ n3657 ;
  assign n4079 = ( x70 & n3800 ) | ( x70 & n3986 ) | ( n3800 & n3986 ) ;
  assign n4080 = n3986 & n4057 ;
  assign n4081 = n4080 ^ n3933 ^ n3749 ;
  assign n4082 = n4049 & ~n4064 ;
  assign n4083 = ( ~n3800 & n3962 ) | ( ~n3800 & n4079 ) | ( n3962 & n4079 ) ;
  assign n4084 = n3986 & n4059 ;
  assign n4085 = n3986 & n4060 ;
  assign n4086 = n4085 ^ n3986 ^ n3952 ;
  assign n4087 = n3986 & n4051 ;
  assign n4088 = n3986 & n4066 ;
  assign n4089 = n3986 & n4056 ;
  assign n4090 = n4088 ^ n3870 ^ n3716 ;
  assign n4091 = n3986 & n4062 ;
  assign n4092 = n3986 ^ n3927 ^ n3464 ;
  assign n4093 = n3986 & n4092 ;
  assign n4094 = n4091 ^ n3986 ^ n3898 ;
  assign n4095 = n4089 ^ n3835 ^ n3720 ;
  assign n4096 = n4084 ^ n3809 ^ n3764 ;
  assign n4097 = n4093 ^ n3924 ^ x75 ;
  assign n4098 = n4087 ^ n3859 ^ n3666 ;
  assign n4099 = n3986 & n4063 ;
  assign n4100 = ~n4079 & n4083 ;
  assign n4101 = n3986 & n4050 ;
  assign n4102 = n4101 ^ n3817 ^ n3678 ;
  assign n4103 = n4072 ^ n3986 ^ n3879 ;
  assign n4104 = n4099 ^ n3841 ^ n3648 ;
  assign n4105 = ~x70 & n3986 ;
  assign n4106 = ( ~x70 & n3804 ) | ( ~x70 & n3986 ) | ( n3804 & n3986 ) ;
  assign n4107 = n4105 ^ x71 ^ 1'b0 ;
  assign n4108 = x68 | x69 ;
  assign n4109 = n4100 | n4107 ;
  assign n4110 = ( x70 & n3804 ) | ( x70 & ~n4108 ) | ( n3804 & ~n4108 ) ;
  assign n4111 = n4106 & n4110 ;
  assign n4112 = n4109 & ~n4111 ;
  assign n4113 = n4074 ^ x73 ^ 1'b0 ;
  assign n4114 = ( ~n3631 & n4112 ) | ( ~n3631 & n4113 ) | ( n4112 & n4113 ) ;
  assign n4115 = ( ~n3464 & n4069 ) | ( ~n3464 & n4114 ) | ( n4069 & n4114 ) ;
  assign n4116 = ( ~n3302 & n4097 ) | ( ~n3302 & n4115 ) | ( n4097 & n4115 ) ;
  assign n4117 = ( ~n3141 & n3992 ) | ( ~n3141 & n4116 ) | ( n3992 & n4116 ) ;
  assign n4118 = ( ~n2995 & n4081 ) | ( ~n2995 & n4117 ) | ( n4081 & n4117 ) ;
  assign n4119 = ( ~n2839 & n4094 ) | ( ~n2839 & n4118 ) | ( n4094 & n4118 ) ;
  assign n4120 = ( ~n2690 & n4096 ) | ( ~n2690 & n4119 ) | ( n4096 & n4119 ) ;
  assign n4121 = ( ~n2544 & n4053 ) | ( ~n2544 & n4120 ) | ( n4053 & n4120 ) ;
  assign n4122 = ( ~n2404 & n4068 ) | ( ~n2404 & n4121 ) | ( n4068 & n4121 ) ;
  assign n4123 = ( ~n2269 & n3996 ) | ( ~n2269 & n4122 ) | ( n3996 & n4122 ) ;
  assign n4124 = ( ~n2139 & n3999 ) | ( ~n2139 & n4123 ) | ( n3999 & n4123 ) ;
  assign n4125 = ( ~n2009 & n4103 ) | ( ~n2009 & n4124 ) | ( n4103 & n4124 ) ;
  assign n4126 = ( ~n1885 & n4104 ) | ( ~n1885 & n4125 ) | ( n4104 & n4125 ) ;
  assign n4127 = ( ~n1766 & n4001 ) | ( ~n1766 & n4126 ) | ( n4001 & n4126 ) ;
  assign n4128 = ( ~n1652 & n4004 ) | ( ~n1652 & n4127 ) | ( n4004 & n4127 ) ;
  assign n4129 = ( ~n1534 & n4007 ) | ( ~n1534 & n4128 ) | ( n4007 & n4128 ) ;
  assign n4130 = ( ~n1416 & n4010 ) | ( ~n1416 & n4129 ) | ( n4010 & n4129 ) ;
  assign n4131 = ( ~n1318 & n4048 ) | ( ~n1318 & n4130 ) | ( n4048 & n4130 ) ;
  assign n4132 = ( ~n1220 & n4013 ) | ( ~n1220 & n4131 ) | ( n4013 & n4131 ) ;
  assign n4133 = ( ~n1118 & n4015 ) | ( ~n1118 & n4132 ) | ( n4015 & n4132 ) ;
  assign n4134 = ( ~n1034 & n4018 ) | ( ~n1034 & n4133 ) | ( n4018 & n4133 ) ;
  assign n4135 = ( ~n941 & n4020 ) | ( ~n941 & n4134 ) | ( n4020 & n4134 ) ;
  assign n4136 = ( ~n859 & n4102 ) | ( ~n859 & n4135 ) | ( n4102 & n4135 ) ;
  assign n4137 = ( ~n785 & n4073 ) | ( ~n785 & n4136 ) | ( n4073 & n4136 ) ;
  assign n4138 = ( ~n716 & n4090 ) | ( ~n716 & n4137 ) | ( n4090 & n4137 ) ;
  assign n4139 = ( ~n640 & n4023 ) | ( ~n640 & n4138 ) | ( n4023 & n4138 ) ;
  assign n4140 = ( ~n572 & n4077 ) | ( ~n572 & n4139 ) | ( n4077 & n4139 ) ;
  assign n4141 = ( ~n514 & n4086 ) | ( ~n514 & n4140 ) | ( n4086 & n4140 ) ;
  assign n4142 = n4134 ^ n941 ^ 1'b0 ;
  assign n4143 = ( ~n458 & n4026 ) | ( ~n458 & n4141 ) | ( n4026 & n4141 ) ;
  assign n4144 = ( n3807 & ~n3980 ) | ( n3807 & n3986 ) | ( ~n3980 & n3986 ) ;
  assign n4145 = n3807 & ~n3980 ;
  assign n4146 = ( n4044 & n4144 ) | ( n4044 & ~n4145 ) | ( n4144 & ~n4145 ) ;
  assign n4147 = n4143 ^ n399 ^ 1'b0 ;
  assign n4148 = ( ~n399 & n4029 ) | ( ~n399 & n4143 ) | ( n4029 & n4143 ) ;
  assign n4149 = ( n3807 & ~n3986 ) | ( n3807 & n4082 ) | ( ~n3986 & n4082 ) ;
  assign n4150 = n4140 ^ n514 ^ 1'b0 ;
  assign n4151 = n4124 ^ n2009 ^ 1'b0 ;
  assign n4152 = n4126 ^ n1766 ^ 1'b0 ;
  assign n4153 = n4116 ^ n3141 ^ 1'b0 ;
  assign n4154 = n4118 ^ n2839 ^ 1'b0 ;
  assign n4155 = ( ~n345 & n4078 ) | ( ~n345 & n4148 ) | ( n4078 & n4148 ) ;
  assign n4156 = ( ~n302 & n4032 ) | ( ~n302 & n4155 ) | ( n4032 & n4155 ) ;
  assign n4157 = ( ~n261 & n4095 ) | ( ~n261 & n4156 ) | ( n4095 & n4156 ) ;
  assign n4158 = ( ~n217 & n4035 ) | ( ~n217 & n4157 ) | ( n4035 & n4157 ) ;
  assign n4159 = ( ~n179 & n4098 ) | ( ~n179 & n4158 ) | ( n4098 & n4158 ) ;
  assign n4160 = ( ~n144 & n4038 ) | ( ~n144 & n4159 ) | ( n4038 & n4159 ) ;
  assign n4161 = ( ~n134 & n4041 ) | ( ~n134 & n4160 ) | ( n4041 & n4160 ) ;
  assign n4162 = ( ~x30 & n4146 ) | ( ~x30 & n4161 ) | ( n4146 & n4161 ) ;
  assign n4163 = ~n136 & n4162 ;
  assign n4164 = ~n4044 & n4161 ;
  assign n4165 = ( n4161 & n4163 ) | ( n4161 & ~n4164 ) | ( n4163 & ~n4164 ) ;
  assign n4166 = n4082 | n4165 ;
  assign n4167 = n4149 | n4166 ;
  assign n4168 = n4167 ^ n4160 ^ n134 ;
  assign n4169 = n4167 & n4168 ;
  assign n4170 = n4169 ^ n4040 ^ n3881 ;
  assign n4171 = ( n4100 & ~n4111 ) | ( n4100 & n4167 ) | ( ~n4111 & n4167 ) ;
  assign n4172 = ~n4100 & n4171 ;
  assign n4173 = n4167 ^ n4114 ^ n3464 ;
  assign n4174 = n4167 & n4173 ;
  assign n4175 = n4174 ^ n3990 ^ n3922 ;
  assign n4176 = n4153 & n4167 ;
  assign n4177 = n4176 ^ n4167 ^ n3992 ;
  assign n4178 = n4167 ^ n4117 ^ n2995 ;
  assign n4179 = n4167 & n4178 ;
  assign n4180 = n4179 ^ n4080 ^ n3934 ;
  assign n4181 = n4154 & n4167 ;
  assign n4182 = n4181 ^ n4167 ^ n4094 ;
  assign n4183 = n4167 ^ n4119 ^ n2690 ;
  assign n4184 = n4167 & n4183 ;
  assign n4185 = n4184 ^ n4084 ^ n3810 ;
  assign n4186 = n4167 ^ n4120 ^ n2544 ;
  assign n4187 = n4167 & n4186 ;
  assign n4188 = n4187 ^ n4052 ^ n3887 ;
  assign n4189 = n4167 ^ n4123 ^ n2139 ;
  assign n4190 = n4167 & n4189 ;
  assign n4191 = n4190 ^ n3998 ^ n3901 ;
  assign n4192 = n4151 & n4167 ;
  assign n4193 = n4192 ^ n4167 ^ n4103 ;
  assign n4194 = n4152 & n4167 ;
  assign n4195 = n4194 ^ n4167 ^ n4001 ;
  assign n4196 = n4167 ^ n4128 ^ n1534 ;
  assign n4197 = n4167 & n4196 ;
  assign n4198 = n4197 ^ n4006 ^ n3907 ;
  assign n4199 = n4167 ^ n4130 ^ n1318 ;
  assign n4200 = n4167 & n4199 ;
  assign n4201 = n4200 ^ n4046 ^ n3815 ;
  assign n4202 = n4167 ^ n4133 ^ n1034 ;
  assign n4203 = n4167 & n4202 ;
  assign n4204 = n4203 ^ n4017 ^ n3906 ;
  assign n4205 = n4142 & n4167 ;
  assign n4206 = n4205 ^ n4167 ^ n4020 ;
  assign n4207 = n4167 ^ n4135 ^ n859 ;
  assign n4208 = n4167 & n4207 ;
  assign n4209 = n4208 ^ n4101 ^ n3818 ;
  assign n4210 = n4167 ^ n4136 ^ n785 ;
  assign n4211 = n4167 & n4210 ;
  assign n4212 = n4211 ^ n4071 ^ n3890 ;
  assign n4213 = n4167 ^ n4137 ^ n716 ;
  assign n4214 = n4167 & n4213 ;
  assign n4215 = n4214 ^ n4088 ^ n3893 ;
  assign n4216 = n4167 ^ n4139 ^ n572 ;
  assign n4217 = n4167 & n4216 ;
  assign n4218 = n4217 ^ n4075 ^ n3824 ;
  assign n4219 = n4150 & n4167 ;
  assign n4220 = n4219 ^ n4167 ^ n4086 ;
  assign n4221 = n4167 ^ n4141 ^ n458 ;
  assign n4222 = n4167 & n4221 ;
  assign n4223 = n4222 ^ n4025 ^ n3827 ;
  assign n4224 = n4147 & n4167 ;
  assign n4225 = n4224 ^ n4167 ^ n4029 ;
  assign n4226 = n4167 ^ n4148 ^ n345 ;
  assign n4227 = n4167 & n4226 ;
  assign n4228 = n4227 ^ n4076 ^ n3830 ;
  assign n4229 = n4167 ^ n4122 ^ n2269 ;
  assign n4230 = n4167 ^ n4138 ^ n640 ;
  assign n4231 = n3986 & ~n4166 ;
  assign n4232 = n4167 & n4229 ;
  assign n4233 = n4232 ^ n3995 ^ n3899 ;
  assign n4234 = ( n4044 & n4161 ) | ( n4044 & ~n4167 ) | ( n4161 & ~n4167 ) ;
  assign n4235 = n4167 ^ n4155 ^ n302 ;
  assign n4236 = n4167 ^ n4157 ^ n217 ;
  assign n4237 = n4167 & n4236 ;
  assign n4238 = n4167 ^ n4156 ^ n261 ;
  assign n4239 = n4237 ^ n4034 ^ n3867 ;
  assign n4240 = n4132 ^ n1118 ^ 1'b0 ;
  assign n4241 = n4167 ^ n4131 ^ n1220 ;
  assign n4242 = n4167 & n4240 ;
  assign n4243 = n4167 & n4241 ;
  assign n4244 = ~n4108 & n4167 ;
  assign n4245 = n4243 ^ n4012 ^ n3904 ;
  assign n4246 = n4044 & ~n4167 ;
  assign n4247 = ( x62 & x63 ) | ( x62 & ~n4246 ) | ( x63 & ~n4246 ) ;
  assign n4248 = n4159 ^ n144 ^ 1'b0 ;
  assign n4249 = n4167 ^ n4129 ^ n1416 ;
  assign n4250 = n4167 & n4235 ;
  assign n4251 = n4250 ^ n4031 ^ n3833 ;
  assign n4252 = ( n4044 & ~n4161 ) | ( n4044 & n4167 ) | ( ~n4161 & n4167 ) ;
  assign n4253 = n4167 & n4238 ;
  assign n4254 = n4253 ^ n4089 ^ n3836 ;
  assign n4255 = ( n136 & n4044 ) | ( n136 & n4161 ) | ( n4044 & n4161 ) ;
  assign n4256 = n4167 ^ n4125 ^ n1885 ;
  assign n4257 = n4167 ^ n4112 ^ n3631 ;
  assign n4258 = n4167 ^ n4127 ^ n1652 ;
  assign n4259 = n4172 ^ n4105 ^ x71 ;
  assign n4260 = n4167 & n4257 ;
  assign n4261 = n4161 ^ n4044 ^ 1'b0 ;
  assign n4262 = n4167 ^ n4158 ^ n179 ;
  assign n4263 = n4167 & n4262 ;
  assign n4264 = n4260 ^ n4074 ^ x73 ;
  assign n4265 = n4263 ^ n4087 ^ n3880 ;
  assign n4266 = n4167 ^ n4115 ^ n3302 ;
  assign n4267 = n4167 & n4230 ;
  assign n4268 = n4167 & n4266 ;
  assign n4269 = n4267 ^ n4022 ^ n3821 ;
  assign n4270 = n4242 ^ n4167 ^ n4015 ;
  assign n4271 = n4167 & n4249 ;
  assign n4272 = n4271 ^ n4009 ^ n3909 ;
  assign n4273 = ( n4161 & n4252 ) | ( n4161 & ~n4261 ) | ( n4252 & ~n4261 ) ;
  assign n4274 = ( x64 & ~n4246 ) | ( x64 & n4247 ) | ( ~n4246 & n4247 ) ;
  assign n4275 = n4167 & n4256 ;
  assign n4276 = n4275 ^ n4099 ^ n3885 ;
  assign n4277 = n4167 & n4248 ;
  assign n4278 = n4161 & n4234 ;
  assign n4279 = ( n4246 & n4255 ) | ( n4246 & ~n4278 ) | ( n4255 & ~n4278 ) ;
  assign n4280 = n4277 ^ n4167 ^ n4038 ;
  assign n4281 = ( n4163 & n4273 ) | ( n4163 & ~n4279 ) | ( n4273 & ~n4279 ) ;
  assign n4282 = n4167 ^ n4121 ^ n2404 ;
  assign n4283 = n4231 | n4244 ;
  assign n4284 = n4167 & n4282 ;
  assign n4285 = n4284 ^ n4067 ^ n3876 ;
  assign n4286 = n4167 & n4258 ;
  assign n4287 = n4286 ^ n4003 ^ n3900 ;
  assign n4288 = n4268 ^ n4093 ^ n3925 ;
  assign n4289 = n4283 ^ x70 ^ 1'b0 ;
  assign n4290 = x68 & n4167 ;
  assign n4291 = x66 | x67 ;
  assign n4292 = x68 | n4291 ;
  assign n4293 = ( n3986 & n4290 ) | ( n3986 & ~n4292 ) | ( n4290 & ~n4292 ) ;
  assign n4294 = n4290 ^ n4167 ^ x69 ;
  assign n4295 = ( x68 & ~n3984 ) | ( x68 & n4291 ) | ( ~n3984 & n4291 ) ;
  assign n4296 = ( ~n3986 & n4290 ) | ( ~n3986 & n4295 ) | ( n4290 & n4295 ) ;
  assign n4297 = ~n4290 & n4296 ;
  assign n4298 = n4294 | n4297 ;
  assign n4299 = ~n4293 & n4298 ;
  assign n4300 = ( ~n3804 & n4289 ) | ( ~n3804 & n4299 ) | ( n4289 & n4299 ) ;
  assign n4301 = ( ~n3631 & n4259 ) | ( ~n3631 & n4300 ) | ( n4259 & n4300 ) ;
  assign n4302 = ( ~n3464 & n4264 ) | ( ~n3464 & n4301 ) | ( n4264 & n4301 ) ;
  assign n4303 = ( ~n3302 & n4175 ) | ( ~n3302 & n4302 ) | ( n4175 & n4302 ) ;
  assign n4304 = ( ~n3141 & n4288 ) | ( ~n3141 & n4303 ) | ( n4288 & n4303 ) ;
  assign n4305 = ( ~n2995 & n4177 ) | ( ~n2995 & n4304 ) | ( n4177 & n4304 ) ;
  assign n4306 = ( ~n2839 & n4180 ) | ( ~n2839 & n4305 ) | ( n4180 & n4305 ) ;
  assign n4307 = ( ~n2690 & n4182 ) | ( ~n2690 & n4306 ) | ( n4182 & n4306 ) ;
  assign n4308 = ( ~n2544 & n4185 ) | ( ~n2544 & n4307 ) | ( n4185 & n4307 ) ;
  assign n4309 = ( ~n2404 & n4188 ) | ( ~n2404 & n4308 ) | ( n4188 & n4308 ) ;
  assign n4310 = ( ~n2269 & n4285 ) | ( ~n2269 & n4309 ) | ( n4285 & n4309 ) ;
  assign n4311 = n4293 | n4297 ;
  assign n4312 = ( ~n2139 & n4233 ) | ( ~n2139 & n4310 ) | ( n4233 & n4310 ) ;
  assign n4313 = ( ~n2009 & n4191 ) | ( ~n2009 & n4312 ) | ( n4191 & n4312 ) ;
  assign n4314 = ( ~n1885 & n4193 ) | ( ~n1885 & n4313 ) | ( n4193 & n4313 ) ;
  assign n4315 = ( ~n1766 & n4276 ) | ( ~n1766 & n4314 ) | ( n4276 & n4314 ) ;
  assign n4316 = ( ~n1652 & n4195 ) | ( ~n1652 & n4315 ) | ( n4195 & n4315 ) ;
  assign n4317 = ( ~n1534 & n4287 ) | ( ~n1534 & n4316 ) | ( n4287 & n4316 ) ;
  assign n4318 = ( ~n1416 & n4198 ) | ( ~n1416 & n4317 ) | ( n4198 & n4317 ) ;
  assign n4319 = ( ~n1318 & n4272 ) | ( ~n1318 & n4318 ) | ( n4272 & n4318 ) ;
  assign n4320 = ( ~n1220 & n4201 ) | ( ~n1220 & n4319 ) | ( n4201 & n4319 ) ;
  assign n4321 = ( ~n1118 & n4245 ) | ( ~n1118 & n4320 ) | ( n4245 & n4320 ) ;
  assign n4322 = ( ~n1034 & n4270 ) | ( ~n1034 & n4321 ) | ( n4270 & n4321 ) ;
  assign n4323 = ( ~n941 & n4204 ) | ( ~n941 & n4322 ) | ( n4204 & n4322 ) ;
  assign n4324 = ( ~n859 & n4206 ) | ( ~n859 & n4323 ) | ( n4206 & n4323 ) ;
  assign n4325 = ( ~n785 & n4209 ) | ( ~n785 & n4324 ) | ( n4209 & n4324 ) ;
  assign n4326 = ( ~n716 & n4212 ) | ( ~n716 & n4325 ) | ( n4212 & n4325 ) ;
  assign n4327 = ( ~n640 & n4215 ) | ( ~n640 & n4326 ) | ( n4215 & n4326 ) ;
  assign n4328 = ( ~n572 & n4269 ) | ( ~n572 & n4327 ) | ( n4269 & n4327 ) ;
  assign n4329 = ( ~n514 & n4218 ) | ( ~n514 & n4328 ) | ( n4218 & n4328 ) ;
  assign n4330 = ( ~n458 & n4220 ) | ( ~n458 & n4329 ) | ( n4220 & n4329 ) ;
  assign n4331 = ( ~n399 & n4223 ) | ( ~n399 & n4330 ) | ( n4223 & n4330 ) ;
  assign n4332 = ( ~n345 & n4225 ) | ( ~n345 & n4331 ) | ( n4225 & n4331 ) ;
  assign n4333 = ( ~n302 & n4228 ) | ( ~n302 & n4332 ) | ( n4228 & n4332 ) ;
  assign n4334 = ( ~n261 & n4251 ) | ( ~n261 & n4333 ) | ( n4251 & n4333 ) ;
  assign n4335 = ( ~n217 & n4254 ) | ( ~n217 & n4334 ) | ( n4254 & n4334 ) ;
  assign n4336 = ( ~n179 & n4239 ) | ( ~n179 & n4335 ) | ( n4239 & n4335 ) ;
  assign n4337 = ( ~n144 & n4265 ) | ( ~n144 & n4336 ) | ( n4265 & n4336 ) ;
  assign n4338 = ( ~n134 & n4280 ) | ( ~n134 & n4337 ) | ( n4280 & n4337 ) ;
  assign n4339 = n4170 & n4338 ;
  assign n4340 = ( n4274 & n4279 ) | ( n4274 & ~n4339 ) | ( n4279 & ~n4339 ) ;
  assign n4341 = ~n4279 & n4340 ;
  assign n4342 = ( ~n136 & n4170 ) | ( ~n136 & n4338 ) | ( n4170 & n4338 ) ;
  assign n4343 = n4273 | n4342 ;
  assign n4344 = ~n136 & n4343 ;
  assign n4345 = n4339 | n4344 ;
  assign n4346 = n4279 | n4345 ;
  assign n4347 = n4346 ^ n4326 ^ n640 ;
  assign n4348 = n4346 & n4347 ;
  assign n4349 = n4346 ^ n4302 ^ n3302 ;
  assign n4350 = n4346 ^ n4301 ^ n3464 ;
  assign n4351 = n4346 ^ n4324 ^ n785 ;
  assign n4352 = n4346 & n4349 ;
  assign n4353 = n4352 ^ n4174 ^ n4069 ;
  assign n4354 = n4346 ^ n4310 ^ n2139 ;
  assign n4355 = n4346 & n4354 ;
  assign n4356 = n4346 ^ n4308 ^ n2404 ;
  assign n4357 = n4346 & n4356 ;
  assign n4358 = ~n4291 & n4346 ;
  assign n4359 = n4311 & n4346 ;
  assign n4360 = n4346 ^ n4328 ^ n514 ;
  assign n4361 = n4345 & ~n4358 ;
  assign n4362 = ( n4281 & n4358 ) | ( n4281 & ~n4361 ) | ( n4358 & ~n4361 ) ;
  assign n4363 = n4357 ^ n4187 ^ n4053 ;
  assign n4364 = n4359 ^ n4346 ^ n4294 ;
  assign n4365 = n4346 ^ n4316 ^ n1534 ;
  assign n4366 = n4346 & n4365 ;
  assign n4367 = n4346 & n4360 ;
  assign n4368 = n4346 ^ n4317 ^ n1416 ;
  assign n4369 = n4346 & n4368 ;
  assign n4370 = n4346 ^ n4318 ^ n1318 ;
  assign n4371 = n4367 ^ n4217 ^ n4077 ;
  assign n4372 = n4346 & n4350 ;
  assign n4373 = n4346 & n4370 ;
  assign n4374 = n4346 & n4351 ;
  assign n4375 = n4366 ^ n4286 ^ n4004 ;
  assign n4376 = n4372 ^ n4260 ^ n4113 ;
  assign n4377 = n4374 ^ n4208 ^ n4102 ;
  assign n4378 = n4355 ^ n4232 ^ n3996 ;
  assign n4379 = n4373 ^ n4271 ^ n4010 ;
  assign n4380 = n4369 ^ n4197 ^ n4007 ;
  assign n4381 = n4348 ^ n4214 ^ n4090 ;
  assign n4382 = n4346 ^ n4314 ^ n1766 ;
  assign n4383 = n4346 ^ n4312 ^ n2009 ;
  assign n4384 = n4346 & n4383 ;
  assign n4385 = n4313 ^ n1885 ^ 1'b0 ;
  assign n4386 = n4346 & n4385 ;
  assign n4387 = n4346 & n4382 ;
  assign n4388 = n4346 ^ n4320 ^ n1118 ;
  assign n4389 = n4306 ^ n2690 ^ 1'b0 ;
  assign n4390 = n4346 & n4389 ;
  assign n4391 = n4390 ^ n4346 ^ n4182 ;
  assign n4392 = n4346 ^ n4300 ^ n3631 ;
  assign n4393 = n4346 ^ n4319 ^ n1220 ;
  assign n4394 = n4329 ^ n458 ^ 1'b0 ;
  assign n4395 = n4346 & n4392 ;
  assign n4396 = n4346 ^ n4336 ^ n144 ;
  assign n4397 = n4346 ^ n4305 ^ n2839 ;
  assign n4398 = n4337 ^ n134 ^ 1'b0 ;
  assign n4399 = n4346 & n4398 ;
  assign n4400 = n4346 & n4397 ;
  assign n4401 = n4321 ^ n1034 ^ 1'b0 ;
  assign n4402 = n4346 ^ n4309 ^ n2269 ;
  assign n4403 = n4346 & n4402 ;
  assign n4404 = n4346 & n4388 ;
  assign n4405 = n4346 & n4401 ;
  assign n4406 = n4304 ^ n2995 ^ 1'b0 ;
  assign n4407 = n4346 ^ n4303 ^ n3141 ;
  assign n4408 = n4399 ^ n4346 ^ n4280 ;
  assign n4409 = n4346 ^ n4333 ^ n261 ;
  assign n4410 = n4346 & n4407 ;
  assign n4411 = n4386 ^ n4346 ^ n4193 ;
  assign n4412 = n4346 & n4406 ;
  assign n4413 = n4412 ^ n4346 ^ n4177 ;
  assign n4414 = n4346 ^ n4335 ^ n179 ;
  assign n4415 = n4315 ^ n1652 ^ 1'b0 ;
  assign n4416 = n4346 ^ n4330 ^ n399 ;
  assign n4417 = n4346 & n4414 ;
  assign n4418 = n4404 ^ n4243 ^ n4013 ;
  assign n4419 = n4346 ^ n4334 ^ n217 ;
  assign n4420 = n4346 & n4415 ;
  assign n4421 = n4405 ^ n4346 ^ n4270 ;
  assign n4422 = n4400 ^ n4179 ^ n4081 ;
  assign n4423 = n4417 ^ n4237 ^ n4035 ;
  assign n4424 = n4346 ^ n4307 ^ n2544 ;
  assign n4425 = n4346 & n4394 ;
  assign n4426 = n4346 & n4424 ;
  assign n4427 = n4426 ^ n4184 ^ n4096 ;
  assign n4428 = n4410 ^ n4268 ^ n4097 ;
  assign n4429 = n4387 ^ n4275 ^ n4104 ;
  assign n4430 = n4384 ^ n4190 ^ n3999 ;
  assign n4431 = n4395 ^ n4172 ^ n4107 ;
  assign n4432 = n4346 ^ n4327 ^ n572 ;
  assign n4433 = n4346 ^ n4322 ^ n941 ;
  assign n4434 = n4346 & n4416 ;
  assign n4435 = n4434 ^ n4222 ^ n4026 ;
  assign n4436 = n4346 & n4433 ;
  assign n4437 = n4346 & n4393 ;
  assign n4438 = n4436 ^ n4203 ^ n4018 ;
  assign n4439 = n4346 & n4419 ;
  assign n4440 = n4439 ^ n4253 ^ n4095 ;
  assign n4441 = n4425 ^ n4346 ^ n4220 ;
  assign n4442 = n4346 ^ n4325 ^ n716 ;
  assign n4443 = n4346 & n4442 ;
  assign n4444 = n4443 ^ n4211 ^ n4073 ;
  assign n4445 = n4323 ^ n859 ^ 1'b0 ;
  assign n4446 = n4346 & n4409 ;
  assign n4447 = n4346 & n4445 ;
  assign n4448 = n4346 & n4432 ;
  assign n4449 = n4448 ^ n4267 ^ n4023 ;
  assign n4450 = n4346 & n4396 ;
  assign n4451 = n4446 ^ n4250 ^ n4032 ;
  assign n4452 = n4450 ^ n4263 ^ n4098 ;
  assign n4453 = n4447 ^ n4346 ^ n4206 ;
  assign n4454 = n4403 ^ n4284 ^ n4068 ;
  assign n4455 = n4437 ^ n4200 ^ n4048 ;
  assign n4456 = n4420 ^ n4346 ^ n4195 ;
  assign n4457 = x66 & n4346 ;
  assign n4458 = n4457 ^ n4346 ^ x67 ;
  assign n4459 = x64 | x65 ;
  assign n4460 = ( x66 & ~n4165 ) | ( x66 & n4459 ) | ( ~n4165 & n4459 ) ;
  assign n4461 = ( ~n4167 & n4457 ) | ( ~n4167 & n4460 ) | ( n4457 & n4460 ) ;
  assign n4462 = n4346 ^ n4299 ^ n3804 ;
  assign n4463 = ~n4457 & n4461 ;
  assign n4464 = n4458 | n4463 ;
  assign n4465 = n4346 & n4462 ;
  assign n4466 = n4465 ^ n4283 ^ x70 ;
  assign n4467 = x66 | n4459 ;
  assign n4468 = ( n4167 & n4457 ) | ( n4167 & ~n4467 ) | ( n4457 & ~n4467 ) ;
  assign n4469 = n4464 & ~n4468 ;
  assign n4470 = n4346 ^ n4332 ^ n302 ;
  assign n4471 = n4362 ^ x68 ^ 1'b0 ;
  assign n4472 = ( ~n3986 & n4469 ) | ( ~n3986 & n4471 ) | ( n4469 & n4471 ) ;
  assign n4473 = ( ~n3804 & n4364 ) | ( ~n3804 & n4472 ) | ( n4364 & n4472 ) ;
  assign n4474 = ( ~n3631 & n4466 ) | ( ~n3631 & n4473 ) | ( n4466 & n4473 ) ;
  assign n4475 = ( ~n3464 & n4431 ) | ( ~n3464 & n4474 ) | ( n4431 & n4474 ) ;
  assign n4476 = ( ~n3302 & n4376 ) | ( ~n3302 & n4475 ) | ( n4376 & n4475 ) ;
  assign n4477 = ( ~n3141 & n4353 ) | ( ~n3141 & n4476 ) | ( n4353 & n4476 ) ;
  assign n4478 = ( ~n2995 & n4428 ) | ( ~n2995 & n4477 ) | ( n4428 & n4477 ) ;
  assign n4479 = ( ~n2839 & n4413 ) | ( ~n2839 & n4478 ) | ( n4413 & n4478 ) ;
  assign n4480 = ( ~n2690 & n4422 ) | ( ~n2690 & n4479 ) | ( n4422 & n4479 ) ;
  assign n4481 = ( ~n2544 & n4391 ) | ( ~n2544 & n4480 ) | ( n4391 & n4480 ) ;
  assign n4482 = ( ~n2404 & n4427 ) | ( ~n2404 & n4481 ) | ( n4427 & n4481 ) ;
  assign n4483 = n4480 ^ n2544 ^ 1'b0 ;
  assign n4484 = n4463 | n4468 ;
  assign n4485 = ( ~n2269 & n4363 ) | ( ~n2269 & n4482 ) | ( n4363 & n4482 ) ;
  assign n4486 = ( ~n2139 & n4454 ) | ( ~n2139 & n4485 ) | ( n4454 & n4485 ) ;
  assign n4487 = ( ~n2009 & n4378 ) | ( ~n2009 & n4486 ) | ( n4378 & n4486 ) ;
  assign n4488 = ( ~n1885 & n4430 ) | ( ~n1885 & n4487 ) | ( n4430 & n4487 ) ;
  assign n4489 = ( ~n1766 & n4411 ) | ( ~n1766 & n4488 ) | ( n4411 & n4488 ) ;
  assign n4490 = ( ~n1652 & n4429 ) | ( ~n1652 & n4489 ) | ( n4429 & n4489 ) ;
  assign n4491 = ( ~n1534 & n4456 ) | ( ~n1534 & n4490 ) | ( n4456 & n4490 ) ;
  assign n4492 = ( ~n1416 & n4375 ) | ( ~n1416 & n4491 ) | ( n4375 & n4491 ) ;
  assign n4493 = ( ~n1318 & n4380 ) | ( ~n1318 & n4492 ) | ( n4380 & n4492 ) ;
  assign n4494 = ( ~n1220 & n4379 ) | ( ~n1220 & n4493 ) | ( n4379 & n4493 ) ;
  assign n4495 = ( ~n1118 & n4455 ) | ( ~n1118 & n4494 ) | ( n4455 & n4494 ) ;
  assign n4496 = ( ~n1034 & n4418 ) | ( ~n1034 & n4495 ) | ( n4418 & n4495 ) ;
  assign n4497 = ( ~n941 & n4421 ) | ( ~n941 & n4496 ) | ( n4421 & n4496 ) ;
  assign n4498 = ( ~n859 & n4438 ) | ( ~n859 & n4497 ) | ( n4438 & n4497 ) ;
  assign n4499 = ( ~n785 & n4453 ) | ( ~n785 & n4498 ) | ( n4453 & n4498 ) ;
  assign n4500 = n4488 ^ n1766 ^ 1'b0 ;
  assign n4501 = ( n4338 & n4342 ) | ( n4338 & n4346 ) | ( n4342 & n4346 ) ;
  assign n4502 = n4170 & ~n4501 ;
  assign n4503 = ( ~n716 & n4377 ) | ( ~n716 & n4499 ) | ( n4377 & n4499 ) ;
  assign n4504 = n4490 ^ n1534 ^ 1'b0 ;
  assign n4505 = n4502 ^ n4501 ^ n4342 ;
  assign n4506 = ( n4170 & ~n4338 ) | ( n4170 & n4346 ) | ( ~n4338 & n4346 ) ;
  assign n4507 = ( ~n640 & n4444 ) | ( ~n640 & n4503 ) | ( n4444 & n4503 ) ;
  assign n4508 = n4496 ^ n941 ^ 1'b0 ;
  assign n4509 = n4170 & ~n4338 ;
  assign n4510 = n4170 & ~n4346 ;
  assign n4511 = ( n4408 & n4506 ) | ( n4408 & ~n4509 ) | ( n4506 & ~n4509 ) ;
  assign n4512 = n4498 ^ n785 ^ 1'b0 ;
  assign n4513 = ( ~n572 & n4381 ) | ( ~n572 & n4507 ) | ( n4381 & n4507 ) ;
  assign n4514 = n4331 ^ n345 ^ 1'b0 ;
  assign n4515 = n4346 & n4470 ;
  assign n4516 = n4515 ^ n4227 ^ n4078 ;
  assign n4517 = ( ~n514 & n4449 ) | ( ~n514 & n4513 ) | ( n4449 & n4513 ) ;
  assign n4518 = n4346 & n4514 ;
  assign n4519 = n4518 ^ n4346 ^ n4225 ;
  assign n4520 = ( ~n458 & n4371 ) | ( ~n458 & n4517 ) | ( n4371 & n4517 ) ;
  assign n4521 = ( ~n399 & n4441 ) | ( ~n399 & n4520 ) | ( n4441 & n4520 ) ;
  assign n4522 = ( ~n345 & n4435 ) | ( ~n345 & n4521 ) | ( n4435 & n4521 ) ;
  assign n4523 = ( ~n302 & n4519 ) | ( ~n302 & n4522 ) | ( n4519 & n4522 ) ;
  assign n4524 = ( ~n261 & n4516 ) | ( ~n261 & n4523 ) | ( n4516 & n4523 ) ;
  assign n4525 = ( ~n217 & n4451 ) | ( ~n217 & n4524 ) | ( n4451 & n4524 ) ;
  assign n4526 = ( ~n179 & n4440 ) | ( ~n179 & n4525 ) | ( n4440 & n4525 ) ;
  assign n4527 = ( ~n144 & n4423 ) | ( ~n144 & n4526 ) | ( n4423 & n4526 ) ;
  assign n4528 = ( ~n134 & n4452 ) | ( ~n134 & n4527 ) | ( n4452 & n4527 ) ;
  assign n4529 = ( ~x30 & n4511 ) | ( ~x30 & n4528 ) | ( n4511 & n4528 ) ;
  assign n4530 = ~n136 & n4529 ;
  assign n4531 = n4408 & n4528 ;
  assign n4532 = n4510 | n4531 ;
  assign n4533 = n4530 | n4532 ;
  assign n4534 = n4505 | n4533 ;
  assign n4535 = n4484 & n4534 ;
  assign n4536 = n4535 ^ n4534 ^ n4458 ;
  assign n4537 = n4534 ^ n4475 ^ n3302 ;
  assign n4538 = n4534 & n4537 ;
  assign n4539 = n4538 ^ n4372 ^ n4264 ;
  assign n4540 = n4534 ^ n4476 ^ n3141 ;
  assign n4541 = n4534 & n4540 ;
  assign n4542 = n4534 ^ n4479 ^ n2690 ;
  assign n4543 = n4534 & n4542 ;
  assign n4544 = n4543 ^ n4400 ^ n4180 ;
  assign n4545 = n4483 & n4534 ;
  assign n4546 = n4545 ^ n4534 ^ n4391 ;
  assign n4547 = n4534 ^ n4482 ^ n2269 ;
  assign n4548 = n4534 & n4547 ;
  assign n4549 = n4548 ^ n4357 ^ n4188 ;
  assign n4550 = n4534 ^ n4485 ^ n2139 ;
  assign n4551 = n4534 & n4550 ;
  assign n4552 = n4551 ^ n4403 ^ n4285 ;
  assign n4553 = n4534 ^ n4486 ^ n2009 ;
  assign n4554 = n4534 & n4553 ;
  assign n4555 = n4554 ^ n4355 ^ n4233 ;
  assign n4556 = n4500 & n4534 ;
  assign n4557 = n4556 ^ n4534 ^ n4411 ;
  assign n4558 = n4504 & n4534 ;
  assign n4559 = n4558 ^ n4534 ^ n4456 ;
  assign n4560 = n4534 ^ n4492 ^ n1318 ;
  assign n4561 = n4534 & n4560 ;
  assign n4562 = n4561 ^ n4369 ^ n4198 ;
  assign n4563 = n4534 ^ n4495 ^ n1034 ;
  assign n4564 = n4541 ^ n4352 ^ n4175 ;
  assign n4565 = n4534 & n4563 ;
  assign n4566 = n4565 ^ n4404 ^ n4245 ;
  assign n4567 = n4508 & n4534 ;
  assign n4568 = n4567 ^ n4534 ^ n4421 ;
  assign n4569 = n4534 ^ n4497 ^ n859 ;
  assign n4570 = n4534 & n4569 ;
  assign n4571 = n4570 ^ n4436 ^ n4204 ;
  assign n4572 = n4512 & n4534 ;
  assign n4573 = n4572 ^ n4534 ^ n4453 ;
  assign n4574 = n4534 ^ n4503 ^ n640 ;
  assign n4575 = n4534 & n4574 ;
  assign n4576 = n4575 ^ n4443 ^ n4212 ;
  assign n4577 = n4534 ^ n4507 ^ n572 ;
  assign n4578 = n4534 & n4577 ;
  assign n4579 = n4578 ^ n4348 ^ n4215 ;
  assign n4580 = n4534 ^ n4517 ^ n458 ;
  assign n4581 = n4534 & n4580 ;
  assign n4582 = n4581 ^ n4367 ^ n4218 ;
  assign n4583 = n4520 ^ n399 ^ 1'b0 ;
  assign n4584 = n4534 & n4583 ;
  assign n4585 = n4584 ^ n4534 ^ n4441 ;
  assign n4586 = n4534 ^ n4521 ^ n345 ;
  assign n4587 = n4534 & n4586 ;
  assign n4588 = n4587 ^ n4434 ^ n4223 ;
  assign n4589 = n4534 ^ n4524 ^ n217 ;
  assign n4590 = n4534 & n4589 ;
  assign n4591 = n4590 ^ n4446 ^ n4251 ;
  assign n4592 = n4534 ^ n4525 ^ n179 ;
  assign n4593 = n4534 & n4592 ;
  assign n4594 = n4593 ^ n4439 ^ n4254 ;
  assign n4595 = n4534 ^ n4527 ^ n134 ;
  assign n4596 = n4534 & n4595 ;
  assign n4597 = n4596 ^ n4450 ^ n4265 ;
  assign n4598 = n4459 & n4534 ;
  assign n4599 = n4534 ^ n4474 ^ n3464 ;
  assign n4600 = n4534 & n4599 ;
  assign n4601 = n4600 ^ n4395 ^ n4259 ;
  assign n4602 = ( x64 & n4344 ) | ( x64 & n4534 ) | ( n4344 & n4534 ) ;
  assign n4603 = ( n4341 & ~n4344 ) | ( n4341 & n4602 ) | ( ~n4344 & n4602 ) ;
  assign n4604 = ~n4602 & n4603 ;
  assign n4605 = n4522 ^ n302 ^ 1'b0 ;
  assign n4606 = n4534 & n4605 ;
  assign n4607 = n4606 ^ n4534 ^ n4519 ;
  assign n4608 = ( n4346 & n4510 ) | ( n4346 & ~n4534 ) | ( n4510 & ~n4534 ) ;
  assign n4609 = n4534 ^ n4499 ^ n716 ;
  assign n4610 = n4505 | n4531 ;
  assign n4611 = ( x59 & x60 ) | ( x59 & ~n4505 ) | ( x60 & ~n4505 ) ;
  assign n4612 = ( x62 & ~n4505 ) | ( x62 & n4611 ) | ( ~n4505 & n4611 ) ;
  assign n4613 = ( ~n4510 & n4610 ) | ( ~n4510 & n4612 ) | ( n4610 & n4612 ) ;
  assign n4614 = ~n4610 & n4613 ;
  assign n4615 = ( n4408 & ~n4505 ) | ( n4408 & n4510 ) | ( ~n4505 & n4510 ) ;
  assign n4616 = ~n4533 & n4615 ;
  assign n4617 = n4534 ^ n4473 ^ n3631 ;
  assign n4618 = n4534 & n4617 ;
  assign n4619 = n4618 ^ n4465 ^ n4289 ;
  assign n4620 = n4478 ^ n2839 ^ 1'b0 ;
  assign n4621 = n4534 & n4620 ;
  assign n4622 = n4534 ^ n4481 ^ n2404 ;
  assign n4623 = n4534 ^ n4523 ^ n261 ;
  assign n4624 = n4534 ^ n4477 ^ n2995 ;
  assign n4625 = n4534 & n4623 ;
  assign n4626 = n4625 ^ n4515 ^ n4228 ;
  assign n4627 = n4534 ^ n4489 ^ n1652 ;
  assign n4628 = n4534 ^ n4526 ^ n144 ;
  assign n4629 = n4534 ^ n4487 ^ n1885 ;
  assign n4630 = n4534 ^ n4493 ^ n1220 ;
  assign n4631 = n4534 & n4609 ;
  assign n4632 = n4621 ^ n4534 ^ n4413 ;
  assign n4633 = n4534 ^ n4494 ^ n1118 ;
  assign n4634 = n4631 ^ n4374 ^ n4209 ;
  assign n4635 = n4534 & n4633 ;
  assign n4636 = n4472 ^ n3804 ^ 1'b0 ;
  assign n4637 = n4635 ^ n4437 ^ n4201 ;
  assign n4638 = n4534 & n4636 ;
  assign n4639 = n4534 & n4628 ;
  assign n4640 = n4639 ^ n4417 ^ n4239 ;
  assign n4641 = n4534 ^ n4513 ^ n514 ;
  assign n4642 = n4534 ^ n4491 ^ n1416 ;
  assign n4643 = n4534 & n4642 ;
  assign n4644 = ( n4528 & n4531 ) | ( n4528 & ~n4534 ) | ( n4531 & ~n4534 ) ;
  assign n4645 = n4638 ^ n4534 ^ n4364 ;
  assign n4646 = n4534 & n4641 ;
  assign n4647 = n4646 ^ n4448 ^ n4269 ;
  assign n4648 = ( n4534 & ~n4598 ) | ( n4534 & n4608 ) | ( ~n4598 & n4608 ) ;
  assign n4649 = n4534 & n4630 ;
  assign n4650 = n4534 & n4629 ;
  assign n4651 = n4650 ^ n4384 ^ n4191 ;
  assign n4652 = n4534 & n4624 ;
  assign n4653 = n4652 ^ n4410 ^ n4288 ;
  assign n4654 = n4534 & n4627 ;
  assign n4655 = n4654 ^ n4387 ^ n4276 ;
  assign n4656 = n4643 ^ n4366 ^ n4287 ;
  assign n4657 = n4649 ^ n4373 ^ n4272 ;
  assign n4658 = n4534 & n4622 ;
  assign n4659 = n4658 ^ n4426 ^ n4185 ;
  assign n4660 = ( ~x64 & n4346 ) | ( ~x64 & n4534 ) | ( n4346 & n4534 ) ;
  assign n4661 = ~x64 & n4534 ;
  assign n4662 = n4661 ^ x65 ^ 1'b0 ;
  assign n4663 = ( n136 & n4408 ) | ( n136 & n4528 ) | ( n4408 & n4528 ) ;
  assign n4664 = n4604 | n4662 ;
  assign n4665 = ~n4644 & n4663 ;
  assign n4666 = n4534 & ~n4616 ;
  assign n4667 = n4616 | n4665 ;
  assign n4668 = x62 | x63 ;
  assign n4669 = ( x64 & n4346 ) | ( x64 & ~n4668 ) | ( n4346 & ~n4668 ) ;
  assign n4670 = n4660 & n4669 ;
  assign n4671 = n4534 ^ n4469 ^ n3986 ;
  assign n4672 = n4534 & n4671 ;
  assign n4673 = n4672 ^ n4362 ^ x68 ;
  assign n4674 = n4648 ^ x66 ^ 1'b0 ;
  assign n4675 = n4664 & ~n4670 ;
  assign n4676 = ( ~n4167 & n4674 ) | ( ~n4167 & n4675 ) | ( n4674 & n4675 ) ;
  assign n4677 = ( ~n3986 & n4536 ) | ( ~n3986 & n4676 ) | ( n4536 & n4676 ) ;
  assign n4678 = ( ~n3804 & n4673 ) | ( ~n3804 & n4677 ) | ( n4673 & n4677 ) ;
  assign n4679 = ( ~n3631 & n4645 ) | ( ~n3631 & n4678 ) | ( n4645 & n4678 ) ;
  assign n4680 = ( ~n3464 & n4619 ) | ( ~n3464 & n4679 ) | ( n4619 & n4679 ) ;
  assign n4681 = ( ~n3302 & n4601 ) | ( ~n3302 & n4680 ) | ( n4601 & n4680 ) ;
  assign n4682 = ( ~n3141 & n4539 ) | ( ~n3141 & n4681 ) | ( n4539 & n4681 ) ;
  assign n4683 = ( ~n2995 & n4564 ) | ( ~n2995 & n4682 ) | ( n4564 & n4682 ) ;
  assign n4684 = ( ~n2839 & n4653 ) | ( ~n2839 & n4683 ) | ( n4653 & n4683 ) ;
  assign n4685 = ( ~n2690 & n4632 ) | ( ~n2690 & n4684 ) | ( n4632 & n4684 ) ;
  assign n4686 = ( ~n2544 & n4544 ) | ( ~n2544 & n4685 ) | ( n4544 & n4685 ) ;
  assign n4687 = ( ~n2404 & n4546 ) | ( ~n2404 & n4686 ) | ( n4546 & n4686 ) ;
  assign n4688 = ( ~n2269 & n4659 ) | ( ~n2269 & n4687 ) | ( n4659 & n4687 ) ;
  assign n4689 = ( ~n2139 & n4549 ) | ( ~n2139 & n4688 ) | ( n4549 & n4688 ) ;
  assign n4690 = ( ~n2009 & n4552 ) | ( ~n2009 & n4689 ) | ( n4552 & n4689 ) ;
  assign n4691 = ( ~n1885 & n4555 ) | ( ~n1885 & n4690 ) | ( n4555 & n4690 ) ;
  assign n4692 = ( ~n1766 & n4651 ) | ( ~n1766 & n4691 ) | ( n4651 & n4691 ) ;
  assign n4693 = ( ~n1652 & n4557 ) | ( ~n1652 & n4692 ) | ( n4557 & n4692 ) ;
  assign n4694 = ( ~n4408 & n4528 ) | ( ~n4408 & n4534 ) | ( n4528 & n4534 ) ;
  assign n4695 = ( ~n1534 & n4655 ) | ( ~n1534 & n4693 ) | ( n4655 & n4693 ) ;
  assign n4696 = ( ~n1416 & n4559 ) | ( ~n1416 & n4695 ) | ( n4559 & n4695 ) ;
  assign n4697 = ( ~n1318 & n4656 ) | ( ~n1318 & n4696 ) | ( n4656 & n4696 ) ;
  assign n4698 = ( ~n1220 & n4562 ) | ( ~n1220 & n4697 ) | ( n4562 & n4697 ) ;
  assign n4699 = ( ~n1118 & n4657 ) | ( ~n1118 & n4698 ) | ( n4657 & n4698 ) ;
  assign n4700 = ( ~n1034 & n4637 ) | ( ~n1034 & n4699 ) | ( n4637 & n4699 ) ;
  assign n4701 = ( ~n941 & n4566 ) | ( ~n941 & n4700 ) | ( n4566 & n4700 ) ;
  assign n4702 = ( ~n859 & n4568 ) | ( ~n859 & n4701 ) | ( n4568 & n4701 ) ;
  assign n4703 = ( ~n785 & n4571 ) | ( ~n785 & n4702 ) | ( n4571 & n4702 ) ;
  assign n4704 = ~n4408 & n4528 ;
  assign n4705 = n4692 ^ n1652 ^ 1'b0 ;
  assign n4706 = n4686 ^ n2404 ^ 1'b0 ;
  assign n4707 = n4701 ^ n859 ^ 1'b0 ;
  assign n4708 = ( ~n716 & n4573 ) | ( ~n716 & n4703 ) | ( n4573 & n4703 ) ;
  assign n4709 = n4695 ^ n1416 ^ 1'b0 ;
  assign n4710 = n4678 ^ n3631 ^ 1'b0 ;
  assign n4711 = n4703 ^ n716 ^ 1'b0 ;
  assign n4712 = n4684 ^ n2690 ^ 1'b0 ;
  assign n4713 = ( ~n640 & n4634 ) | ( ~n640 & n4708 ) | ( n4634 & n4708 ) ;
  assign n4714 = ( ~n572 & n4576 ) | ( ~n572 & n4713 ) | ( n4576 & n4713 ) ;
  assign n4715 = ( ~n514 & n4579 ) | ( ~n514 & n4714 ) | ( n4579 & n4714 ) ;
  assign n4716 = ( ~n458 & n4647 ) | ( ~n458 & n4715 ) | ( n4647 & n4715 ) ;
  assign n4717 = ( ~n399 & n4582 ) | ( ~n399 & n4716 ) | ( n4582 & n4716 ) ;
  assign n4718 = ( ~n345 & n4585 ) | ( ~n345 & n4717 ) | ( n4585 & n4717 ) ;
  assign n4719 = ( ~n302 & n4588 ) | ( ~n302 & n4718 ) | ( n4588 & n4718 ) ;
  assign n4720 = ( ~n261 & n4607 ) | ( ~n261 & n4719 ) | ( n4607 & n4719 ) ;
  assign n4721 = ( ~n217 & n4626 ) | ( ~n217 & n4720 ) | ( n4626 & n4720 ) ;
  assign n4722 = ( ~n179 & n4591 ) | ( ~n179 & n4721 ) | ( n4591 & n4721 ) ;
  assign n4723 = ( ~n144 & n4594 ) | ( ~n144 & n4722 ) | ( n4594 & n4722 ) ;
  assign n4724 = ( ~n134 & n4640 ) | ( ~n134 & n4723 ) | ( n4640 & n4723 ) ;
  assign n4725 = ( ~n136 & n4597 ) | ( ~n136 & n4724 ) | ( n4597 & n4724 ) ;
  assign n4726 = ( ~n136 & n4694 ) | ( ~n136 & n4725 ) | ( n4694 & n4725 ) ;
  assign n4727 = ( ~n4704 & n4725 ) | ( ~n4704 & n4726 ) | ( n4725 & n4726 ) ;
  assign n4728 = n4667 | n4727 ;
  assign n4729 = n4728 ^ n4723 ^ n134 ;
  assign n4730 = n4728 & n4729 ;
  assign n4731 = n4730 ^ n4639 ^ n4423 ;
  assign n4732 = ~n4668 & n4728 ;
  assign n4733 = ( n4665 & n4727 ) | ( n4665 & ~n4732 ) | ( n4727 & ~n4732 ) ;
  assign n4734 = n4666 | n4732 ;
  assign n4735 = ( n4732 & ~n4733 ) | ( n4732 & n4734 ) | ( ~n4733 & n4734 ) ;
  assign n4736 = ( x62 & n4530 ) | ( x62 & n4728 ) | ( n4530 & n4728 ) ;
  assign n4737 = ( ~n4530 & n4614 ) | ( ~n4530 & n4736 ) | ( n4614 & n4736 ) ;
  assign n4738 = ~n4736 & n4737 ;
  assign n4739 = ( n4604 & ~n4670 ) | ( n4604 & n4728 ) | ( ~n4670 & n4728 ) ;
  assign n4740 = ~n4604 & n4739 ;
  assign n4741 = n4728 ^ n4677 ^ n3804 ;
  assign n4742 = n4728 & n4741 ;
  assign n4743 = n4742 ^ n4672 ^ n4471 ;
  assign n4744 = n4710 & n4728 ;
  assign n4745 = n4744 ^ n4728 ^ n4645 ;
  assign n4746 = n4728 ^ n4679 ^ n3464 ;
  assign n4747 = n4728 & n4746 ;
  assign n4748 = n4747 ^ n4618 ^ n4466 ;
  assign n4749 = n4728 ^ n4681 ^ n3141 ;
  assign n4750 = n4728 & n4749 ;
  assign n4751 = n4750 ^ n4538 ^ n4376 ;
  assign n4752 = n4712 & n4728 ;
  assign n4753 = n4752 ^ n4728 ^ n4632 ;
  assign n4754 = n4706 & n4728 ;
  assign n4755 = n4754 ^ n4728 ^ n4546 ;
  assign n4756 = n4728 ^ n4688 ^ n2139 ;
  assign n4757 = n4728 & n4756 ;
  assign n4758 = n4757 ^ n4548 ^ n4363 ;
  assign n4759 = n4728 ^ n4690 ^ n1885 ;
  assign n4760 = n4728 & n4759 ;
  assign n4761 = n4760 ^ n4554 ^ n4378 ;
  assign n4762 = n4705 & n4728 ;
  assign n4763 = n4762 ^ n4728 ^ n4557 ;
  assign n4764 = n4728 ^ n4693 ^ n1534 ;
  assign n4765 = n4728 & n4764 ;
  assign n4766 = n4765 ^ n4654 ^ n4429 ;
  assign n4767 = n4709 & n4728 ;
  assign n4768 = n4767 ^ n4728 ^ n4559 ;
  assign n4769 = n4728 ^ n4696 ^ n1318 ;
  assign n4770 = n4728 & n4769 ;
  assign n4771 = n4770 ^ n4643 ^ n4375 ;
  assign n4772 = n4728 ^ n4697 ^ n1220 ;
  assign n4773 = n4728 & n4772 ;
  assign n4774 = n4773 ^ n4561 ^ n4380 ;
  assign n4775 = n4728 ^ n4698 ^ n1118 ;
  assign n4776 = n4728 & n4775 ;
  assign n4777 = n4776 ^ n4649 ^ n4379 ;
  assign n4778 = n4728 ^ n4700 ^ n941 ;
  assign n4779 = n4728 & n4778 ;
  assign n4780 = n4779 ^ n4565 ^ n4418 ;
  assign n4781 = n4707 & n4728 ;
  assign n4782 = n4781 ^ n4728 ^ n4568 ;
  assign n4783 = n4711 & n4728 ;
  assign n4784 = n4783 ^ n4728 ^ n4573 ;
  assign n4785 = n4728 ^ n4722 ^ n144 ;
  assign n4786 = n4728 & n4785 ;
  assign n4787 = n4786 ^ n4593 ^ n4440 ;
  assign n4788 = n4740 ^ n4661 ^ x65 ;
  assign n4789 = n4728 ^ n4675 ^ n4167 ;
  assign n4790 = n4728 & n4789 ;
  assign n4791 = n4790 ^ n4648 ^ x66 ;
  assign n4792 = n4676 ^ n3986 ^ 1'b0 ;
  assign n4793 = n4728 & n4792 ;
  assign n4794 = n4793 ^ n4728 ^ n4536 ;
  assign n4795 = n4728 ^ n4680 ^ n3302 ;
  assign n4796 = n4728 & n4795 ;
  assign n4797 = n4796 ^ n4600 ^ n4431 ;
  assign n4798 = n4728 ^ n4682 ^ n2995 ;
  assign n4799 = n4728 & n4798 ;
  assign n4800 = n4799 ^ n4541 ^ n4353 ;
  assign n4801 = n4728 ^ n4683 ^ n2839 ;
  assign n4802 = n4728 & n4801 ;
  assign n4803 = n4802 ^ n4652 ^ n4428 ;
  assign n4804 = n4728 ^ n4685 ^ n2544 ;
  assign n4805 = n4728 & n4804 ;
  assign n4806 = n4805 ^ n4543 ^ n4422 ;
  assign n4807 = n4728 ^ n4687 ^ n2269 ;
  assign n4808 = n4728 & n4807 ;
  assign n4809 = n4808 ^ n4658 ^ n4427 ;
  assign n4810 = n4728 ^ n4689 ^ n2009 ;
  assign n4811 = n4728 & n4810 ;
  assign n4812 = n4811 ^ n4551 ^ n4454 ;
  assign n4813 = n4728 ^ n4691 ^ n1766 ;
  assign n4814 = n4728 & n4813 ;
  assign n4815 = n4814 ^ n4650 ^ n4430 ;
  assign n4816 = n4728 ^ n4699 ^ n1034 ;
  assign n4817 = n4728 & n4816 ;
  assign n4818 = n4817 ^ n4635 ^ n4455 ;
  assign n4819 = n4728 ^ n4702 ^ n785 ;
  assign n4820 = n4728 & n4819 ;
  assign n4821 = n4820 ^ n4570 ^ n4438 ;
  assign n4822 = n4728 ^ n4708 ^ n640 ;
  assign n4823 = n4728 & n4822 ;
  assign n4824 = n4823 ^ n4631 ^ n4377 ;
  assign n4825 = n4728 ^ n4713 ^ n572 ;
  assign n4826 = n4728 & n4825 ;
  assign n4827 = n4728 ^ n4714 ^ n514 ;
  assign n4828 = n4728 & n4827 ;
  assign n4829 = n4828 ^ n4578 ^ n4381 ;
  assign n4830 = n4728 ^ n4715 ^ n458 ;
  assign n4831 = n4728 & n4830 ;
  assign n4832 = n4831 ^ n4646 ^ n4449 ;
  assign n4833 = n4728 ^ n4716 ^ n399 ;
  assign n4834 = n4826 ^ n4575 ^ n4444 ;
  assign n4835 = n4728 & n4833 ;
  assign n4836 = n4835 ^ n4581 ^ n4371 ;
  assign n4837 = n4717 ^ n345 ^ 1'b0 ;
  assign n4838 = n4728 & n4837 ;
  assign n4839 = n4838 ^ n4728 ^ n4585 ;
  assign n4840 = n4728 ^ n4718 ^ n302 ;
  assign n4841 = n4728 & n4840 ;
  assign n4842 = n4841 ^ n4587 ^ n4435 ;
  assign n4843 = n4719 ^ n261 ^ 1'b0 ;
  assign n4844 = n4728 & n4843 ;
  assign n4845 = n4844 ^ n4728 ^ n4607 ;
  assign n4846 = n4728 ^ n4720 ^ n217 ;
  assign n4847 = n4728 & n4846 ;
  assign n4848 = n4847 ^ n4625 ^ n4516 ;
  assign n4849 = n4728 ^ n4721 ^ n179 ;
  assign n4850 = n4728 & n4849 ;
  assign n4851 = n4850 ^ n4590 ^ n4451 ;
  assign n4852 = ~x62 & n4728 ;
  assign n4853 = x59 | x60 ;
  assign n4854 = ( x62 & n4534 ) | ( x62 & ~n4853 ) | ( n4534 & ~n4853 ) ;
  assign n4855 = n4852 ^ x63 ^ 1'b0 ;
  assign n4856 = n4738 | n4855 ;
  assign n4857 = ( ~x62 & n4534 ) | ( ~x62 & n4728 ) | ( n4534 & n4728 ) ;
  assign n4858 = n4854 & n4857 ;
  assign n4859 = n4856 & ~n4858 ;
  assign n4860 = n4735 ^ x64 ^ 1'b0 ;
  assign n4861 = ( ~n4346 & n4859 ) | ( ~n4346 & n4860 ) | ( n4859 & n4860 ) ;
  assign n4862 = ( ~n4167 & n4788 ) | ( ~n4167 & n4861 ) | ( n4788 & n4861 ) ;
  assign n4863 = ( ~n3986 & n4791 ) | ( ~n3986 & n4862 ) | ( n4791 & n4862 ) ;
  assign n4864 = ( ~n3804 & n4794 ) | ( ~n3804 & n4863 ) | ( n4794 & n4863 ) ;
  assign n4865 = ( ~n3631 & n4743 ) | ( ~n3631 & n4864 ) | ( n4743 & n4864 ) ;
  assign n4866 = ( ~n3464 & n4745 ) | ( ~n3464 & n4865 ) | ( n4745 & n4865 ) ;
  assign n4867 = ( ~n3302 & n4748 ) | ( ~n3302 & n4866 ) | ( n4748 & n4866 ) ;
  assign n4868 = ( ~n3141 & n4797 ) | ( ~n3141 & n4867 ) | ( n4797 & n4867 ) ;
  assign n4869 = ( ~n2995 & n4751 ) | ( ~n2995 & n4868 ) | ( n4751 & n4868 ) ;
  assign n4870 = ( ~n2839 & n4800 ) | ( ~n2839 & n4869 ) | ( n4800 & n4869 ) ;
  assign n4871 = ( ~n2690 & n4803 ) | ( ~n2690 & n4870 ) | ( n4803 & n4870 ) ;
  assign n4872 = ( ~n2544 & n4753 ) | ( ~n2544 & n4871 ) | ( n4753 & n4871 ) ;
  assign n4873 = ( ~n2404 & n4806 ) | ( ~n2404 & n4872 ) | ( n4806 & n4872 ) ;
  assign n4874 = ( ~n2269 & n4755 ) | ( ~n2269 & n4873 ) | ( n4755 & n4873 ) ;
  assign n4875 = ( ~n2139 & n4809 ) | ( ~n2139 & n4874 ) | ( n4809 & n4874 ) ;
  assign n4876 = ( ~n4597 & n4724 ) | ( ~n4597 & n4728 ) | ( n4724 & n4728 ) ;
  assign n4877 = ~n4597 & n4724 ;
  assign n4878 = ( ~n2009 & n4758 ) | ( ~n2009 & n4875 ) | ( n4758 & n4875 ) ;
  assign n4879 = ( ~n1885 & n4812 ) | ( ~n1885 & n4878 ) | ( n4812 & n4878 ) ;
  assign n4880 = ( ~n1766 & n4761 ) | ( ~n1766 & n4879 ) | ( n4761 & n4879 ) ;
  assign n4881 = ( n4597 & n4724 ) | ( n4597 & ~n4728 ) | ( n4724 & ~n4728 ) ;
  assign n4882 = ( ~n1652 & n4815 ) | ( ~n1652 & n4880 ) | ( n4815 & n4880 ) ;
  assign n4883 = ( ~n1534 & n4763 ) | ( ~n1534 & n4882 ) | ( n4763 & n4882 ) ;
  assign n4884 = ( ~n1416 & n4766 ) | ( ~n1416 & n4883 ) | ( n4766 & n4883 ) ;
  assign n4885 = ( ~n1318 & n4768 ) | ( ~n1318 & n4884 ) | ( n4768 & n4884 ) ;
  assign n4886 = ( ~n1220 & n4771 ) | ( ~n1220 & n4885 ) | ( n4771 & n4885 ) ;
  assign n4887 = ( ~n1118 & n4774 ) | ( ~n1118 & n4886 ) | ( n4774 & n4886 ) ;
  assign n4888 = ( ~n1034 & n4777 ) | ( ~n1034 & n4887 ) | ( n4777 & n4887 ) ;
  assign n4889 = ( ~n941 & n4818 ) | ( ~n941 & n4888 ) | ( n4818 & n4888 ) ;
  assign n4890 = ( ~n859 & n4780 ) | ( ~n859 & n4889 ) | ( n4780 & n4889 ) ;
  assign n4891 = ( ~n785 & n4782 ) | ( ~n785 & n4890 ) | ( n4782 & n4890 ) ;
  assign n4892 = ( n4731 & n4876 ) | ( n4731 & ~n4877 ) | ( n4876 & ~n4877 ) ;
  assign n4893 = ( n136 & n4597 ) | ( n136 & n4724 ) | ( n4597 & n4724 ) ;
  assign n4894 = ~n4724 & n4893 ;
  assign n4895 = ( ~n4881 & n4893 ) | ( ~n4881 & n4894 ) | ( n4893 & n4894 ) ;
  assign n4896 = ( ~n716 & n4821 ) | ( ~n716 & n4891 ) | ( n4821 & n4891 ) ;
  assign n4897 = ( ~n640 & n4784 ) | ( ~n640 & n4896 ) | ( n4784 & n4896 ) ;
  assign n4898 = ( ~n572 & n4824 ) | ( ~n572 & n4897 ) | ( n4824 & n4897 ) ;
  assign n4899 = ( ~n514 & n4834 ) | ( ~n514 & n4898 ) | ( n4834 & n4898 ) ;
  assign n4900 = ( ~n458 & n4829 ) | ( ~n458 & n4899 ) | ( n4829 & n4899 ) ;
  assign n4901 = ( ~n399 & n4832 ) | ( ~n399 & n4900 ) | ( n4832 & n4900 ) ;
  assign n4902 = ( ~n345 & n4836 ) | ( ~n345 & n4901 ) | ( n4836 & n4901 ) ;
  assign n4903 = ( ~n302 & n4839 ) | ( ~n302 & n4902 ) | ( n4839 & n4902 ) ;
  assign n4904 = ( ~n261 & n4842 ) | ( ~n261 & n4903 ) | ( n4842 & n4903 ) ;
  assign n4905 = ( ~n217 & n4845 ) | ( ~n217 & n4904 ) | ( n4845 & n4904 ) ;
  assign n4906 = ( ~n179 & n4848 ) | ( ~n179 & n4905 ) | ( n4848 & n4905 ) ;
  assign n4907 = ( ~n144 & n4851 ) | ( ~n144 & n4906 ) | ( n4851 & n4906 ) ;
  assign n4908 = ( ~n134 & n4787 ) | ( ~n134 & n4907 ) | ( n4787 & n4907 ) ;
  assign n4909 = n4731 & n4908 ;
  assign n4910 = ( n4597 & ~n4728 ) | ( n4597 & n4909 ) | ( ~n4728 & n4909 ) ;
  assign n4911 = ( ~x30 & n4892 ) | ( ~x30 & n4908 ) | ( n4892 & n4908 ) ;
  assign n4912 = ~n136 & n4911 ;
  assign n4913 = n4909 | n4912 ;
  assign n4914 = ( n4895 & ~n4910 ) | ( n4895 & n4913 ) | ( ~n4910 & n4913 ) ;
  assign n4915 = n4910 | n4914 ;
  assign n4916 = n4915 ^ n4907 ^ n134 ;
  assign n4917 = n4915 & n4916 ;
  assign n4918 = n4917 ^ n4786 ^ n4594 ;
  assign n4919 = ( n4738 & ~n4858 ) | ( n4738 & n4915 ) | ( ~n4858 & n4915 ) ;
  assign n4920 = ~n4738 & n4919 ;
  assign n4921 = n4915 ^ n4861 ^ n4167 ;
  assign n4922 = n4915 & n4921 ;
  assign n4923 = n4922 ^ n4740 ^ n4662 ;
  assign n4924 = n4915 ^ n4864 ^ n3631 ;
  assign n4925 = n4915 & n4924 ;
  assign n4926 = n4925 ^ n4742 ^ n4673 ;
  assign n4927 = n4915 ^ n4868 ^ n2995 ;
  assign n4928 = n4915 & n4927 ;
  assign n4929 = n4928 ^ n4750 ^ n4539 ;
  assign n4930 = n4915 ^ n4869 ^ n2839 ;
  assign n4931 = n4915 & n4930 ;
  assign n4932 = n4931 ^ n4799 ^ n4564 ;
  assign n4933 = n4915 ^ n4875 ^ n2009 ;
  assign n4934 = n4915 & n4933 ;
  assign n4935 = n4934 ^ n4757 ^ n4549 ;
  assign n4936 = n4915 ^ n4878 ^ n1885 ;
  assign n4937 = n4915 & n4936 ;
  assign n4938 = n4937 ^ n4811 ^ n4552 ;
  assign n4939 = n4915 ^ n4879 ^ n1766 ;
  assign n4940 = n4915 & n4939 ;
  assign n4941 = n4940 ^ n4760 ^ n4555 ;
  assign n4942 = n4915 ^ n4885 ^ n1220 ;
  assign n4943 = n4915 & n4942 ;
  assign n4944 = n4943 ^ n4770 ^ n4656 ;
  assign n4945 = n4915 ^ n4886 ^ n1118 ;
  assign n4946 = n4915 & n4945 ;
  assign n4947 = n4946 ^ n4773 ^ n4562 ;
  assign n4948 = n4915 ^ n4898 ^ n514 ;
  assign n4949 = n4915 & n4948 ;
  assign n4950 = n4949 ^ n4826 ^ n4576 ;
  assign n4951 = n4915 ^ n4903 ^ n261 ;
  assign n4952 = n4915 & n4951 ;
  assign n4953 = n4952 ^ n4841 ^ n4588 ;
  assign n4954 = n4915 ^ n4862 ^ n3986 ;
  assign n4955 = n4863 ^ n3804 ^ 1'b0 ;
  assign n4956 = n4915 & n4955 ;
  assign n4957 = n4956 ^ n4915 ^ n4794 ;
  assign n4958 = n4865 ^ n3464 ^ 1'b0 ;
  assign n4959 = n4915 & n4958 ;
  assign n4960 = n4959 ^ n4915 ^ n4745 ;
  assign n4961 = n4871 ^ n2544 ^ 1'b0 ;
  assign n4962 = n4915 & n4961 ;
  assign n4963 = n4962 ^ n4915 ^ n4753 ;
  assign n4964 = n4915 ^ n4872 ^ n2404 ;
  assign n4965 = n4915 & n4964 ;
  assign n4966 = n4965 ^ n4805 ^ n4544 ;
  assign n4967 = n4873 ^ n2269 ^ 1'b0 ;
  assign n4968 = n4915 & n4967 ;
  assign n4969 = n4968 ^ n4915 ^ n4755 ;
  assign n4970 = n4915 ^ n4880 ^ n1652 ;
  assign n4971 = n4915 & n4954 ;
  assign n4972 = n4971 ^ n4790 ^ n4674 ;
  assign n4973 = n4915 & n4970 ;
  assign n4974 = n4973 ^ n4814 ^ n4651 ;
  assign n4975 = n4882 ^ n1534 ^ 1'b0 ;
  assign n4976 = n4915 & n4975 ;
  assign n4977 = n4976 ^ n4915 ^ n4763 ;
  assign n4978 = n4884 ^ n1318 ^ 1'b0 ;
  assign n4979 = n4915 & n4978 ;
  assign n4980 = n4915 ^ n4888 ^ n941 ;
  assign n4981 = n4915 & n4980 ;
  assign n4982 = n4981 ^ n4817 ^ n4637 ;
  assign n4983 = n4890 ^ n785 ^ 1'b0 ;
  assign n4984 = n4915 & n4983 ;
  assign n4985 = n4984 ^ n4915 ^ n4782 ;
  assign n4986 = n4896 ^ n640 ^ 1'b0 ;
  assign n4987 = n4915 & n4986 ;
  assign n4988 = n4987 ^ n4915 ^ n4784 ;
  assign n4989 = n4979 ^ n4915 ^ n4768 ;
  assign n4990 = n4915 ^ n4897 ^ n572 ;
  assign n4991 = n4915 & n4990 ;
  assign n4992 = n4991 ^ n4823 ^ n4634 ;
  assign n4993 = n4902 ^ n302 ^ 1'b0 ;
  assign n4994 = n4915 & n4993 ;
  assign n4995 = n4994 ^ n4915 ^ n4839 ;
  assign n4996 = n4904 ^ n217 ^ 1'b0 ;
  assign n4997 = n4915 & n4996 ;
  assign n4998 = n4997 ^ n4915 ^ n4845 ;
  assign n4999 = n4915 ^ n4906 ^ n144 ;
  assign n5000 = n4915 ^ n4866 ^ n3302 ;
  assign n5001 = n4915 & n5000 ;
  assign n5002 = n5001 ^ n4747 ^ n4619 ;
  assign n5003 = n4915 ^ n4867 ^ n3141 ;
  assign n5004 = n4915 & n5003 ;
  assign n5005 = n5004 ^ n4796 ^ n4601 ;
  assign n5006 = n4915 ^ n4870 ^ n2690 ;
  assign n5007 = n4915 & n5006 ;
  assign n5008 = n5007 ^ n4802 ^ n4653 ;
  assign n5009 = n4915 ^ n4874 ^ n2139 ;
  assign n5010 = n4915 & n5009 ;
  assign n5011 = n5010 ^ n4808 ^ n4659 ;
  assign n5012 = n4915 ^ n4887 ^ n1034 ;
  assign n5013 = n4915 & n5012 ;
  assign n5014 = n5013 ^ n4776 ^ n4657 ;
  assign n5015 = n4915 ^ n4889 ^ n859 ;
  assign n5016 = n4915 & n5015 ;
  assign n5017 = n5016 ^ n4779 ^ n4566 ;
  assign n5018 = n4915 ^ n4891 ^ n716 ;
  assign n5019 = n4915 & n5018 ;
  assign n5020 = n5019 ^ n4820 ^ n4571 ;
  assign n5021 = n4915 ^ n4899 ^ n458 ;
  assign n5022 = n4915 & n5021 ;
  assign n5023 = n5022 ^ n4828 ^ n4579 ;
  assign n5024 = n4915 ^ n4900 ^ n399 ;
  assign n5025 = n4915 & n5024 ;
  assign n5026 = n5025 ^ n4831 ^ n4647 ;
  assign n5027 = n4915 ^ n4901 ^ n345 ;
  assign n5028 = n4915 ^ n4883 ^ n1416 ;
  assign n5029 = n4915 & n5028 ;
  assign n5030 = n5029 ^ n4765 ^ n4655 ;
  assign n5031 = n4915 & n5027 ;
  assign n5032 = n5031 ^ n4835 ^ n4582 ;
  assign n5033 = n4915 ^ n4905 ^ n179 ;
  assign n5034 = n4915 & n5033 ;
  assign n5035 = n5034 ^ n4847 ^ n4626 ;
  assign n5036 = n4915 & n4999 ;
  assign n5037 = n5036 ^ n4850 ^ n4591 ;
  assign n5038 = n4915 ^ n4859 ^ n4346 ;
  assign n5039 = n4915 & n5038 ;
  assign n5040 = x57 | x58 ;
  assign n5041 = ( x59 & ~n4727 ) | ( x59 & n5040 ) | ( ~n4727 & n5040 ) ;
  assign n5042 = x59 & n4915 ;
  assign n5043 = ~n4853 & n4915 ;
  assign n5044 = n5039 ^ n4735 ^ x64 ;
  assign n5045 = ( n4728 & ~n4913 ) | ( n4728 & n5043 ) | ( ~n4913 & n5043 ) ;
  assign n5046 = n4895 & ~n5043 ;
  assign n5047 = n4920 ^ n4852 ^ x63 ;
  assign n5048 = ( n5043 & n5045 ) | ( n5043 & ~n5046 ) | ( n5045 & ~n5046 ) ;
  assign n5049 = ( ~n4728 & n5041 ) | ( ~n4728 & n5042 ) | ( n5041 & n5042 ) ;
  assign n5050 = n5048 ^ x62 ^ 1'b0 ;
  assign n5051 = ~n5042 & n5049 ;
  assign n5052 = n5042 ^ n4915 ^ x60 ;
  assign n5053 = n5051 | n5052 ;
  assign n5054 = ( ~x59 & n4728 ) | ( ~x59 & n4915 ) | ( n4728 & n4915 ) ;
  assign n5055 = ( x59 & n4728 ) | ( x59 & ~n5040 ) | ( n4728 & ~n5040 ) ;
  assign n5056 = ( n136 & n4731 ) | ( n136 & n4908 ) | ( n4731 & n4908 ) ;
  assign n5057 = n5054 & n5055 ;
  assign n5058 = n5053 & ~n5057 ;
  assign n5059 = ( ~n4534 & n5050 ) | ( ~n4534 & n5058 ) | ( n5050 & n5058 ) ;
  assign n5060 = ( ~n4346 & n5047 ) | ( ~n4346 & n5059 ) | ( n5047 & n5059 ) ;
  assign n5061 = ( ~n4167 & n5044 ) | ( ~n4167 & n5060 ) | ( n5044 & n5060 ) ;
  assign n5062 = ( ~n3986 & n4923 ) | ( ~n3986 & n5061 ) | ( n4923 & n5061 ) ;
  assign n5063 = ( ~n3804 & n4972 ) | ( ~n3804 & n5062 ) | ( n4972 & n5062 ) ;
  assign n5064 = ( ~n3631 & n4957 ) | ( ~n3631 & n5063 ) | ( n4957 & n5063 ) ;
  assign n5065 = ( n4908 & n4909 ) | ( n4908 & ~n4915 ) | ( n4909 & ~n4915 ) ;
  assign n5066 = n5056 & ~n5065 ;
  assign n5067 = ( ~n4731 & n4909 ) | ( ~n4731 & n4915 ) | ( n4909 & n4915 ) ;
  assign n5068 = n4731 & ~n4915 ;
  assign n5069 = ( ~n3464 & n4926 ) | ( ~n3464 & n5064 ) | ( n4926 & n5064 ) ;
  assign n5070 = ( ~n3302 & n4960 ) | ( ~n3302 & n5069 ) | ( n4960 & n5069 ) ;
  assign n5071 = n5069 ^ n3302 ^ 1'b0 ;
  assign n5072 = ( ~n3141 & n5002 ) | ( ~n3141 & n5070 ) | ( n5002 & n5070 ) ;
  assign n5073 = n4908 & ~n4909 ;
  assign n5074 = ( ~n2995 & n5005 ) | ( ~n2995 & n5072 ) | ( n5005 & n5072 ) ;
  assign n5075 = ( ~n2839 & n4929 ) | ( ~n2839 & n5074 ) | ( n4929 & n5074 ) ;
  assign n5076 = ( ~n2690 & n4932 ) | ( ~n2690 & n5075 ) | ( n4932 & n5075 ) ;
  assign n5077 = ( ~n2544 & n5008 ) | ( ~n2544 & n5076 ) | ( n5008 & n5076 ) ;
  assign n5078 = ( ~n2404 & n4963 ) | ( ~n2404 & n5077 ) | ( n4963 & n5077 ) ;
  assign n5079 = ( ~n2269 & n4966 ) | ( ~n2269 & n5078 ) | ( n4966 & n5078 ) ;
  assign n5080 = ( ~n2139 & n4969 ) | ( ~n2139 & n5079 ) | ( n4969 & n5079 ) ;
  assign n5081 = ( ~n2009 & n5011 ) | ( ~n2009 & n5080 ) | ( n5011 & n5080 ) ;
  assign n5082 = ( ~n1885 & n4935 ) | ( ~n1885 & n5081 ) | ( n4935 & n5081 ) ;
  assign n5083 = ( ~n1766 & n4938 ) | ( ~n1766 & n5082 ) | ( n4938 & n5082 ) ;
  assign n5084 = ( ~n1652 & n4941 ) | ( ~n1652 & n5083 ) | ( n4941 & n5083 ) ;
  assign n5085 = ( ~n1534 & n4974 ) | ( ~n1534 & n5084 ) | ( n4974 & n5084 ) ;
  assign n5086 = ( ~n1416 & n4977 ) | ( ~n1416 & n5085 ) | ( n4977 & n5085 ) ;
  assign n5087 = ( ~n1318 & n5030 ) | ( ~n1318 & n5086 ) | ( n5030 & n5086 ) ;
  assign n5088 = ( ~n1220 & n4989 ) | ( ~n1220 & n5087 ) | ( n4989 & n5087 ) ;
  assign n5089 = ( ~n1118 & n4944 ) | ( ~n1118 & n5088 ) | ( n4944 & n5088 ) ;
  assign n5090 = ( ~n1034 & n4947 ) | ( ~n1034 & n5089 ) | ( n4947 & n5089 ) ;
  assign n5091 = ( ~n941 & n5014 ) | ( ~n941 & n5090 ) | ( n5014 & n5090 ) ;
  assign n5092 = n5077 ^ n2404 ^ 1'b0 ;
  assign n5093 = n5079 ^ n2139 ^ 1'b0 ;
  assign n5094 = ( ~n859 & n4982 ) | ( ~n859 & n5091 ) | ( n4982 & n5091 ) ;
  assign n5095 = ( n4909 & n5067 ) | ( n4909 & ~n5073 ) | ( n5067 & ~n5073 ) ;
  assign n5096 = ( ~n785 & n5017 ) | ( ~n785 & n5094 ) | ( n5017 & n5094 ) ;
  assign n5097 = n5051 | n5057 ;
  assign n5098 = ( ~n716 & n4985 ) | ( ~n716 & n5096 ) | ( n4985 & n5096 ) ;
  assign n5099 = ( ~n640 & n5020 ) | ( ~n640 & n5098 ) | ( n5020 & n5098 ) ;
  assign n5100 = n5087 ^ n1220 ^ 1'b0 ;
  assign n5101 = ( x53 & x54 ) | ( x53 & ~n5066 ) | ( x54 & ~n5066 ) ;
  assign n5102 = ( x55 & ~n5066 ) | ( x55 & n5101 ) | ( ~n5066 & n5101 ) ;
  assign n5103 = n5066 | n5068 ;
  assign n5104 = n5099 ^ n572 ^ 1'b0 ;
  assign n5105 = ( n4912 & n5095 ) | ( n4912 & ~n5103 ) | ( n5095 & ~n5103 ) ;
  assign n5106 = ( ~n572 & n4988 ) | ( ~n572 & n5099 ) | ( n4988 & n5099 ) ;
  assign n5107 = ( ~n514 & n4992 ) | ( ~n514 & n5106 ) | ( n4992 & n5106 ) ;
  assign n5108 = ( ~n458 & n4950 ) | ( ~n458 & n5107 ) | ( n4950 & n5107 ) ;
  assign n5109 = ( ~n399 & n5023 ) | ( ~n399 & n5108 ) | ( n5023 & n5108 ) ;
  assign n5110 = ( ~n345 & n5026 ) | ( ~n345 & n5109 ) | ( n5026 & n5109 ) ;
  assign n5111 = ( ~n302 & n5032 ) | ( ~n302 & n5110 ) | ( n5032 & n5110 ) ;
  assign n5112 = ( ~n261 & n4995 ) | ( ~n261 & n5111 ) | ( n4995 & n5111 ) ;
  assign n5113 = ( ~n217 & n4953 ) | ( ~n217 & n5112 ) | ( n4953 & n5112 ) ;
  assign n5114 = ( ~n179 & n4998 ) | ( ~n179 & n5113 ) | ( n4998 & n5113 ) ;
  assign n5115 = ( ~n144 & n5035 ) | ( ~n144 & n5114 ) | ( n5035 & n5114 ) ;
  assign n5116 = ( ~n134 & n5037 ) | ( ~n134 & n5115 ) | ( n5037 & n5115 ) ;
  assign n5117 = ( ~n136 & n4918 ) | ( ~n136 & n5116 ) | ( n4918 & n5116 ) ;
  assign n5118 = n4918 & n5116 ;
  assign n5119 = ( n5102 & n5103 ) | ( n5102 & ~n5118 ) | ( n5103 & ~n5118 ) ;
  assign n5120 = ~n5103 & n5119 ;
  assign n5121 = n5095 | n5117 ;
  assign n5122 = ~n136 & n5121 ;
  assign n5123 = n5118 | n5122 ;
  assign n5124 = n5103 | n5123 ;
  assign n5125 = n5124 ^ n5115 ^ n134 ;
  assign n5126 = n5124 ^ n5098 ^ n640 ;
  assign n5127 = n5124 & n5126 ;
  assign n5128 = ~n5040 & n5124 ;
  assign n5129 = n5123 & ~n5128 ;
  assign n5130 = ( n5105 & n5128 ) | ( n5105 & ~n5129 ) | ( n5128 & ~n5129 ) ;
  assign n5131 = n5124 ^ n5106 ^ n514 ;
  assign n5132 = n5124 & n5125 ;
  assign n5133 = n5124 ^ n5059 ^ n4346 ;
  assign n5134 = n5132 ^ n5036 ^ n4851 ;
  assign n5135 = n5124 & n5131 ;
  assign n5136 = n5093 & n5124 ;
  assign n5137 = n5135 ^ n4991 ^ n4824 ;
  assign n5138 = n5104 & n5124 ;
  assign n5139 = n5071 & n5124 ;
  assign n5140 = n5136 ^ n5124 ^ n4969 ;
  assign n5141 = n5100 & n5124 ;
  assign n5142 = n5138 ^ n5124 ^ n4988 ;
  assign n5143 = n5097 & n5124 ;
  assign n5144 = n5141 ^ n5124 ^ n4989 ;
  assign n5145 = n5143 ^ n5124 ^ n5052 ;
  assign n5146 = n5092 & n5124 ;
  assign n5147 = n5127 ^ n5019 ^ n4821 ;
  assign n5148 = n5139 ^ n5124 ^ n4960 ;
  assign n5149 = n5146 ^ n5124 ^ n4963 ;
  assign n5150 = n5124 & n5133 ;
  assign n5151 = n5150 ^ n4920 ^ n4855 ;
  assign n5152 = n5124 ^ n5061 ^ n3986 ;
  assign n5153 = n5124 & n5152 ;
  assign n5154 = n5153 ^ n4922 ^ n4788 ;
  assign n5155 = n5124 ^ n5064 ^ n3464 ;
  assign n5156 = n5124 & n5155 ;
  assign n5157 = n5156 ^ n4925 ^ n4743 ;
  assign n5158 = n5124 ^ n5070 ^ n3141 ;
  assign n5159 = n5124 ^ n5074 ^ n2839 ;
  assign n5160 = n5124 & n5159 ;
  assign n5161 = n5160 ^ n4928 ^ n4751 ;
  assign n5162 = n5124 ^ n5076 ^ n2544 ;
  assign n5163 = n5124 & n5162 ;
  assign n5164 = n5163 ^ n5007 ^ n4803 ;
  assign n5165 = n5124 ^ n5078 ^ n2269 ;
  assign n5166 = n5124 & n5165 ;
  assign n5167 = n5166 ^ n4965 ^ n4806 ;
  assign n5168 = n5124 ^ n5086 ^ n1318 ;
  assign n5169 = n5124 & n5168 ;
  assign n5170 = n5124 & n5158 ;
  assign n5171 = n5170 ^ n5001 ^ n4748 ;
  assign n5172 = n5169 ^ n5029 ^ n4766 ;
  assign n5173 = n5124 ^ n5088 ^ n1118 ;
  assign n5174 = n5124 & n5173 ;
  assign n5175 = n5174 ^ n4943 ^ n4771 ;
  assign n5176 = n5124 ^ n5089 ^ n1034 ;
  assign n5177 = n5124 & n5176 ;
  assign n5178 = n5177 ^ n4946 ^ n4774 ;
  assign n5179 = n5124 ^ n5091 ^ n859 ;
  assign n5180 = n5124 & n5179 ;
  assign n5181 = n5180 ^ n4981 ^ n4818 ;
  assign n5182 = n5124 ^ n5075 ^ n2690 ;
  assign n5183 = n5124 & n5182 ;
  assign n5184 = n5183 ^ n4931 ^ n4800 ;
  assign n5185 = n5124 ^ n5094 ^ n785 ;
  assign n5186 = n5124 & n5185 ;
  assign n5187 = n5186 ^ n5016 ^ n4780 ;
  assign n5188 = n5124 ^ n5110 ^ n302 ;
  assign n5189 = n5124 & n5188 ;
  assign n5190 = n5189 ^ n5031 ^ n4836 ;
  assign n5191 = n5096 ^ n716 ^ 1'b0 ;
  assign n5192 = n5124 & n5191 ;
  assign n5193 = n5192 ^ n5124 ^ n4985 ;
  assign n5194 = n5130 ^ x59 ^ 1'b0 ;
  assign n5195 = n5124 ^ n5109 ^ n345 ;
  assign n5196 = n5124 ^ n5062 ^ n3804 ;
  assign n5197 = n5124 ^ n5082 ^ n1766 ;
  assign n5198 = n5063 ^ n3631 ^ 1'b0 ;
  assign n5199 = n5124 ^ n5107 ^ n458 ;
  assign n5200 = n5124 ^ n5081 ^ n1885 ;
  assign n5201 = n5124 ^ n5083 ^ n1652 ;
  assign n5202 = n5124 ^ n5108 ^ n399 ;
  assign n5203 = n5124 ^ n5072 ^ n2995 ;
  assign n5204 = n5124 ^ n5058 ^ n4534 ;
  assign n5205 = n5124 ^ n5090 ^ n941 ;
  assign n5206 = n5124 ^ n5060 ^ n4167 ;
  assign n5207 = n5124 & n5206 ;
  assign n5208 = n5207 ^ n5039 ^ n4860 ;
  assign n5209 = n4918 & ~n5124 ;
  assign n5210 = n5111 ^ n261 ^ 1'b0 ;
  assign n5211 = n5124 & n5204 ;
  assign n5212 = n5211 ^ n5048 ^ x62 ;
  assign n5213 = n5124 & n5196 ;
  assign n5214 = n5213 ^ n4971 ^ n4791 ;
  assign n5215 = n5124 & n5210 ;
  assign n5216 = n5215 ^ n5124 ^ n4995 ;
  assign n5217 = n5124 & n5200 ;
  assign n5218 = n5217 ^ n4934 ^ n4758 ;
  assign n5219 = n5124 & n5203 ;
  assign n5220 = n5219 ^ n5004 ^ n4797 ;
  assign n5221 = n5124 & n5199 ;
  assign n5222 = n5124 ^ n5112 ^ n217 ;
  assign n5223 = n5124 & n5198 ;
  assign n5224 = n5223 ^ n5124 ^ n4957 ;
  assign n5225 = n5221 ^ n4949 ^ n4834 ;
  assign n5226 = n5124 ^ n5080 ^ n2009 ;
  assign n5227 = n5124 & n5197 ;
  assign n5228 = n5227 ^ n4937 ^ n4812 ;
  assign n5229 = n5124 & n5202 ;
  assign n5230 = n5229 ^ n5022 ^ n4829 ;
  assign n5231 = n5124 & n5205 ;
  assign n5232 = n5231 ^ n5013 ^ n4777 ;
  assign n5233 = n5124 ^ n5084 ^ n1534 ;
  assign n5234 = n5124 & n5222 ;
  assign n5235 = n5085 ^ n1416 ^ 1'b0 ;
  assign n5236 = n5234 ^ n4952 ^ n4842 ;
  assign n5237 = n5124 & n5233 ;
  assign n5238 = n5237 ^ n4973 ^ n4815 ;
  assign n5239 = n5124 & n5235 ;
  assign n5240 = n5239 ^ n5124 ^ n4977 ;
  assign n5241 = n5124 & n5201 ;
  assign n5242 = n5241 ^ n4940 ^ n4761 ;
  assign n5243 = n5124 & n5195 ;
  assign n5244 = n5243 ^ n5025 ^ n4832 ;
  assign n5245 = ( n5116 & n5117 ) | ( n5116 & n5124 ) | ( n5117 & n5124 ) ;
  assign n5246 = n4918 & ~n5245 ;
  assign n5247 = n4918 & ~n5116 ;
  assign n5248 = ( n4918 & ~n5116 ) | ( n4918 & n5124 ) | ( ~n5116 & n5124 ) ;
  assign n5249 = n5124 & n5226 ;
  assign n5250 = n5249 ^ n5010 ^ n4809 ;
  assign n5251 = n5124 ^ n5114 ^ n144 ;
  assign n5252 = ( n5134 & ~n5247 ) | ( n5134 & n5248 ) | ( ~n5247 & n5248 ) ;
  assign n5253 = n5246 ^ n5245 ^ n5117 ;
  assign n5254 = n5113 ^ n179 ^ 1'b0 ;
  assign n5255 = n5124 & n5254 ;
  assign n5256 = n5255 ^ n5124 ^ n4998 ;
  assign n5257 = n5124 & n5251 ;
  assign n5258 = n5257 ^ n5034 ^ n4848 ;
  assign n5259 = x57 & n5124 ;
  assign n5260 = x55 | x56 ;
  assign n5261 = x57 | n5260 ;
  assign n5262 = n5259 ^ n5124 ^ x58 ;
  assign n5263 = ( x57 & ~n4913 ) | ( x57 & n5260 ) | ( ~n4913 & n5260 ) ;
  assign n5264 = ( ~n4915 & n5259 ) | ( ~n4915 & n5263 ) | ( n5259 & n5263 ) ;
  assign n5265 = ~n5259 & n5264 ;
  assign n5266 = ( n4915 & n5259 ) | ( n4915 & ~n5261 ) | ( n5259 & ~n5261 ) ;
  assign n5267 = n5262 | n5265 ;
  assign n5268 = ~n5266 & n5267 ;
  assign n5269 = ( ~n4728 & n5194 ) | ( ~n4728 & n5268 ) | ( n5194 & n5268 ) ;
  assign n5270 = ( ~n4534 & n5145 ) | ( ~n4534 & n5269 ) | ( n5145 & n5269 ) ;
  assign n5271 = ( ~n4346 & n5212 ) | ( ~n4346 & n5270 ) | ( n5212 & n5270 ) ;
  assign n5272 = ( ~n4167 & n5151 ) | ( ~n4167 & n5271 ) | ( n5151 & n5271 ) ;
  assign n5273 = ( ~n3986 & n5208 ) | ( ~n3986 & n5272 ) | ( n5208 & n5272 ) ;
  assign n5274 = ( ~n3804 & n5154 ) | ( ~n3804 & n5273 ) | ( n5154 & n5273 ) ;
  assign n5275 = ( ~n3631 & n5214 ) | ( ~n3631 & n5274 ) | ( n5214 & n5274 ) ;
  assign n5276 = ( ~n3464 & n5224 ) | ( ~n3464 & n5275 ) | ( n5224 & n5275 ) ;
  assign n5277 = ( ~n3302 & n5157 ) | ( ~n3302 & n5276 ) | ( n5157 & n5276 ) ;
  assign n5278 = ( ~n3141 & n5148 ) | ( ~n3141 & n5277 ) | ( n5148 & n5277 ) ;
  assign n5279 = ( ~n2995 & n5171 ) | ( ~n2995 & n5278 ) | ( n5171 & n5278 ) ;
  assign n5280 = ( ~n2839 & n5220 ) | ( ~n2839 & n5279 ) | ( n5220 & n5279 ) ;
  assign n5281 = ( ~n2690 & n5161 ) | ( ~n2690 & n5280 ) | ( n5161 & n5280 ) ;
  assign n5282 = ( ~n2544 & n5184 ) | ( ~n2544 & n5281 ) | ( n5184 & n5281 ) ;
  assign n5283 = ( ~n2404 & n5164 ) | ( ~n2404 & n5282 ) | ( n5164 & n5282 ) ;
  assign n5284 = ( ~n2269 & n5149 ) | ( ~n2269 & n5283 ) | ( n5149 & n5283 ) ;
  assign n5285 = ( ~n2139 & n5167 ) | ( ~n2139 & n5284 ) | ( n5167 & n5284 ) ;
  assign n5286 = ( ~n2009 & n5140 ) | ( ~n2009 & n5285 ) | ( n5140 & n5285 ) ;
  assign n5287 = ( ~n1885 & n5250 ) | ( ~n1885 & n5286 ) | ( n5250 & n5286 ) ;
  assign n5288 = ( ~n1766 & n5218 ) | ( ~n1766 & n5287 ) | ( n5218 & n5287 ) ;
  assign n5289 = ( ~n1652 & n5228 ) | ( ~n1652 & n5288 ) | ( n5228 & n5288 ) ;
  assign n5290 = ( ~n1534 & n5242 ) | ( ~n1534 & n5289 ) | ( n5242 & n5289 ) ;
  assign n5291 = ( ~n1416 & n5238 ) | ( ~n1416 & n5290 ) | ( n5238 & n5290 ) ;
  assign n5292 = ( ~n1318 & n5240 ) | ( ~n1318 & n5291 ) | ( n5240 & n5291 ) ;
  assign n5293 = ( ~n1220 & n5172 ) | ( ~n1220 & n5292 ) | ( n5172 & n5292 ) ;
  assign n5294 = n5265 | n5266 ;
  assign n5295 = ( ~n1118 & n5144 ) | ( ~n1118 & n5293 ) | ( n5144 & n5293 ) ;
  assign n5296 = ( ~n1034 & n5175 ) | ( ~n1034 & n5295 ) | ( n5175 & n5295 ) ;
  assign n5297 = ( ~n941 & n5178 ) | ( ~n941 & n5296 ) | ( n5178 & n5296 ) ;
  assign n5298 = ( ~n859 & n5232 ) | ( ~n859 & n5297 ) | ( n5232 & n5297 ) ;
  assign n5299 = ( ~n785 & n5181 ) | ( ~n785 & n5298 ) | ( n5181 & n5298 ) ;
  assign n5300 = ( ~n716 & n5187 ) | ( ~n716 & n5299 ) | ( n5187 & n5299 ) ;
  assign n5301 = ( ~n640 & n5193 ) | ( ~n640 & n5300 ) | ( n5193 & n5300 ) ;
  assign n5302 = ( ~n572 & n5147 ) | ( ~n572 & n5301 ) | ( n5147 & n5301 ) ;
  assign n5303 = ( ~n514 & n5142 ) | ( ~n514 & n5302 ) | ( n5142 & n5302 ) ;
  assign n5304 = ( ~n458 & n5137 ) | ( ~n458 & n5303 ) | ( n5137 & n5303 ) ;
  assign n5305 = ( ~n399 & n5225 ) | ( ~n399 & n5304 ) | ( n5225 & n5304 ) ;
  assign n5306 = ( ~n345 & n5230 ) | ( ~n345 & n5305 ) | ( n5230 & n5305 ) ;
  assign n5307 = ( ~n302 & n5244 ) | ( ~n302 & n5306 ) | ( n5244 & n5306 ) ;
  assign n5308 = ( ~n261 & n5190 ) | ( ~n261 & n5307 ) | ( n5190 & n5307 ) ;
  assign n5309 = ( ~n217 & n5216 ) | ( ~n217 & n5308 ) | ( n5216 & n5308 ) ;
  assign n5310 = ( ~n179 & n5236 ) | ( ~n179 & n5309 ) | ( n5236 & n5309 ) ;
  assign n5311 = ( ~n144 & n5256 ) | ( ~n144 & n5310 ) | ( n5256 & n5310 ) ;
  assign n5312 = ( ~n134 & n5258 ) | ( ~n134 & n5311 ) | ( n5258 & n5311 ) ;
  assign n5313 = n5134 & n5312 ;
  assign n5314 = n5253 | n5313 ;
  assign n5315 = n5308 ^ n217 ^ 1'b0 ;
  assign n5316 = ( ~x30 & n5252 ) | ( ~x30 & n5312 ) | ( n5252 & n5312 ) ;
  assign n5317 = ~n136 & n5316 ;
  assign n5318 = n5314 | n5317 ;
  assign n5319 = n5209 | n5318 ;
  assign n5320 = n5294 & n5319 ;
  assign n5321 = n5315 & n5319 ;
  assign n5322 = n5320 ^ n5319 ^ n5262 ;
  assign n5323 = n5319 ^ n5311 ^ n134 ;
  assign n5324 = n5319 ^ n5307 ^ n261 ;
  assign n5325 = n5319 & n5324 ;
  assign n5326 = n5319 ^ n5305 ^ n345 ;
  assign n5327 = n5319 & n5326 ;
  assign n5328 = n5327 ^ n5229 ^ n5023 ;
  assign n5329 = n5325 ^ n5189 ^ n5032 ;
  assign n5330 = n5319 & n5323 ;
  assign n5331 = n5330 ^ n5257 ^ n5035 ;
  assign n5332 = n5319 ^ n5306 ^ n302 ;
  assign n5333 = n5319 & n5332 ;
  assign n5334 = n5333 ^ n5243 ^ n5026 ;
  assign n5335 = n5321 ^ n5319 ^ n5216 ;
  assign n5336 = n5319 ^ n5309 ^ n179 ;
  assign n5337 = n5319 & n5336 ;
  assign n5338 = n5337 ^ n5234 ^ n4953 ;
  assign n5339 = n5310 ^ n144 ^ 1'b0 ;
  assign n5340 = n5319 & n5339 ;
  assign n5341 = n5340 ^ n5319 ^ n5256 ;
  assign n5342 = n5319 ^ n5270 ^ n4346 ;
  assign n5343 = n5319 & n5342 ;
  assign n5344 = n5343 ^ n5211 ^ n5050 ;
  assign n5345 = n5319 ^ n5271 ^ n4167 ;
  assign n5346 = n5319 & n5345 ;
  assign n5347 = n5346 ^ n5150 ^ n5047 ;
  assign n5348 = n5319 ^ n5273 ^ n3804 ;
  assign n5349 = n5319 & n5348 ;
  assign n5350 = n5349 ^ n5153 ^ n4923 ;
  assign n5351 = n5319 ^ n5274 ^ n3631 ;
  assign n5352 = n5319 & n5351 ;
  assign n5353 = n5352 ^ n5213 ^ n4972 ;
  assign n5354 = n5319 ^ n5276 ^ n3302 ;
  assign n5355 = n5319 & n5354 ;
  assign n5356 = n5355 ^ n5156 ^ n4926 ;
  assign n5357 = n5319 ^ n5278 ^ n2995 ;
  assign n5358 = n5319 & n5357 ;
  assign n5359 = n5358 ^ n5170 ^ n5002 ;
  assign n5360 = n5319 ^ n5280 ^ n2690 ;
  assign n5361 = n5319 & n5360 ;
  assign n5362 = n5361 ^ n5160 ^ n4929 ;
  assign n5363 = n5319 ^ n5281 ^ n2544 ;
  assign n5364 = n5319 & n5363 ;
  assign n5365 = n5364 ^ n5183 ^ n4932 ;
  assign n5366 = n5319 ^ n5284 ^ n2139 ;
  assign n5367 = n5319 & n5366 ;
  assign n5368 = n5367 ^ n5166 ^ n4966 ;
  assign n5369 = n5319 ^ n5287 ^ n1766 ;
  assign n5370 = n5319 & n5369 ;
  assign n5371 = n5370 ^ n5217 ^ n4935 ;
  assign n5372 = n5319 ^ n5288 ^ n1652 ;
  assign n5373 = n5319 & n5372 ;
  assign n5374 = n5373 ^ n5227 ^ n4938 ;
  assign n5375 = n5319 ^ n5289 ^ n1534 ;
  assign n5376 = n5319 & n5375 ;
  assign n5377 = n5376 ^ n5241 ^ n4941 ;
  assign n5378 = n5319 ^ n5290 ^ n1416 ;
  assign n5379 = n5319 & n5378 ;
  assign n5380 = n5379 ^ n5237 ^ n4974 ;
  assign n5381 = n5291 ^ n1318 ^ 1'b0 ;
  assign n5382 = n5319 & n5381 ;
  assign n5383 = n5382 ^ n5319 ^ n5240 ;
  assign n5384 = n5319 ^ n5292 ^ n1220 ;
  assign n5385 = n5319 & n5384 ;
  assign n5386 = n5385 ^ n5169 ^ n5030 ;
  assign n5387 = n5293 ^ n1118 ^ 1'b0 ;
  assign n5388 = n5319 & n5387 ;
  assign n5389 = n5388 ^ n5319 ^ n5144 ;
  assign n5390 = n5319 ^ n5295 ^ n1034 ;
  assign n5391 = n5319 & n5390 ;
  assign n5392 = n5391 ^ n5174 ^ n4944 ;
  assign n5393 = n5319 ^ n5296 ^ n941 ;
  assign n5394 = n5319 & n5393 ;
  assign n5395 = n5394 ^ n5177 ^ n4947 ;
  assign n5396 = n5319 ^ n5297 ^ n859 ;
  assign n5397 = n5319 & n5396 ;
  assign n5398 = n5397 ^ n5231 ^ n5014 ;
  assign n5399 = n5319 ^ n5298 ^ n785 ;
  assign n5400 = n5319 & n5399 ;
  assign n5401 = n5400 ^ n5180 ^ n4982 ;
  assign n5402 = n5319 ^ n5299 ^ n716 ;
  assign n5403 = n5319 & n5402 ;
  assign n5404 = n5403 ^ n5186 ^ n5017 ;
  assign n5405 = n5319 ^ n5301 ^ n572 ;
  assign n5406 = n5319 & n5405 ;
  assign n5407 = n5406 ^ n5127 ^ n5020 ;
  assign n5408 = n5319 ^ n5304 ^ n399 ;
  assign n5409 = n5319 & n5408 ;
  assign n5410 = n5409 ^ n5221 ^ n4950 ;
  assign n5411 = n5260 & n5319 ;
  assign n5412 = n5319 ^ n5303 ^ n458 ;
  assign n5413 = n5319 ^ n5279 ^ n2839 ;
  assign n5414 = n5277 ^ n3141 ^ 1'b0 ;
  assign n5415 = n5285 ^ n2009 ^ 1'b0 ;
  assign n5416 = n5275 ^ n3464 ^ 1'b0 ;
  assign n5417 = n5319 & n5412 ;
  assign n5418 = n5417 ^ n5135 ^ n4992 ;
  assign n5419 = ( x55 & n5122 ) | ( x55 & n5319 ) | ( n5122 & n5319 ) ;
  assign n5420 = n5319 ^ n5282 ^ n2404 ;
  assign n5421 = ( n5120 & ~n5122 ) | ( n5120 & n5419 ) | ( ~n5122 & n5419 ) ;
  assign n5422 = ( ~n5134 & n5312 ) | ( ~n5134 & n5319 ) | ( n5312 & n5319 ) ;
  assign n5423 = n5319 & n5416 ;
  assign n5424 = n5423 ^ n5319 ^ n5224 ;
  assign n5425 = n5319 & n5420 ;
  assign n5426 = n5300 ^ n640 ^ 1'b0 ;
  assign n5427 = n5319 ^ n5286 ^ n1885 ;
  assign n5428 = ~n5419 & n5421 ;
  assign n5429 = n5209 | n5313 ;
  assign n5430 = ( n5312 & n5313 ) | ( n5312 & ~n5319 ) | ( n5313 & ~n5319 ) ;
  assign n5431 = n5319 & n5414 ;
  assign n5432 = ( x51 & x52 ) | ( x51 & ~n5209 ) | ( x52 & ~n5209 ) ;
  assign n5433 = ( x53 & ~n5209 ) | ( x53 & n5432 ) | ( ~n5209 & n5432 ) ;
  assign n5434 = n5425 ^ n5163 ^ n5008 ;
  assign n5435 = ~n5134 & n5312 ;
  assign n5436 = ( ~n5253 & n5429 ) | ( ~n5253 & n5433 ) | ( n5429 & n5433 ) ;
  assign n5437 = ( n136 & n5134 ) | ( n136 & n5312 ) | ( n5134 & n5312 ) ;
  assign n5438 = n5319 ^ n5272 ^ n3986 ;
  assign n5439 = n5269 ^ n4534 ^ 1'b0 ;
  assign n5440 = n5319 & n5415 ;
  assign n5441 = n5283 ^ n2269 ^ 1'b0 ;
  assign n5442 = n5440 ^ n5319 ^ n5140 ;
  assign n5443 = n5124 & ~n5318 ;
  assign n5444 = n5431 ^ n5319 ^ n5148 ;
  assign n5445 = ( n5134 & ~n5209 ) | ( n5134 & n5253 ) | ( ~n5209 & n5253 ) ;
  assign n5446 = ~n5318 & n5445 ;
  assign n5447 = ( n5331 & n5422 ) | ( n5331 & ~n5435 ) | ( n5422 & ~n5435 ) ;
  assign n5448 = ~n5429 & n5436 ;
  assign n5449 = n5319 & n5441 ;
  assign n5450 = n5319 & n5438 ;
  assign n5451 = n5449 ^ n5319 ^ n5149 ;
  assign n5452 = n5319 ^ n5268 ^ n4728 ;
  assign n5453 = n5302 ^ n514 ^ 1'b0 ;
  assign n5454 = ( n5319 & ~n5411 ) | ( n5319 & n5443 ) | ( ~n5411 & n5443 ) ;
  assign n5455 = n5319 & n5413 ;
  assign n5456 = n5319 & n5439 ;
  assign n5457 = n5456 ^ n5319 ^ n5145 ;
  assign n5458 = n5455 ^ n5219 ^ n5005 ;
  assign n5459 = n5319 & n5452 ;
  assign n5460 = n5319 & n5427 ;
  assign n5461 = n5459 ^ n5130 ^ x59 ;
  assign n5462 = n5319 & n5426 ;
  assign n5463 = ~n5430 & n5437 ;
  assign n5464 = n5462 ^ n5319 ^ n5193 ;
  assign n5465 = n5460 ^ n5249 ^ n5011 ;
  assign n5466 = n5319 & n5453 ;
  assign n5467 = n5466 ^ n5319 ^ n5142 ;
  assign n5468 = n5450 ^ n5207 ^ n5044 ;
  assign n5469 = n5454 ^ x57 ^ 1'b0 ;
  assign n5470 = x53 | x54 ;
  assign n5471 = ( x55 & n5124 ) | ( x55 & ~n5470 ) | ( n5124 & ~n5470 ) ;
  assign n5472 = ( ~x55 & n5124 ) | ( ~x55 & n5319 ) | ( n5124 & n5319 ) ;
  assign n5473 = n5471 & n5472 ;
  assign n5474 = ~x55 & n5319 ;
  assign n5475 = n5474 ^ x56 ^ 1'b0 ;
  assign n5476 = n5428 | n5475 ;
  assign n5477 = ~n5473 & n5476 ;
  assign n5478 = ( ~n4915 & n5469 ) | ( ~n4915 & n5477 ) | ( n5469 & n5477 ) ;
  assign n5479 = ( ~n4728 & n5322 ) | ( ~n4728 & n5478 ) | ( n5322 & n5478 ) ;
  assign n5480 = ( ~n4534 & n5461 ) | ( ~n4534 & n5479 ) | ( n5461 & n5479 ) ;
  assign n5481 = ( ~n4346 & n5457 ) | ( ~n4346 & n5480 ) | ( n5457 & n5480 ) ;
  assign n5482 = ( ~n4167 & n5344 ) | ( ~n4167 & n5481 ) | ( n5344 & n5481 ) ;
  assign n5483 = ( ~n3986 & n5347 ) | ( ~n3986 & n5482 ) | ( n5347 & n5482 ) ;
  assign n5484 = ( ~n3804 & n5468 ) | ( ~n3804 & n5483 ) | ( n5468 & n5483 ) ;
  assign n5485 = ( ~n3631 & n5350 ) | ( ~n3631 & n5484 ) | ( n5350 & n5484 ) ;
  assign n5486 = ( ~n3464 & n5353 ) | ( ~n3464 & n5485 ) | ( n5353 & n5485 ) ;
  assign n5487 = ( ~n3302 & n5424 ) | ( ~n3302 & n5486 ) | ( n5424 & n5486 ) ;
  assign n5488 = ( ~n3141 & n5356 ) | ( ~n3141 & n5487 ) | ( n5356 & n5487 ) ;
  assign n5489 = ( ~n2995 & n5444 ) | ( ~n2995 & n5488 ) | ( n5444 & n5488 ) ;
  assign n5490 = ( ~n2839 & n5359 ) | ( ~n2839 & n5489 ) | ( n5359 & n5489 ) ;
  assign n5491 = ( ~n2690 & n5458 ) | ( ~n2690 & n5490 ) | ( n5458 & n5490 ) ;
  assign n5492 = ( ~n2544 & n5362 ) | ( ~n2544 & n5491 ) | ( n5362 & n5491 ) ;
  assign n5493 = ( ~n2404 & n5365 ) | ( ~n2404 & n5492 ) | ( n5365 & n5492 ) ;
  assign n5494 = ( ~n2269 & n5434 ) | ( ~n2269 & n5493 ) | ( n5434 & n5493 ) ;
  assign n5495 = ( ~n2139 & n5451 ) | ( ~n2139 & n5494 ) | ( n5451 & n5494 ) ;
  assign n5496 = ( ~n2009 & n5368 ) | ( ~n2009 & n5495 ) | ( n5368 & n5495 ) ;
  assign n5497 = ( ~n1885 & n5442 ) | ( ~n1885 & n5496 ) | ( n5442 & n5496 ) ;
  assign n5498 = ( ~n1766 & n5465 ) | ( ~n1766 & n5497 ) | ( n5465 & n5497 ) ;
  assign n5499 = ( ~n1652 & n5371 ) | ( ~n1652 & n5498 ) | ( n5371 & n5498 ) ;
  assign n5500 = ( ~n1534 & n5374 ) | ( ~n1534 & n5499 ) | ( n5374 & n5499 ) ;
  assign n5501 = ( ~n1416 & n5377 ) | ( ~n1416 & n5500 ) | ( n5377 & n5500 ) ;
  assign n5502 = ( ~n1318 & n5380 ) | ( ~n1318 & n5501 ) | ( n5380 & n5501 ) ;
  assign n5503 = ( ~n1220 & n5383 ) | ( ~n1220 & n5502 ) | ( n5383 & n5502 ) ;
  assign n5504 = ( ~n1118 & n5386 ) | ( ~n1118 & n5503 ) | ( n5386 & n5503 ) ;
  assign n5505 = ( ~n1034 & n5389 ) | ( ~n1034 & n5504 ) | ( n5389 & n5504 ) ;
  assign n5506 = ( ~n941 & n5392 ) | ( ~n941 & n5505 ) | ( n5392 & n5505 ) ;
  assign n5507 = ( ~n859 & n5395 ) | ( ~n859 & n5506 ) | ( n5395 & n5506 ) ;
  assign n5508 = ( ~n785 & n5398 ) | ( ~n785 & n5507 ) | ( n5398 & n5507 ) ;
  assign n5509 = ( ~n716 & n5401 ) | ( ~n716 & n5508 ) | ( n5401 & n5508 ) ;
  assign n5510 = ( ~n640 & n5404 ) | ( ~n640 & n5509 ) | ( n5404 & n5509 ) ;
  assign n5511 = ( ~n572 & n5464 ) | ( ~n572 & n5510 ) | ( n5464 & n5510 ) ;
  assign n5512 = ( ~n514 & n5407 ) | ( ~n514 & n5511 ) | ( n5407 & n5511 ) ;
  assign n5513 = ( ~n458 & n5467 ) | ( ~n458 & n5512 ) | ( n5467 & n5512 ) ;
  assign n5514 = ( ~n399 & n5418 ) | ( ~n399 & n5513 ) | ( n5418 & n5513 ) ;
  assign n5515 = ( ~n345 & n5410 ) | ( ~n345 & n5514 ) | ( n5410 & n5514 ) ;
  assign n5516 = ( ~n302 & n5328 ) | ( ~n302 & n5515 ) | ( n5328 & n5515 ) ;
  assign n5517 = ( ~n261 & n5334 ) | ( ~n261 & n5516 ) | ( n5334 & n5516 ) ;
  assign n5518 = ( ~n217 & n5329 ) | ( ~n217 & n5517 ) | ( n5329 & n5517 ) ;
  assign n5519 = ( ~n179 & n5335 ) | ( ~n179 & n5518 ) | ( n5335 & n5518 ) ;
  assign n5520 = ( ~n144 & n5338 ) | ( ~n144 & n5519 ) | ( n5338 & n5519 ) ;
  assign n5521 = ( ~n134 & n5341 ) | ( ~n134 & n5520 ) | ( n5341 & n5520 ) ;
  assign n5522 = ( ~x30 & n5447 ) | ( ~x30 & n5521 ) | ( n5447 & n5521 ) ;
  assign n5523 = n5331 & n5521 ;
  assign n5524 = ~n136 & n5522 ;
  assign n5525 = n5523 | n5524 ;
  assign n5526 = n5463 | n5525 ;
  assign n5527 = n5446 | n5526 ;
  assign n5528 = n5527 ^ n5501 ^ n1318 ;
  assign n5529 = n5527 ^ n5493 ^ n2269 ;
  assign n5530 = n5527 & n5529 ;
  assign n5531 = n5527 ^ n5487 ^ n3141 ;
  assign n5532 = n5527 ^ n5497 ^ n1766 ;
  assign n5533 = ( n5428 & ~n5473 ) | ( n5428 & n5527 ) | ( ~n5473 & n5527 ) ;
  assign n5534 = n5530 ^ n5425 ^ n5164 ;
  assign n5535 = n5527 ^ n5492 ^ n2404 ;
  assign n5536 = n5527 & n5535 ;
  assign n5537 = ~n5428 & n5533 ;
  assign n5538 = n5527 ^ n5499 ^ n1534 ;
  assign n5539 = n5536 ^ n5364 ^ n5184 ;
  assign n5540 = n5527 ^ n5498 ^ n1652 ;
  assign n5541 = n5527 ^ n5505 ^ n941 ;
  assign n5542 = n5527 & n5532 ;
  assign n5543 = n5527 & n5531 ;
  assign n5544 = n5543 ^ n5355 ^ n5157 ;
  assign n5545 = ~n5470 & n5527 ;
  assign n5546 = n5527 & n5540 ;
  assign n5547 = ( n5446 & n5463 ) | ( n5446 & ~n5545 ) | ( n5463 & ~n5545 ) ;
  assign n5548 = n5542 ^ n5460 ^ n5250 ;
  assign n5549 = n5527 & n5538 ;
  assign n5550 = n5549 ^ n5373 ^ n5228 ;
  assign n5551 = n5546 ^ n5370 ^ n5218 ;
  assign n5552 = n5527 ^ n5500 ^ n1416 ;
  assign n5553 = n5527 & n5528 ;
  assign n5554 = n5553 ^ n5379 ^ n5238 ;
  assign n5555 = n5527 ^ n5490 ^ n2690 ;
  assign n5556 = n5527 & n5555 ;
  assign n5557 = n5527 ^ n5491 ^ n2544 ;
  assign n5558 = n5527 & n5557 ;
  assign n5559 = n5558 ^ n5361 ^ n5161 ;
  assign n5560 = n5527 & n5552 ;
  assign n5561 = n5560 ^ n5376 ^ n5242 ;
  assign n5562 = n5556 ^ n5455 ^ n5220 ;
  assign n5563 = n5527 & n5541 ;
  assign n5564 = n5563 ^ n5391 ^ n5175 ;
  assign n5565 = n5527 ^ n5508 ^ n716 ;
  assign n5566 = n5527 & n5565 ;
  assign n5567 = n5566 ^ n5400 ^ n5181 ;
  assign n5568 = n5527 ^ n5511 ^ n514 ;
  assign n5569 = n5527 & n5568 ;
  assign n5570 = n5569 ^ n5406 ^ n5147 ;
  assign n5571 = n5527 ^ n5513 ^ n399 ;
  assign n5572 = n5527 & n5571 ;
  assign n5573 = n5572 ^ n5417 ^ n5137 ;
  assign n5574 = n5478 ^ n4728 ^ 1'b0 ;
  assign n5575 = n5527 & n5574 ;
  assign n5576 = n5575 ^ n5527 ^ n5322 ;
  assign n5577 = n5480 ^ n4346 ^ 1'b0 ;
  assign n5578 = n5527 & n5577 ;
  assign n5579 = n5578 ^ n5527 ^ n5457 ;
  assign n5580 = n5527 ^ n5482 ^ n3986 ;
  assign n5581 = n5527 & n5580 ;
  assign n5582 = n5581 ^ n5346 ^ n5151 ;
  assign n5583 = n5486 ^ n3302 ^ 1'b0 ;
  assign n5584 = n5527 & n5583 ;
  assign n5585 = n5584 ^ n5527 ^ n5424 ;
  assign n5586 = n5488 ^ n2995 ^ 1'b0 ;
  assign n5587 = n5527 & n5586 ;
  assign n5588 = n5527 ^ n5489 ^ n2839 ;
  assign n5589 = n5527 & n5588 ;
  assign n5590 = n5589 ^ n5358 ^ n5171 ;
  assign n5591 = n5494 ^ n2139 ^ 1'b0 ;
  assign n5592 = n5527 & n5591 ;
  assign n5593 = n5592 ^ n5527 ^ n5451 ;
  assign n5594 = n5496 ^ n1885 ^ 1'b0 ;
  assign n5595 = n5527 & n5594 ;
  assign n5596 = n5595 ^ n5527 ^ n5442 ;
  assign n5597 = n5502 ^ n1220 ^ 1'b0 ;
  assign n5598 = n5527 & n5597 ;
  assign n5599 = n5598 ^ n5527 ^ n5383 ;
  assign n5600 = n5504 ^ n1034 ^ 1'b0 ;
  assign n5601 = n5527 & n5600 ;
  assign n5602 = n5601 ^ n5527 ^ n5389 ;
  assign n5603 = n5527 ^ n5479 ^ n4534 ;
  assign n5604 = n5527 & n5603 ;
  assign n5605 = n5604 ^ n5459 ^ n5194 ;
  assign n5606 = n5527 ^ n5507 ^ n785 ;
  assign n5607 = n5527 & n5606 ;
  assign n5608 = n5587 ^ n5527 ^ n5444 ;
  assign n5609 = n5607 ^ n5397 ^ n5232 ;
  assign n5610 = n5512 ^ n458 ^ 1'b0 ;
  assign n5611 = n5527 & n5610 ;
  assign n5612 = n5611 ^ n5527 ^ n5467 ;
  assign n5613 = n5527 ^ n5515 ^ n302 ;
  assign n5614 = n5527 & n5613 ;
  assign n5615 = n5614 ^ n5327 ^ n5230 ;
  assign n5616 = n5518 ^ n179 ^ 1'b0 ;
  assign n5617 = n5527 & n5616 ;
  assign n5618 = n5617 ^ n5527 ^ n5335 ;
  assign n5619 = n5520 ^ n134 ^ 1'b0 ;
  assign n5620 = n5527 & n5619 ;
  assign n5621 = n5620 ^ n5527 ^ n5341 ;
  assign n5622 = n5527 ^ n5481 ^ n4167 ;
  assign n5623 = n5527 ^ n5503 ^ n1118 ;
  assign n5624 = n5527 & n5622 ;
  assign n5625 = n5527 ^ n5519 ^ n144 ;
  assign n5626 = n5624 ^ n5343 ^ n5212 ;
  assign n5627 = n5527 ^ n5495 ^ n2009 ;
  assign n5628 = n5527 ^ n5483 ^ n3804 ;
  assign n5629 = n5527 ^ n5484 ^ n3631 ;
  assign n5630 = n5319 & ~n5525 ;
  assign n5631 = n5527 ^ n5485 ^ n3464 ;
  assign n5632 = n5527 & n5629 ;
  assign n5633 = n5527 ^ n5506 ^ n859 ;
  assign n5634 = n5527 ^ n5514 ^ n345 ;
  assign n5635 = n5527 ^ n5516 ^ n261 ;
  assign n5636 = n5632 ^ n5349 ^ n5154 ;
  assign n5637 = ( x53 & n5317 ) | ( x53 & n5527 ) | ( n5317 & n5527 ) ;
  assign n5638 = ( ~n5317 & n5448 ) | ( ~n5317 & n5637 ) | ( n5448 & n5637 ) ;
  assign n5639 = n5527 ^ n5517 ^ n217 ;
  assign n5640 = n5527 & n5634 ;
  assign n5641 = n5527 & n5627 ;
  assign n5642 = n5640 ^ n5409 ^ n5225 ;
  assign n5643 = n5527 & n5623 ;
  assign n5644 = n5641 ^ n5367 ^ n5167 ;
  assign n5645 = n5545 | n5630 ;
  assign n5646 = n5527 & n5631 ;
  assign n5647 = n5646 ^ n5352 ^ n5214 ;
  assign n5648 = n5643 ^ n5385 ^ n5172 ;
  assign n5649 = n5527 & n5633 ;
  assign n5650 = n5527 & n5625 ;
  assign n5651 = n5527 & n5635 ;
  assign n5652 = n5650 ^ n5337 ^ n5236 ;
  assign n5653 = n5649 ^ n5394 ^ n5178 ;
  assign n5654 = n5527 & n5639 ;
  assign n5655 = n5654 ^ n5325 ^ n5190 ;
  assign n5656 = ( n5545 & ~n5547 ) | ( n5545 & n5645 ) | ( ~n5547 & n5645 ) ;
  assign n5657 = n5527 & n5628 ;
  assign n5658 = ~n5637 & n5638 ;
  assign n5659 = n5651 ^ n5333 ^ n5244 ;
  assign n5660 = n5657 ^ n5450 ^ n5208 ;
  assign n5661 = x51 | x52 ;
  assign n5662 = ( x53 & n5319 ) | ( x53 & ~n5661 ) | ( n5319 & ~n5661 ) ;
  assign n5663 = n4915 & n5477 ;
  assign n5664 = ~x53 & n5527 ;
  assign n5665 = n5664 ^ x54 ^ 1'b0 ;
  assign n5666 = n5658 | n5665 ;
  assign n5667 = n5527 ^ n5509 ^ n640 ;
  assign n5668 = n5527 & n5667 ;
  assign n5669 = n5510 ^ n572 ^ 1'b0 ;
  assign n5670 = n5656 ^ x55 ^ 1'b0 ;
  assign n5671 = ( n5521 & n5523 ) | ( n5521 & ~n5527 ) | ( n5523 & ~n5527 ) ;
  assign n5672 = ( ~x53 & n5319 ) | ( ~x53 & n5527 ) | ( n5319 & n5527 ) ;
  assign n5673 = n5662 & n5672 ;
  assign n5674 = n5666 & ~n5673 ;
  assign n5675 = ( ~n4915 & n5527 ) | ( ~n4915 & n5663 ) | ( n5527 & n5663 ) ;
  assign n5676 = ( ~n5124 & n5670 ) | ( ~n5124 & n5674 ) | ( n5670 & n5674 ) ;
  assign n5677 = n5537 ^ n5474 ^ x56 ;
  assign n5678 = ( ~n4915 & n5676 ) | ( ~n4915 & n5677 ) | ( n5676 & n5677 ) ;
  assign n5679 = ( ~n5477 & n5663 ) | ( ~n5477 & n5675 ) | ( n5663 & n5675 ) ;
  assign n5680 = n5679 ^ n5454 ^ x57 ;
  assign n5681 = ( ~n4728 & n5678 ) | ( ~n4728 & n5680 ) | ( n5678 & n5680 ) ;
  assign n5682 = ( ~n4534 & n5576 ) | ( ~n4534 & n5681 ) | ( n5576 & n5681 ) ;
  assign n5683 = ( ~n4346 & n5605 ) | ( ~n4346 & n5682 ) | ( n5605 & n5682 ) ;
  assign n5684 = ( n5331 & ~n5521 ) | ( n5331 & n5527 ) | ( ~n5521 & n5527 ) ;
  assign n5685 = n5527 & n5669 ;
  assign n5686 = ( n136 & n5331 ) | ( n136 & n5521 ) | ( n5331 & n5521 ) ;
  assign n5687 = ~n5671 & n5686 ;
  assign n5688 = n5668 ^ n5403 ^ n5187 ;
  assign n5689 = ( ~n4167 & n5579 ) | ( ~n4167 & n5683 ) | ( n5579 & n5683 ) ;
  assign n5690 = ( ~n3986 & n5626 ) | ( ~n3986 & n5689 ) | ( n5626 & n5689 ) ;
  assign n5691 = ( ~n3804 & n5582 ) | ( ~n3804 & n5690 ) | ( n5582 & n5690 ) ;
  assign n5692 = ( ~n3631 & n5660 ) | ( ~n3631 & n5691 ) | ( n5660 & n5691 ) ;
  assign n5693 = ( ~n3464 & n5636 ) | ( ~n3464 & n5692 ) | ( n5636 & n5692 ) ;
  assign n5694 = ( ~n3302 & n5647 ) | ( ~n3302 & n5693 ) | ( n5647 & n5693 ) ;
  assign n5695 = ( n5331 & ~n5527 ) | ( n5331 & n5687 ) | ( ~n5527 & n5687 ) ;
  assign n5696 = ( ~n3141 & n5585 ) | ( ~n3141 & n5694 ) | ( n5585 & n5694 ) ;
  assign n5697 = ( ~n2995 & n5544 ) | ( ~n2995 & n5696 ) | ( n5544 & n5696 ) ;
  assign n5698 = ( ~n2839 & n5608 ) | ( ~n2839 & n5697 ) | ( n5608 & n5697 ) ;
  assign n5699 = ( ~n2690 & n5590 ) | ( ~n2690 & n5698 ) | ( n5590 & n5698 ) ;
  assign n5700 = ( ~n2544 & n5562 ) | ( ~n2544 & n5699 ) | ( n5562 & n5699 ) ;
  assign n5701 = ( ~n2404 & n5559 ) | ( ~n2404 & n5700 ) | ( n5559 & n5700 ) ;
  assign n5702 = ( ~n2269 & n5539 ) | ( ~n2269 & n5701 ) | ( n5539 & n5701 ) ;
  assign n5703 = ( ~n2139 & n5534 ) | ( ~n2139 & n5702 ) | ( n5534 & n5702 ) ;
  assign n5704 = ( ~n2009 & n5593 ) | ( ~n2009 & n5703 ) | ( n5593 & n5703 ) ;
  assign n5705 = ( ~n1885 & n5644 ) | ( ~n1885 & n5704 ) | ( n5644 & n5704 ) ;
  assign n5706 = n5703 ^ n2009 ^ 1'b0 ;
  assign n5707 = ( ~n1766 & n5596 ) | ( ~n1766 & n5705 ) | ( n5596 & n5705 ) ;
  assign n5708 = ( ~n1652 & n5548 ) | ( ~n1652 & n5707 ) | ( n5548 & n5707 ) ;
  assign n5709 = ( ~n1534 & n5551 ) | ( ~n1534 & n5708 ) | ( n5551 & n5708 ) ;
  assign n5710 = ( ~n1416 & n5550 ) | ( ~n1416 & n5709 ) | ( n5550 & n5709 ) ;
  assign n5711 = ( ~n1318 & n5561 ) | ( ~n1318 & n5710 ) | ( n5561 & n5710 ) ;
  assign n5712 = ( ~n1220 & n5554 ) | ( ~n1220 & n5711 ) | ( n5554 & n5711 ) ;
  assign n5713 = ( ~n1118 & n5599 ) | ( ~n1118 & n5712 ) | ( n5599 & n5712 ) ;
  assign n5714 = ( ~n1034 & n5648 ) | ( ~n1034 & n5713 ) | ( n5648 & n5713 ) ;
  assign n5715 = ( ~n941 & n5602 ) | ( ~n941 & n5714 ) | ( n5602 & n5714 ) ;
  assign n5716 = ( ~n859 & n5564 ) | ( ~n859 & n5715 ) | ( n5564 & n5715 ) ;
  assign n5717 = n5331 & ~n5521 ;
  assign n5718 = ( n5621 & n5684 ) | ( n5621 & ~n5717 ) | ( n5684 & ~n5717 ) ;
  assign n5719 = ( ~n785 & n5653 ) | ( ~n785 & n5716 ) | ( n5653 & n5716 ) ;
  assign n5720 = n5712 ^ n1118 ^ 1'b0 ;
  assign n5721 = ( ~n716 & n5609 ) | ( ~n716 & n5719 ) | ( n5609 & n5719 ) ;
  assign n5722 = n5681 ^ n4534 ^ 1'b0 ;
  assign n5723 = n5694 ^ n3141 ^ 1'b0 ;
  assign n5724 = n5685 ^ n5527 ^ n5464 ;
  assign n5725 = ( ~n640 & n5567 ) | ( ~n640 & n5721 ) | ( n5567 & n5721 ) ;
  assign n5726 = n5697 ^ n2839 ^ 1'b0 ;
  assign n5727 = ( ~n572 & n5688 ) | ( ~n572 & n5725 ) | ( n5688 & n5725 ) ;
  assign n5728 = ( ~n514 & n5724 ) | ( ~n514 & n5727 ) | ( n5724 & n5727 ) ;
  assign n5729 = ( ~n458 & n5570 ) | ( ~n458 & n5728 ) | ( n5570 & n5728 ) ;
  assign n5730 = ( ~n399 & n5612 ) | ( ~n399 & n5729 ) | ( n5612 & n5729 ) ;
  assign n5731 = ( ~n345 & n5573 ) | ( ~n345 & n5730 ) | ( n5573 & n5730 ) ;
  assign n5732 = ( ~n302 & n5642 ) | ( ~n302 & n5731 ) | ( n5642 & n5731 ) ;
  assign n5733 = ( ~n261 & n5615 ) | ( ~n261 & n5732 ) | ( n5615 & n5732 ) ;
  assign n5734 = ( ~n217 & n5659 ) | ( ~n217 & n5733 ) | ( n5659 & n5733 ) ;
  assign n5735 = ( ~n179 & n5655 ) | ( ~n179 & n5734 ) | ( n5655 & n5734 ) ;
  assign n5736 = ( ~n144 & n5618 ) | ( ~n144 & n5735 ) | ( n5618 & n5735 ) ;
  assign n5737 = ( ~n134 & n5652 ) | ( ~n134 & n5736 ) | ( n5652 & n5736 ) ;
  assign n5738 = ( ~x30 & n5718 ) | ( ~x30 & n5737 ) | ( n5718 & n5737 ) ;
  assign n5739 = ~n136 & n5738 ;
  assign n5740 = ~n5621 & n5737 ;
  assign n5741 = ( n5737 & n5739 ) | ( n5737 & ~n5740 ) | ( n5739 & ~n5740 ) ;
  assign n5742 = n5687 | n5741 ;
  assign n5743 = n5695 | n5742 ;
  assign n5744 = n5743 ^ n5736 ^ n134 ;
  assign n5745 = n5743 & n5744 ;
  assign n5746 = n5745 ^ n5650 ^ n5338 ;
  assign n5747 = ( n5658 & ~n5673 ) | ( n5658 & n5743 ) | ( ~n5673 & n5743 ) ;
  assign n5748 = ~n5658 & n5747 ;
  assign n5749 = n5743 ^ n5676 ^ n4915 ;
  assign n5750 = n5743 & n5749 ;
  assign n5751 = n5750 ^ n5537 ^ n5475 ;
  assign n5752 = n5722 & n5743 ;
  assign n5753 = n5752 ^ n5743 ^ n5576 ;
  assign n5754 = n5723 & n5743 ;
  assign n5755 = n5754 ^ n5743 ^ n5585 ;
  assign n5756 = n5743 ^ n5696 ^ n2995 ;
  assign n5757 = n5743 & n5756 ;
  assign n5758 = n5757 ^ n5543 ^ n5356 ;
  assign n5759 = n5726 & n5743 ;
  assign n5760 = n5759 ^ n5743 ^ n5608 ;
  assign n5761 = n5743 ^ n5702 ^ n2139 ;
  assign n5762 = n5743 & n5761 ;
  assign n5763 = n5762 ^ n5530 ^ n5434 ;
  assign n5764 = n5706 & n5743 ;
  assign n5765 = n5764 ^ n5743 ^ n5593 ;
  assign n5766 = n5743 ^ n5707 ^ n1652 ;
  assign n5767 = n5743 & n5766 ;
  assign n5768 = n5767 ^ n5542 ^ n5465 ;
  assign n5769 = n5743 ^ n5710 ^ n1318 ;
  assign n5770 = n5743 & n5769 ;
  assign n5771 = n5770 ^ n5560 ^ n5377 ;
  assign n5772 = n5720 & n5743 ;
  assign n5773 = n5772 ^ n5743 ^ n5599 ;
  assign n5774 = n5743 ^ n5725 ^ n572 ;
  assign n5775 = n5743 & n5774 ;
  assign n5776 = n5775 ^ n5668 ^ n5404 ;
  assign n5777 = n5743 ^ n5734 ^ n179 ;
  assign n5778 = n5743 & n5777 ;
  assign n5779 = n5778 ^ n5654 ^ n5329 ;
  assign n5780 = n5743 ^ n5678 ^ n4728 ;
  assign n5781 = n5743 & n5780 ;
  assign n5782 = n5781 ^ n5679 ^ n5469 ;
  assign n5783 = n5743 ^ n5690 ^ n3804 ;
  assign n5784 = n5743 & n5783 ;
  assign n5785 = n5784 ^ n5581 ^ n5347 ;
  assign n5786 = n5743 ^ n5698 ^ n2690 ;
  assign n5787 = n5743 ^ n5700 ^ n2404 ;
  assign n5788 = n5743 & n5787 ;
  assign n5789 = n5788 ^ n5558 ^ n5362 ;
  assign n5790 = n5743 ^ n5711 ^ n1220 ;
  assign n5791 = n5743 & n5790 ;
  assign n5792 = n5791 ^ n5553 ^ n5380 ;
  assign n5793 = n5743 ^ n5713 ^ n1034 ;
  assign n5794 = n5743 & n5793 ;
  assign n5795 = n5794 ^ n5643 ^ n5386 ;
  assign n5796 = n5743 ^ n5715 ^ n859 ;
  assign n5797 = n5743 & n5796 ;
  assign n5798 = n5743 & n5786 ;
  assign n5799 = n5798 ^ n5589 ^ n5359 ;
  assign n5800 = n5797 ^ n5563 ^ n5392 ;
  assign n5801 = n5743 ^ n5716 ^ n785 ;
  assign n5802 = n5743 & n5801 ;
  assign n5803 = n5802 ^ n5649 ^ n5395 ;
  assign n5804 = n5743 ^ n5719 ^ n716 ;
  assign n5805 = n5743 & n5804 ;
  assign n5806 = n5805 ^ n5607 ^ n5398 ;
  assign n5807 = n5743 ^ n5728 ^ n458 ;
  assign n5808 = n5743 & n5807 ;
  assign n5809 = n5808 ^ n5569 ^ n5407 ;
  assign n5810 = n5743 ^ n5704 ^ n1885 ;
  assign n5811 = n5743 & n5810 ;
  assign n5812 = n5811 ^ n5641 ^ n5368 ;
  assign n5813 = n5743 ^ n5730 ^ n345 ;
  assign n5814 = n5743 & n5813 ;
  assign n5815 = n5814 ^ n5572 ^ n5418 ;
  assign n5816 = n5743 ^ n5733 ^ n217 ;
  assign n5817 = n5743 & n5816 ;
  assign n5818 = n5817 ^ n5651 ^ n5334 ;
  assign n5819 = ~n5661 & n5743 ;
  assign n5820 = n5527 & ~n5742 ;
  assign n5821 = n5819 | n5820 ;
  assign n5822 = n5748 ^ n5664 ^ x54 ;
  assign n5823 = n5743 ^ n5674 ^ n5124 ;
  assign n5824 = n5743 & n5823 ;
  assign n5825 = n5824 ^ n5656 ^ x55 ;
  assign n5826 = n5743 ^ n5682 ^ n4346 ;
  assign n5827 = n5743 & n5826 ;
  assign n5828 = n5827 ^ n5604 ^ n5461 ;
  assign n5829 = n5683 ^ n4167 ^ 1'b0 ;
  assign n5830 = n5743 & n5829 ;
  assign n5831 = n5830 ^ n5743 ^ n5579 ;
  assign n5832 = n5743 ^ n5689 ^ n3986 ;
  assign n5833 = n5743 & n5832 ;
  assign n5834 = n5833 ^ n5624 ^ n5344 ;
  assign n5835 = n5743 ^ n5691 ^ n3631 ;
  assign n5836 = n5743 & n5835 ;
  assign n5837 = n5836 ^ n5657 ^ n5468 ;
  assign n5838 = n5743 ^ n5692 ^ n3464 ;
  assign n5839 = n5743 & n5838 ;
  assign n5840 = n5839 ^ n5632 ^ n5350 ;
  assign n5841 = n5743 ^ n5693 ^ n3302 ;
  assign n5842 = n5743 & n5841 ;
  assign n5843 = n5743 ^ n5699 ^ n2544 ;
  assign n5844 = n5743 & n5843 ;
  assign n5845 = n5844 ^ n5556 ^ n5458 ;
  assign n5846 = n5842 ^ n5646 ^ n5353 ;
  assign n5847 = n5705 ^ n1766 ^ 1'b0 ;
  assign n5848 = n5743 & n5847 ;
  assign n5849 = n5848 ^ n5743 ^ n5596 ;
  assign n5850 = n5743 ^ n5708 ^ n1534 ;
  assign n5851 = n5743 & n5850 ;
  assign n5852 = n5851 ^ n5546 ^ n5371 ;
  assign n5853 = n5743 ^ n5709 ^ n1416 ;
  assign n5854 = n5743 & n5853 ;
  assign n5855 = n5854 ^ n5549 ^ n5374 ;
  assign n5856 = n5714 ^ n941 ^ 1'b0 ;
  assign n5857 = n5743 & n5856 ;
  assign n5858 = n5857 ^ n5743 ^ n5602 ;
  assign n5859 = n5743 ^ n5721 ^ n640 ;
  assign n5860 = n5743 & n5859 ;
  assign n5861 = n5860 ^ n5566 ^ n5401 ;
  assign n5862 = n5727 ^ n514 ^ 1'b0 ;
  assign n5863 = n5743 & n5862 ;
  assign n5864 = n5863 ^ n5743 ^ n5724 ;
  assign n5865 = n5729 ^ n399 ^ 1'b0 ;
  assign n5866 = n5743 & n5865 ;
  assign n5867 = n5866 ^ n5743 ^ n5612 ;
  assign n5868 = n5743 ^ n5701 ^ n2269 ;
  assign n5869 = n5743 & n5868 ;
  assign n5870 = n5869 ^ n5536 ^ n5365 ;
  assign n5871 = n5743 ^ n5731 ^ n302 ;
  assign n5872 = n5743 & n5871 ;
  assign n5873 = n5872 ^ n5640 ^ n5410 ;
  assign n5874 = n5743 ^ n5732 ^ n261 ;
  assign n5875 = n5743 & n5874 ;
  assign n5876 = n5875 ^ n5614 ^ n5328 ;
  assign n5877 = n5735 ^ n144 ^ 1'b0 ;
  assign n5878 = n5743 & n5877 ;
  assign n5879 = n5878 ^ n5743 ^ n5618 ;
  assign n5880 = n5737 ^ n5621 ^ 1'b0 ;
  assign n5881 = x48 | x49 ;
  assign n5882 = ( x51 & ~n5525 ) | ( x51 & n5881 ) | ( ~n5525 & n5881 ) ;
  assign n5883 = x51 & n5743 ;
  assign n5884 = ( ~n5527 & n5882 ) | ( ~n5527 & n5883 ) | ( n5882 & n5883 ) ;
  assign n5885 = ~n5883 & n5884 ;
  assign n5886 = n5883 ^ n5743 ^ x52 ;
  assign n5887 = n5621 & ~n5743 ;
  assign n5888 = n5885 | n5886 ;
  assign n5889 = x51 | n5881 ;
  assign n5890 = n5821 ^ x53 ^ 1'b0 ;
  assign n5891 = ( n5527 & n5883 ) | ( n5527 & ~n5889 ) | ( n5883 & ~n5889 ) ;
  assign n5892 = n5888 & ~n5891 ;
  assign n5893 = ( ~n5319 & n5890 ) | ( ~n5319 & n5892 ) | ( n5890 & n5892 ) ;
  assign n5894 = ( ~n5124 & n5822 ) | ( ~n5124 & n5893 ) | ( n5822 & n5893 ) ;
  assign n5895 = ( ~n4915 & n5825 ) | ( ~n4915 & n5894 ) | ( n5825 & n5894 ) ;
  assign n5896 = ( ~n4728 & n5751 ) | ( ~n4728 & n5895 ) | ( n5751 & n5895 ) ;
  assign n5897 = ( ~n4534 & n5782 ) | ( ~n4534 & n5896 ) | ( n5782 & n5896 ) ;
  assign n5898 = ( ~n4346 & n5753 ) | ( ~n4346 & n5897 ) | ( n5753 & n5897 ) ;
  assign n5899 = ( ~n4167 & n5828 ) | ( ~n4167 & n5898 ) | ( n5828 & n5898 ) ;
  assign n5900 = ( ~n3986 & n5831 ) | ( ~n3986 & n5899 ) | ( n5831 & n5899 ) ;
  assign n5901 = ( ~n3804 & n5834 ) | ( ~n3804 & n5900 ) | ( n5834 & n5900 ) ;
  assign n5902 = ( ~n3631 & n5785 ) | ( ~n3631 & n5901 ) | ( n5785 & n5901 ) ;
  assign n5903 = ( ~n3464 & n5837 ) | ( ~n3464 & n5902 ) | ( n5837 & n5902 ) ;
  assign n5904 = ( ~n3302 & n5840 ) | ( ~n3302 & n5903 ) | ( n5840 & n5903 ) ;
  assign n5905 = ( ~n3141 & n5846 ) | ( ~n3141 & n5904 ) | ( n5846 & n5904 ) ;
  assign n5906 = ( n136 & n5621 ) | ( n136 & n5737 ) | ( n5621 & n5737 ) ;
  assign n5907 = ( ~n2995 & n5755 ) | ( ~n2995 & n5905 ) | ( n5755 & n5905 ) ;
  assign n5908 = ( ~n2839 & n5758 ) | ( ~n2839 & n5907 ) | ( n5758 & n5907 ) ;
  assign n5909 = ( ~n2690 & n5760 ) | ( ~n2690 & n5908 ) | ( n5760 & n5908 ) ;
  assign n5910 = ( ~n2544 & n5799 ) | ( ~n2544 & n5909 ) | ( n5799 & n5909 ) ;
  assign n5911 = ( ~n2404 & n5845 ) | ( ~n2404 & n5910 ) | ( n5845 & n5910 ) ;
  assign n5912 = ( ~n2269 & n5789 ) | ( ~n2269 & n5911 ) | ( n5789 & n5911 ) ;
  assign n5913 = ( ~n2139 & n5870 ) | ( ~n2139 & n5912 ) | ( n5870 & n5912 ) ;
  assign n5914 = ( n5621 & n5737 ) | ( n5621 & ~n5743 ) | ( n5737 & ~n5743 ) ;
  assign n5915 = n5908 ^ n2690 ^ 1'b0 ;
  assign n5916 = ( ~n2009 & n5763 ) | ( ~n2009 & n5913 ) | ( n5763 & n5913 ) ;
  assign n5917 = n5905 ^ n2995 ^ 1'b0 ;
  assign n5918 = ( ~n1885 & n5765 ) | ( ~n1885 & n5916 ) | ( n5765 & n5916 ) ;
  assign n5919 = n5897 ^ n4346 ^ 1'b0 ;
  assign n5920 = ( ~n1766 & n5812 ) | ( ~n1766 & n5918 ) | ( n5812 & n5918 ) ;
  assign n5921 = n5920 ^ n1652 ^ 1'b0 ;
  assign n5922 = ( x44 & x45 ) | ( x44 & ~n5887 ) | ( x45 & ~n5887 ) ;
  assign n5923 = ( ~n1652 & n5849 ) | ( ~n1652 & n5920 ) | ( n5849 & n5920 ) ;
  assign n5924 = ( ~n1534 & n5768 ) | ( ~n1534 & n5923 ) | ( n5768 & n5923 ) ;
  assign n5925 = ( ~n1416 & n5852 ) | ( ~n1416 & n5924 ) | ( n5852 & n5924 ) ;
  assign n5926 = ( n5621 & ~n5737 ) | ( n5621 & n5743 ) | ( ~n5737 & n5743 ) ;
  assign n5927 = ( ~n1318 & n5855 ) | ( ~n1318 & n5925 ) | ( n5855 & n5925 ) ;
  assign n5928 = ( ~n1220 & n5771 ) | ( ~n1220 & n5927 ) | ( n5771 & n5927 ) ;
  assign n5929 = n5737 & n5914 ;
  assign n5930 = ( x46 & ~n5887 ) | ( x46 & n5922 ) | ( ~n5887 & n5922 ) ;
  assign n5931 = ( ~n1118 & n5792 ) | ( ~n1118 & n5928 ) | ( n5792 & n5928 ) ;
  assign n5932 = n5885 | n5891 ;
  assign n5933 = ( n5737 & ~n5880 ) | ( n5737 & n5926 ) | ( ~n5880 & n5926 ) ;
  assign n5934 = ( ~n1034 & n5773 ) | ( ~n1034 & n5931 ) | ( n5773 & n5931 ) ;
  assign n5935 = ( ~n941 & n5795 ) | ( ~n941 & n5934 ) | ( n5795 & n5934 ) ;
  assign n5936 = ( n5887 & n5906 ) | ( n5887 & ~n5929 ) | ( n5906 & ~n5929 ) ;
  assign n5937 = ( n5739 & n5933 ) | ( n5739 & ~n5936 ) | ( n5933 & ~n5936 ) ;
  assign n5938 = n5935 ^ n859 ^ 1'b0 ;
  assign n5939 = n5916 ^ n1885 ^ 1'b0 ;
  assign n5940 = n5931 ^ n1034 ^ 1'b0 ;
  assign n5941 = ( ~n859 & n5858 ) | ( ~n859 & n5935 ) | ( n5858 & n5935 ) ;
  assign n5942 = ( ~n785 & n5800 ) | ( ~n785 & n5941 ) | ( n5800 & n5941 ) ;
  assign n5943 = ( ~n716 & n5803 ) | ( ~n716 & n5942 ) | ( n5803 & n5942 ) ;
  assign n5944 = ( ~n640 & n5806 ) | ( ~n640 & n5943 ) | ( n5806 & n5943 ) ;
  assign n5945 = ( ~n572 & n5861 ) | ( ~n572 & n5944 ) | ( n5861 & n5944 ) ;
  assign n5946 = ( ~n514 & n5776 ) | ( ~n514 & n5945 ) | ( n5776 & n5945 ) ;
  assign n5947 = ( ~n458 & n5864 ) | ( ~n458 & n5946 ) | ( n5864 & n5946 ) ;
  assign n5948 = n5946 ^ n458 ^ 1'b0 ;
  assign n5949 = ( ~n399 & n5809 ) | ( ~n399 & n5947 ) | ( n5809 & n5947 ) ;
  assign n5950 = ( ~n345 & n5867 ) | ( ~n345 & n5949 ) | ( n5867 & n5949 ) ;
  assign n5951 = ( ~n302 & n5815 ) | ( ~n302 & n5950 ) | ( n5815 & n5950 ) ;
  assign n5952 = ( ~n261 & n5873 ) | ( ~n261 & n5951 ) | ( n5873 & n5951 ) ;
  assign n5953 = ( ~n217 & n5876 ) | ( ~n217 & n5952 ) | ( n5876 & n5952 ) ;
  assign n5954 = ( ~n179 & n5818 ) | ( ~n179 & n5953 ) | ( n5818 & n5953 ) ;
  assign n5955 = ( ~n144 & n5779 ) | ( ~n144 & n5954 ) | ( n5779 & n5954 ) ;
  assign n5956 = ( ~n134 & n5879 ) | ( ~n134 & n5955 ) | ( n5879 & n5955 ) ;
  assign n5957 = ( ~n136 & n5746 ) | ( ~n136 & n5956 ) | ( n5746 & n5956 ) ;
  assign n5958 = n5933 | n5957 ;
  assign n5959 = ~n136 & n5958 ;
  assign n5960 = n5746 & n5956 ;
  assign n5961 = ( n5930 & n5936 ) | ( n5930 & ~n5960 ) | ( n5936 & ~n5960 ) ;
  assign n5962 = ~n5936 & n5961 ;
  assign n5963 = n5959 | n5960 ;
  assign n5964 = n5936 | n5963 ;
  assign n5965 = n5948 & n5964 ;
  assign n5966 = n5940 & n5964 ;
  assign n5967 = n5966 ^ n5964 ^ n5773 ;
  assign n5968 = n5915 & n5964 ;
  assign n5969 = n5964 ^ n5944 ^ n572 ;
  assign n5970 = n5919 & n5964 ;
  assign n5971 = n5964 ^ n5934 ^ n941 ;
  assign n5972 = n5938 & n5964 ;
  assign n5973 = n5964 & n5971 ;
  assign n5974 = n5973 ^ n5794 ^ n5648 ;
  assign n5975 = n5964 & n5969 ;
  assign n5976 = n5975 ^ n5860 ^ n5567 ;
  assign n5977 = ~n5881 & n5964 ;
  assign n5978 = n5963 & ~n5977 ;
  assign n5979 = n5921 & n5964 ;
  assign n5980 = n5964 ^ n5923 ^ n1534 ;
  assign n5981 = n5964 & n5980 ;
  assign n5982 = n5917 & n5964 ;
  assign n5983 = n5981 ^ n5767 ^ n5548 ;
  assign n5984 = n5932 & n5964 ;
  assign n5985 = n5979 ^ n5964 ^ n5849 ;
  assign n5986 = n5939 & n5964 ;
  assign n5987 = n5965 ^ n5964 ^ n5864 ;
  assign n5988 = n5970 ^ n5964 ^ n5753 ;
  assign n5989 = n5968 ^ n5964 ^ n5760 ;
  assign n5990 = n5982 ^ n5964 ^ n5755 ;
  assign n5991 = n5986 ^ n5964 ^ n5765 ;
  assign n5992 = n5972 ^ n5964 ^ n5858 ;
  assign n5993 = n5984 ^ n5964 ^ n5886 ;
  assign n5994 = ( n5937 & n5977 ) | ( n5937 & ~n5978 ) | ( n5977 & ~n5978 ) ;
  assign n5995 = n5964 ^ n5895 ^ n4728 ;
  assign n5996 = n5964 & n5995 ;
  assign n5997 = n5996 ^ n5750 ^ n5677 ;
  assign n5998 = n5964 ^ n5896 ^ n4534 ;
  assign n5999 = n5964 & n5998 ;
  assign n6000 = n5999 ^ n5781 ^ n5680 ;
  assign n6001 = n5964 ^ n5898 ^ n4167 ;
  assign n6002 = n5964 ^ n5910 ^ n2404 ;
  assign n6003 = n5964 & n6002 ;
  assign n6004 = n6003 ^ n5844 ^ n5562 ;
  assign n6005 = n5964 ^ n5918 ^ n1766 ;
  assign n6006 = n5964 & n6005 ;
  assign n6007 = n6006 ^ n5811 ^ n5644 ;
  assign n6008 = n5964 ^ n5924 ^ n1416 ;
  assign n6009 = n5964 & n6008 ;
  assign n6010 = n6009 ^ n5851 ^ n5551 ;
  assign n6011 = n5964 ^ n5927 ^ n1220 ;
  assign n6012 = n5964 & n6011 ;
  assign n6013 = n5964 & n6001 ;
  assign n6014 = n6013 ^ n5827 ^ n5605 ;
  assign n6015 = n6012 ^ n5770 ^ n5561 ;
  assign n6016 = n5964 ^ n5943 ^ n640 ;
  assign n6017 = n5964 & n6016 ;
  assign n6018 = n6017 ^ n5805 ^ n5609 ;
  assign n6019 = n5964 ^ n5947 ^ n399 ;
  assign n6020 = n5964 & n6019 ;
  assign n6021 = n6020 ^ n5808 ^ n5570 ;
  assign n6022 = n5964 ^ n5950 ^ n302 ;
  assign n6023 = n5964 & n6022 ;
  assign n6024 = n6023 ^ n5814 ^ n5573 ;
  assign n6025 = n5964 ^ n5913 ^ n2009 ;
  assign n6026 = n5964 & n6025 ;
  assign n6027 = n6026 ^ n5762 ^ n5534 ;
  assign n6028 = n5964 ^ n5952 ^ n217 ;
  assign n6029 = n5964 & n6028 ;
  assign n6030 = n6029 ^ n5875 ^ n5615 ;
  assign n6031 = n5964 ^ n5953 ^ n179 ;
  assign n6032 = n5964 & n6031 ;
  assign n6033 = n6032 ^ n5817 ^ n5659 ;
  assign n6034 = n5899 ^ n3986 ^ 1'b0 ;
  assign n6035 = n5964 ^ n5903 ^ n3302 ;
  assign n6036 = n5964 ^ n5945 ^ n514 ;
  assign n6037 = n5949 ^ n345 ^ 1'b0 ;
  assign n6038 = n5964 & n6034 ;
  assign n6039 = n5964 & n6037 ;
  assign n6040 = n6039 ^ n5964 ^ n5867 ;
  assign n6041 = n5964 ^ n5941 ^ n785 ;
  assign n6042 = n5964 & n6041 ;
  assign n6043 = n6042 ^ n5797 ^ n5564 ;
  assign n6044 = n5964 ^ n5893 ^ n5124 ;
  assign n6045 = n5964 ^ n5942 ^ n716 ;
  assign n6046 = n5964 ^ n5902 ^ n3464 ;
  assign n6047 = n5964 ^ n5909 ^ n2544 ;
  assign n6048 = n5964 & n6047 ;
  assign n6049 = n5964 ^ n5901 ^ n3631 ;
  assign n6050 = n5964 & n6046 ;
  assign n6051 = ( n5746 & ~n5956 ) | ( n5746 & n5964 ) | ( ~n5956 & n5964 ) ;
  assign n6052 = n5964 ^ n5894 ^ n4915 ;
  assign n6053 = n5964 ^ n5907 ^ n2839 ;
  assign n6054 = n5964 ^ n5904 ^ n3141 ;
  assign n6055 = n5964 ^ n5892 ^ n5319 ;
  assign n6056 = n5964 & n6054 ;
  assign n6057 = n5746 & ~n5964 ;
  assign n6058 = n6050 ^ n5836 ^ n5660 ;
  assign n6059 = n5964 ^ n5925 ^ n1318 ;
  assign n6060 = n6048 ^ n5798 ^ n5590 ;
  assign n6061 = n5964 ^ n5900 ^ n3804 ;
  assign n6062 = n6056 ^ n5842 ^ n5647 ;
  assign n6063 = n5964 & n6055 ;
  assign n6064 = n5964 ^ n5911 ^ n2269 ;
  assign n6065 = n6063 ^ n5821 ^ x53 ;
  assign n6066 = n5964 & n6049 ;
  assign n6067 = n5964 ^ n5912 ^ n2139 ;
  assign n6068 = n6066 ^ n5784 ^ n5582 ;
  assign n6069 = n5964 & n6067 ;
  assign n6070 = n6069 ^ n5869 ^ n5539 ;
  assign n6071 = n5964 & n6053 ;
  assign n6072 = n6071 ^ n5757 ^ n5544 ;
  assign n6073 = n5964 & n6035 ;
  assign n6074 = n6073 ^ n5839 ^ n5636 ;
  assign n6075 = n5964 & n6061 ;
  assign n6076 = n6075 ^ n5833 ^ n5626 ;
  assign n6077 = n5964 & n6064 ;
  assign n6078 = n6077 ^ n5788 ^ n5559 ;
  assign n6079 = n5964 & n6044 ;
  assign n6080 = n6079 ^ n5748 ^ n5665 ;
  assign n6081 = n5964 & n6045 ;
  assign n6082 = n6081 ^ n5802 ^ n5653 ;
  assign n6083 = n5964 & n6052 ;
  assign n6084 = ( n5956 & n5957 ) | ( n5956 & n5964 ) | ( n5957 & n5964 ) ;
  assign n6085 = n5746 & ~n6084 ;
  assign n6086 = n5746 & ~n5956 ;
  assign n6087 = n5955 ^ n134 ^ 1'b0 ;
  assign n6088 = n5964 & n6087 ;
  assign n6089 = n5964 & n6036 ;
  assign n6090 = n6089 ^ n5775 ^ n5688 ;
  assign n6091 = n6088 ^ n5964 ^ n5879 ;
  assign n6092 = n6083 ^ n5824 ^ n5670 ;
  assign n6093 = ( n6051 & ~n6086 ) | ( n6051 & n6091 ) | ( ~n6086 & n6091 ) ;
  assign n6094 = n6085 ^ n6084 ^ n5957 ;
  assign n6095 = n6038 ^ n5964 ^ n5831 ;
  assign n6096 = n5964 ^ n5954 ^ n144 ;
  assign n6097 = n5964 & n6096 ;
  assign n6098 = n5964 ^ n5951 ^ n261 ;
  assign n6099 = n5964 & n6098 ;
  assign n6100 = n6097 ^ n5778 ^ n5655 ;
  assign n6101 = n5964 ^ n5928 ^ n1118 ;
  assign n6102 = n6099 ^ n5872 ^ n5642 ;
  assign n6103 = n5964 & n6101 ;
  assign n6104 = n5964 & n6059 ;
  assign n6105 = n6103 ^ n5791 ^ n5554 ;
  assign n6106 = n6104 ^ n5854 ^ n5550 ;
  assign n6107 = n5994 ^ x51 ^ 1'b0 ;
  assign n6108 = x48 & n5964 ;
  assign n6109 = x46 | x47 ;
  assign n6110 = x48 | n6109 ;
  assign n6111 = n6108 ^ n5964 ^ x49 ;
  assign n6112 = ( x48 & ~n5741 ) | ( x48 & n6109 ) | ( ~n5741 & n6109 ) ;
  assign n6113 = ( ~n5743 & n6108 ) | ( ~n5743 & n6112 ) | ( n6108 & n6112 ) ;
  assign n6114 = ( n5743 & n6108 ) | ( n5743 & ~n6110 ) | ( n6108 & ~n6110 ) ;
  assign n6115 = ~n6108 & n6113 ;
  assign n6116 = n6111 | n6115 ;
  assign n6117 = ~n6114 & n6116 ;
  assign n6118 = ( ~n5527 & n6107 ) | ( ~n5527 & n6117 ) | ( n6107 & n6117 ) ;
  assign n6119 = ( ~n5319 & n5993 ) | ( ~n5319 & n6118 ) | ( n5993 & n6118 ) ;
  assign n6120 = ( ~n5124 & n6065 ) | ( ~n5124 & n6119 ) | ( n6065 & n6119 ) ;
  assign n6121 = ( ~n4915 & n6080 ) | ( ~n4915 & n6120 ) | ( n6080 & n6120 ) ;
  assign n6122 = ( ~n4728 & n6092 ) | ( ~n4728 & n6121 ) | ( n6092 & n6121 ) ;
  assign n6123 = ( ~n4534 & n5997 ) | ( ~n4534 & n6122 ) | ( n5997 & n6122 ) ;
  assign n6124 = ( ~n4346 & n6000 ) | ( ~n4346 & n6123 ) | ( n6000 & n6123 ) ;
  assign n6125 = ( ~n4167 & n5988 ) | ( ~n4167 & n6124 ) | ( n5988 & n6124 ) ;
  assign n6126 = ( ~n3986 & n6014 ) | ( ~n3986 & n6125 ) | ( n6014 & n6125 ) ;
  assign n6127 = ( ~n3804 & n6095 ) | ( ~n3804 & n6126 ) | ( n6095 & n6126 ) ;
  assign n6128 = ( ~n3631 & n6076 ) | ( ~n3631 & n6127 ) | ( n6076 & n6127 ) ;
  assign n6129 = ( ~n3464 & n6068 ) | ( ~n3464 & n6128 ) | ( n6068 & n6128 ) ;
  assign n6130 = ( ~n3302 & n6058 ) | ( ~n3302 & n6129 ) | ( n6058 & n6129 ) ;
  assign n6131 = ( ~n3141 & n6074 ) | ( ~n3141 & n6130 ) | ( n6074 & n6130 ) ;
  assign n6132 = ( ~n2995 & n6062 ) | ( ~n2995 & n6131 ) | ( n6062 & n6131 ) ;
  assign n6133 = n6114 | n6115 ;
  assign n6134 = ( ~n2839 & n5990 ) | ( ~n2839 & n6132 ) | ( n5990 & n6132 ) ;
  assign n6135 = ( ~n2690 & n6072 ) | ( ~n2690 & n6134 ) | ( n6072 & n6134 ) ;
  assign n6136 = ( ~n2544 & n5989 ) | ( ~n2544 & n6135 ) | ( n5989 & n6135 ) ;
  assign n6137 = ( ~n2404 & n6060 ) | ( ~n2404 & n6136 ) | ( n6060 & n6136 ) ;
  assign n6138 = ( ~n2269 & n6004 ) | ( ~n2269 & n6137 ) | ( n6004 & n6137 ) ;
  assign n6139 = ( ~n2139 & n6078 ) | ( ~n2139 & n6138 ) | ( n6078 & n6138 ) ;
  assign n6140 = ( ~n2009 & n6070 ) | ( ~n2009 & n6139 ) | ( n6070 & n6139 ) ;
  assign n6141 = ( ~n1885 & n6027 ) | ( ~n1885 & n6140 ) | ( n6027 & n6140 ) ;
  assign n6142 = ( ~n1766 & n5991 ) | ( ~n1766 & n6141 ) | ( n5991 & n6141 ) ;
  assign n6143 = ( ~n1652 & n6007 ) | ( ~n1652 & n6142 ) | ( n6007 & n6142 ) ;
  assign n6144 = ( ~n1534 & n5985 ) | ( ~n1534 & n6143 ) | ( n5985 & n6143 ) ;
  assign n6145 = ( ~n1416 & n5983 ) | ( ~n1416 & n6144 ) | ( n5983 & n6144 ) ;
  assign n6146 = ( ~n1318 & n6010 ) | ( ~n1318 & n6145 ) | ( n6010 & n6145 ) ;
  assign n6147 = ( ~n1220 & n6106 ) | ( ~n1220 & n6146 ) | ( n6106 & n6146 ) ;
  assign n6148 = ( ~n1118 & n6015 ) | ( ~n1118 & n6147 ) | ( n6015 & n6147 ) ;
  assign n6149 = ( ~n1034 & n6105 ) | ( ~n1034 & n6148 ) | ( n6105 & n6148 ) ;
  assign n6150 = ( ~n941 & n5967 ) | ( ~n941 & n6149 ) | ( n5967 & n6149 ) ;
  assign n6151 = ( ~n859 & n5974 ) | ( ~n859 & n6150 ) | ( n5974 & n6150 ) ;
  assign n6152 = ( ~n785 & n5992 ) | ( ~n785 & n6151 ) | ( n5992 & n6151 ) ;
  assign n6153 = ( ~n716 & n6043 ) | ( ~n716 & n6152 ) | ( n6043 & n6152 ) ;
  assign n6154 = ( ~n640 & n6082 ) | ( ~n640 & n6153 ) | ( n6082 & n6153 ) ;
  assign n6155 = ( ~n572 & n6018 ) | ( ~n572 & n6154 ) | ( n6018 & n6154 ) ;
  assign n6156 = ( ~n514 & n5976 ) | ( ~n514 & n6155 ) | ( n5976 & n6155 ) ;
  assign n6157 = ( ~n458 & n6090 ) | ( ~n458 & n6156 ) | ( n6090 & n6156 ) ;
  assign n6158 = ( ~n399 & n5987 ) | ( ~n399 & n6157 ) | ( n5987 & n6157 ) ;
  assign n6159 = ( ~n345 & n6021 ) | ( ~n345 & n6158 ) | ( n6021 & n6158 ) ;
  assign n6160 = ( ~n302 & n6040 ) | ( ~n302 & n6159 ) | ( n6040 & n6159 ) ;
  assign n6161 = ( ~n261 & n6024 ) | ( ~n261 & n6160 ) | ( n6024 & n6160 ) ;
  assign n6162 = ( ~n217 & n6102 ) | ( ~n217 & n6161 ) | ( n6102 & n6161 ) ;
  assign n6163 = ( ~n179 & n6030 ) | ( ~n179 & n6162 ) | ( n6030 & n6162 ) ;
  assign n6164 = ( ~n144 & n6033 ) | ( ~n144 & n6163 ) | ( n6033 & n6163 ) ;
  assign n6165 = ( ~n134 & n6100 ) | ( ~n134 & n6164 ) | ( n6100 & n6164 ) ;
  assign n6166 = n6091 & n6165 ;
  assign n6167 = ( ~x30 & n6093 ) | ( ~x30 & n6165 ) | ( n6093 & n6165 ) ;
  assign n6168 = ~n136 & n6167 ;
  assign n6169 = n6057 | n6168 ;
  assign n6170 = n6166 | n6169 ;
  assign n6171 = n6094 | n6170 ;
  assign n6172 = n6171 ^ n6119 ^ n5124 ;
  assign n6173 = n6171 & n6172 ;
  assign n6174 = n6173 ^ n6063 ^ n5890 ;
  assign n6175 = n6133 & n6171 ;
  assign n6176 = n6175 ^ n6171 ^ n6111 ;
  assign n6177 = n6171 ^ n6127 ^ n3631 ;
  assign n6178 = n6171 & n6177 ;
  assign n6179 = n6178 ^ n6075 ^ n5834 ;
  assign n6180 = n6171 ^ n6128 ^ n3464 ;
  assign n6181 = n6171 & n6180 ;
  assign n6182 = n6181 ^ n6066 ^ n5785 ;
  assign n6183 = n6171 ^ n6134 ^ n2690 ;
  assign n6184 = n6171 & n6183 ;
  assign n6185 = n6184 ^ n6071 ^ n5758 ;
  assign n6186 = n6171 ^ n6137 ^ n2269 ;
  assign n6187 = n6171 & n6186 ;
  assign n6188 = n6187 ^ n6003 ^ n5845 ;
  assign n6189 = n6171 ^ n6138 ^ n2139 ;
  assign n6190 = n6171 & n6189 ;
  assign n6191 = n6190 ^ n6077 ^ n5789 ;
  assign n6192 = n6171 ^ n6140 ^ n1885 ;
  assign n6193 = n6171 & n6192 ;
  assign n6194 = n6193 ^ n6026 ^ n5763 ;
  assign n6195 = n6171 ^ n6142 ^ n1652 ;
  assign n6196 = n6171 & n6195 ;
  assign n6197 = n6196 ^ n6006 ^ n5812 ;
  assign n6198 = n6171 ^ n6144 ^ n1416 ;
  assign n6199 = n6171 & n6198 ;
  assign n6200 = n6199 ^ n5981 ^ n5768 ;
  assign n6201 = n6171 ^ n6146 ^ n1220 ;
  assign n6202 = n6171 & n6201 ;
  assign n6203 = n6202 ^ n6104 ^ n5855 ;
  assign n6204 = n6171 ^ n6154 ^ n572 ;
  assign n6205 = n6171 & n6204 ;
  assign n6206 = n6205 ^ n6017 ^ n5806 ;
  assign n6207 = n6171 ^ n6155 ^ n514 ;
  assign n6208 = n6171 & n6207 ;
  assign n6209 = n6208 ^ n5975 ^ n5861 ;
  assign n6210 = n6171 ^ n6156 ^ n458 ;
  assign n6211 = n6171 & n6210 ;
  assign n6212 = n6211 ^ n6089 ^ n5776 ;
  assign n6213 = n6171 ^ n6164 ^ n134 ;
  assign n6214 = n6171 & n6213 ;
  assign n6215 = n6214 ^ n6097 ^ n5779 ;
  assign n6216 = n6171 ^ n6152 ^ n716 ;
  assign n6217 = n6171 ^ n6145 ^ n1318 ;
  assign n6218 = n6171 & n6217 ;
  assign n6219 = n6171 & n6216 ;
  assign n6220 = n6171 ^ n6158 ^ n345 ;
  assign n6221 = n6171 ^ n6123 ^ n4346 ;
  assign n6222 = n6171 ^ n6161 ^ n217 ;
  assign n6223 = n6171 ^ n6131 ^ n2995 ;
  assign n6224 = n6171 ^ n6136 ^ n2404 ;
  assign n6225 = n6171 ^ n6121 ^ n4728 ;
  assign n6226 = n6171 ^ n6148 ^ n1034 ;
  assign n6227 = n6171 ^ n6147 ^ n1118 ;
  assign n6228 = n6171 ^ n6130 ^ n3141 ;
  assign n6229 = n6171 ^ n6139 ^ n2009 ;
  assign n6230 = n6218 ^ n6009 ^ n5852 ;
  assign n6231 = ( x46 & n5959 ) | ( x46 & n6171 ) | ( n5959 & n6171 ) ;
  assign n6232 = ( ~n5959 & n5962 ) | ( ~n5959 & n6231 ) | ( n5962 & n6231 ) ;
  assign n6233 = n6171 & n6224 ;
  assign n6234 = n6171 & n6225 ;
  assign n6235 = n6171 ^ n6160 ^ n261 ;
  assign n6236 = n6171 & n6223 ;
  assign n6237 = n6171 & n6220 ;
  assign n6238 = n6171 & n6228 ;
  assign n6239 = n6238 ^ n6073 ^ n5840 ;
  assign n6240 = n6237 ^ n6020 ^ n5809 ;
  assign n6241 = n6219 ^ n6042 ^ n5800 ;
  assign n6242 = n6236 ^ n6056 ^ n5846 ;
  assign n6243 = n6234 ^ n6083 ^ n5825 ;
  assign n6244 = n6233 ^ n6048 ^ n5799 ;
  assign n6245 = n6171 & n6229 ;
  assign n6246 = n6171 ^ n6129 ^ n3302 ;
  assign n6247 = n6171 ^ n6122 ^ n4534 ;
  assign n6248 = n6171 & n6247 ;
  assign n6249 = n6171 & n6235 ;
  assign n6250 = n6249 ^ n6023 ^ n5815 ;
  assign n6251 = n6171 & n6246 ;
  assign n6252 = n6171 ^ n6153 ^ n640 ;
  assign n6253 = n6171 & n6252 ;
  assign n6254 = n6248 ^ n5996 ^ n5751 ;
  assign n6255 = n6171 & n6221 ;
  assign n6256 = n6251 ^ n6050 ^ n5837 ;
  assign n6257 = n6255 ^ n5999 ^ n5782 ;
  assign n6258 = n6253 ^ n6081 ^ n5803 ;
  assign n6259 = n6171 & n6222 ;
  assign n6260 = n6171 & n6227 ;
  assign n6261 = n6259 ^ n6099 ^ n5873 ;
  assign n6262 = n6171 & n6226 ;
  assign n6263 = n6260 ^ n6012 ^ n5771 ;
  assign n6264 = n6262 ^ n6103 ^ n5792 ;
  assign n6265 = ~n6231 & n6232 ;
  assign n6266 = n6245 ^ n6069 ^ n5870 ;
  assign n6267 = n6143 ^ n1534 ^ 1'b0 ;
  assign n6268 = n6149 ^ n941 ^ 1'b0 ;
  assign n6269 = n6141 ^ n1766 ^ 1'b0 ;
  assign n6270 = n6118 ^ n5319 ^ 1'b0 ;
  assign n6271 = n6135 ^ n2544 ^ 1'b0 ;
  assign n6272 = n6171 & n6270 ;
  assign n6273 = n6272 ^ n6171 ^ n5993 ;
  assign n6274 = n6171 & n6267 ;
  assign n6275 = n6274 ^ n6171 ^ n5985 ;
  assign n6276 = n6171 & n6271 ;
  assign n6277 = n6171 & n6268 ;
  assign n6278 = n6276 ^ n6171 ^ n5989 ;
  assign n6279 = n6171 & n6269 ;
  assign n6280 = n6171 ^ n6162 ^ n179 ;
  assign n6281 = n6171 ^ n6125 ^ n3986 ;
  assign n6282 = n6277 ^ n6171 ^ n5967 ;
  assign n6283 = n6279 ^ n6171 ^ n5991 ;
  assign n6284 = n6171 ^ n6163 ^ n144 ;
  assign n6285 = n6124 ^ n4167 ^ 1'b0 ;
  assign n6286 = n6171 & n6285 ;
  assign n6287 = n6286 ^ n6171 ^ n5988 ;
  assign n6288 = n6171 ^ n6120 ^ n4915 ;
  assign n6289 = n6151 ^ n785 ^ 1'b0 ;
  assign n6290 = n6132 ^ n2839 ^ 1'b0 ;
  assign n6291 = n6171 & n6289 ;
  assign n6292 = n6291 ^ n6171 ^ n5992 ;
  assign n6293 = n6157 ^ n399 ^ 1'b0 ;
  assign n6294 = n6171 & n6293 ;
  assign n6295 = n6294 ^ n6171 ^ n5987 ;
  assign n6296 = n6171 & n6290 ;
  assign n6297 = n6296 ^ n6171 ^ n5990 ;
  assign n6298 = n6126 ^ n3804 ^ 1'b0 ;
  assign n6299 = n6171 & n6298 ;
  assign n6300 = n6171 & n6281 ;
  assign n6301 = n6299 ^ n6171 ^ n6095 ;
  assign n6302 = n6300 ^ n6013 ^ n5828 ;
  assign n6303 = n6171 & n6280 ;
  assign n6304 = n6171 & n6284 ;
  assign n6305 = n6304 ^ n6032 ^ n5818 ;
  assign n6306 = n6171 & n6288 ;
  assign n6307 = n6306 ^ n6079 ^ n5822 ;
  assign n6308 = n6109 & n6171 ;
  assign n6309 = ( ~x46 & n5964 ) | ( ~x46 & n6171 ) | ( n5964 & n6171 ) ;
  assign n6310 = x44 | x45 ;
  assign n6311 = ( n5964 & n6057 ) | ( n5964 & ~n6171 ) | ( n6057 & ~n6171 ) ;
  assign n6312 = ~x46 & n6171 ;
  assign n6313 = ( x46 & n5964 ) | ( x46 & ~n6310 ) | ( n5964 & ~n6310 ) ;
  assign n6314 = n6312 ^ x47 ^ 1'b0 ;
  assign n6315 = n6309 & n6313 ;
  assign n6316 = n6171 ^ n6117 ^ n5527 ;
  assign n6317 = ( n6171 & ~n6308 ) | ( n6171 & n6311 ) | ( ~n6308 & n6311 ) ;
  assign n6318 = n6265 | n6314 ;
  assign n6319 = ~n6315 & n6318 ;
  assign n6320 = n6171 & n6316 ;
  assign n6321 = ( n6165 & n6166 ) | ( n6165 & ~n6171 ) | ( n6166 & ~n6171 ) ;
  assign n6322 = ( n6057 & n6091 ) | ( n6057 & ~n6094 ) | ( n6091 & ~n6094 ) ;
  assign n6323 = n6317 ^ x48 ^ 1'b0 ;
  assign n6324 = ~n6170 & n6322 ;
  assign n6325 = ( ~n6091 & n6165 ) | ( ~n6091 & n6171 ) | ( n6165 & n6171 ) ;
  assign n6326 = ( ~n5743 & n6319 ) | ( ~n5743 & n6323 ) | ( n6319 & n6323 ) ;
  assign n6327 = ( n136 & n6091 ) | ( n136 & n6165 ) | ( n6091 & n6165 ) ;
  assign n6328 = n6320 ^ n5994 ^ x51 ;
  assign n6329 = n6303 ^ n6029 ^ n5876 ;
  assign n6330 = n6171 & ~n6324 ;
  assign n6331 = ( ~n5527 & n6176 ) | ( ~n5527 & n6326 ) | ( n6176 & n6326 ) ;
  assign n6332 = ( ~n5319 & n6328 ) | ( ~n5319 & n6331 ) | ( n6328 & n6331 ) ;
  assign n6333 = n6332 ^ n5124 ^ 1'b0 ;
  assign n6334 = n6159 ^ n302 ^ 1'b0 ;
  assign n6335 = ( ~n5124 & n6273 ) | ( ~n5124 & n6332 ) | ( n6273 & n6332 ) ;
  assign n6336 = ( ~n4915 & n6174 ) | ( ~n4915 & n6335 ) | ( n6174 & n6335 ) ;
  assign n6337 = ( ~n4728 & n6307 ) | ( ~n4728 & n6336 ) | ( n6307 & n6336 ) ;
  assign n6338 = ( ~n4534 & n6243 ) | ( ~n4534 & n6337 ) | ( n6243 & n6337 ) ;
  assign n6339 = ( ~n4346 & n6254 ) | ( ~n4346 & n6338 ) | ( n6254 & n6338 ) ;
  assign n6340 = ( ~n4167 & n6257 ) | ( ~n4167 & n6339 ) | ( n6257 & n6339 ) ;
  assign n6341 = ( ~n3986 & n6287 ) | ( ~n3986 & n6340 ) | ( n6287 & n6340 ) ;
  assign n6342 = ( ~n3804 & n6302 ) | ( ~n3804 & n6341 ) | ( n6302 & n6341 ) ;
  assign n6343 = ( ~n3631 & n6301 ) | ( ~n3631 & n6342 ) | ( n6301 & n6342 ) ;
  assign n6344 = ( ~n3464 & n6179 ) | ( ~n3464 & n6343 ) | ( n6179 & n6343 ) ;
  assign n6345 = ( ~n3302 & n6182 ) | ( ~n3302 & n6344 ) | ( n6182 & n6344 ) ;
  assign n6346 = n6342 ^ n3631 ^ 1'b0 ;
  assign n6347 = ( ~n3141 & n6256 ) | ( ~n3141 & n6345 ) | ( n6256 & n6345 ) ;
  assign n6348 = ~n6321 & n6327 ;
  assign n6349 = n6324 | n6348 ;
  assign n6350 = ( ~n2995 & n6239 ) | ( ~n2995 & n6347 ) | ( n6239 & n6347 ) ;
  assign n6351 = ( ~n2839 & n6242 ) | ( ~n2839 & n6350 ) | ( n6242 & n6350 ) ;
  assign n6352 = n6326 ^ n5527 ^ 1'b0 ;
  assign n6353 = n6171 & n6334 ;
  assign n6354 = n6057 | n6094 ;
  assign n6355 = ( x42 & x43 ) | ( x42 & ~n6094 ) | ( x43 & ~n6094 ) ;
  assign n6356 = n6171 ^ n6150 ^ n859 ;
  assign n6357 = n6171 & n6356 ;
  assign n6358 = n6357 ^ n5973 ^ n5795 ;
  assign n6359 = n6340 ^ n3986 ^ 1'b0 ;
  assign n6360 = ( x44 & ~n6094 ) | ( x44 & n6355 ) | ( ~n6094 & n6355 ) ;
  assign n6361 = n6351 ^ n2690 ^ 1'b0 ;
  assign n6362 = ( ~n2690 & n6297 ) | ( ~n2690 & n6351 ) | ( n6297 & n6351 ) ;
  assign n6363 = ( ~n2544 & n6185 ) | ( ~n2544 & n6362 ) | ( n6185 & n6362 ) ;
  assign n6364 = ( ~n2404 & n6278 ) | ( ~n2404 & n6363 ) | ( n6278 & n6363 ) ;
  assign n6365 = ( ~n2269 & n6244 ) | ( ~n2269 & n6364 ) | ( n6244 & n6364 ) ;
  assign n6366 = ( ~n6166 & n6354 ) | ( ~n6166 & n6360 ) | ( n6354 & n6360 ) ;
  assign n6367 = ~n6354 & n6366 ;
  assign n6368 = ( ~n2139 & n6188 ) | ( ~n2139 & n6365 ) | ( n6188 & n6365 ) ;
  assign n6369 = ( ~n2009 & n6191 ) | ( ~n2009 & n6368 ) | ( n6191 & n6368 ) ;
  assign n6370 = ( ~n1885 & n6266 ) | ( ~n1885 & n6369 ) | ( n6266 & n6369 ) ;
  assign n6371 = ( ~n1766 & n6194 ) | ( ~n1766 & n6370 ) | ( n6194 & n6370 ) ;
  assign n6372 = ( ~n1652 & n6283 ) | ( ~n1652 & n6371 ) | ( n6283 & n6371 ) ;
  assign n6373 = ( ~n1534 & n6197 ) | ( ~n1534 & n6372 ) | ( n6197 & n6372 ) ;
  assign n6374 = n6353 ^ n6171 ^ n6040 ;
  assign n6375 = ( ~n1416 & n6275 ) | ( ~n1416 & n6373 ) | ( n6275 & n6373 ) ;
  assign n6376 = ( ~n1318 & n6200 ) | ( ~n1318 & n6375 ) | ( n6200 & n6375 ) ;
  assign n6377 = ( ~n1220 & n6230 ) | ( ~n1220 & n6376 ) | ( n6230 & n6376 ) ;
  assign n6378 = ( ~n1118 & n6203 ) | ( ~n1118 & n6377 ) | ( n6203 & n6377 ) ;
  assign n6379 = ~n6091 & n6165 ;
  assign n6380 = ( ~n1034 & n6263 ) | ( ~n1034 & n6378 ) | ( n6263 & n6378 ) ;
  assign n6381 = ( ~n941 & n6264 ) | ( ~n941 & n6380 ) | ( n6264 & n6380 ) ;
  assign n6382 = n6373 ^ n1416 ^ 1'b0 ;
  assign n6383 = ( ~n859 & n6282 ) | ( ~n859 & n6381 ) | ( n6282 & n6381 ) ;
  assign n6384 = ( ~n785 & n6358 ) | ( ~n785 & n6383 ) | ( n6358 & n6383 ) ;
  assign n6385 = ( ~n716 & n6292 ) | ( ~n716 & n6384 ) | ( n6292 & n6384 ) ;
  assign n6386 = ( ~n640 & n6241 ) | ( ~n640 & n6385 ) | ( n6241 & n6385 ) ;
  assign n6387 = ( ~n572 & n6258 ) | ( ~n572 & n6386 ) | ( n6258 & n6386 ) ;
  assign n6388 = ( ~n514 & n6206 ) | ( ~n514 & n6387 ) | ( n6206 & n6387 ) ;
  assign n6389 = ( ~n458 & n6209 ) | ( ~n458 & n6388 ) | ( n6209 & n6388 ) ;
  assign n6390 = ( ~n399 & n6212 ) | ( ~n399 & n6389 ) | ( n6212 & n6389 ) ;
  assign n6391 = ( ~n345 & n6295 ) | ( ~n345 & n6390 ) | ( n6295 & n6390 ) ;
  assign n6392 = ( ~n302 & n6240 ) | ( ~n302 & n6391 ) | ( n6240 & n6391 ) ;
  assign n6393 = ( ~n261 & n6374 ) | ( ~n261 & n6392 ) | ( n6374 & n6392 ) ;
  assign n6394 = ( ~n217 & n6250 ) | ( ~n217 & n6393 ) | ( n6250 & n6393 ) ;
  assign n6395 = ( ~n179 & n6261 ) | ( ~n179 & n6394 ) | ( n6261 & n6394 ) ;
  assign n6396 = ( ~n144 & n6329 ) | ( ~n144 & n6395 ) | ( n6329 & n6395 ) ;
  assign n6397 = ( ~n134 & n6305 ) | ( ~n134 & n6396 ) | ( n6305 & n6396 ) ;
  assign n6398 = ( ~n136 & n6215 ) | ( ~n136 & n6397 ) | ( n6215 & n6397 ) ;
  assign n6399 = ( ~n136 & n6325 ) | ( ~n136 & n6398 ) | ( n6325 & n6398 ) ;
  assign n6400 = ( ~n6379 & n6398 ) | ( ~n6379 & n6399 ) | ( n6398 & n6399 ) ;
  assign n6401 = n6349 | n6400 ;
  assign n6402 = n6401 ^ n6385 ^ n640 ;
  assign n6403 = n6401 & n6402 ;
  assign n6404 = n6403 ^ n6219 ^ n6043 ;
  assign n6405 = n6352 & n6401 ;
  assign n6406 = n6392 ^ n261 ^ 1'b0 ;
  assign n6407 = n6401 & n6406 ;
  assign n6408 = n6407 ^ n6401 ^ n6374 ;
  assign n6409 = n6361 & n6401 ;
  assign n6410 = ~n6310 & n6401 ;
  assign n6411 = n6330 | n6410 ;
  assign n6412 = ( n6348 & n6400 ) | ( n6348 & ~n6410 ) | ( n6400 & ~n6410 ) ;
  assign n6413 = n6409 ^ n6401 ^ n6297 ;
  assign n6414 = ( n6410 & n6411 ) | ( n6410 & ~n6412 ) | ( n6411 & ~n6412 ) ;
  assign n6415 = n6405 ^ n6401 ^ n6176 ;
  assign n6416 = n6382 & n6401 ;
  assign n6417 = n6401 ^ n6344 ^ n3302 ;
  assign n6418 = n6346 & n6401 ;
  assign n6419 = n6416 ^ n6401 ^ n6275 ;
  assign n6420 = ( n6265 & ~n6315 ) | ( n6265 & n6401 ) | ( ~n6315 & n6401 ) ;
  assign n6421 = n6359 & n6401 ;
  assign n6422 = n6333 & n6401 ;
  assign n6423 = ~n6265 & n6420 ;
  assign n6424 = n6422 ^ n6401 ^ n6273 ;
  assign n6425 = n6421 ^ n6401 ^ n6287 ;
  assign n6426 = n6418 ^ n6401 ^ n6301 ;
  assign n6427 = n6401 & n6417 ;
  assign n6428 = n6427 ^ n6181 ^ n6068 ;
  assign n6429 = n6401 ^ n6396 ^ n134 ;
  assign n6430 = n6401 & n6429 ;
  assign n6431 = n6430 ^ n6304 ^ n6033 ;
  assign n6432 = n6401 ^ n6345 ^ n3141 ;
  assign n6433 = n6401 & n6432 ;
  assign n6434 = n6433 ^ n6251 ^ n6058 ;
  assign n6435 = n6401 ^ n6347 ^ n2995 ;
  assign n6436 = n6401 & n6435 ;
  assign n6437 = n6436 ^ n6238 ^ n6074 ;
  assign n6438 = n6401 ^ n6350 ^ n2839 ;
  assign n6439 = n6401 & n6438 ;
  assign n6440 = n6439 ^ n6236 ^ n6062 ;
  assign n6441 = n6401 ^ n6362 ^ n2544 ;
  assign n6442 = n6401 & n6441 ;
  assign n6443 = n6442 ^ n6184 ^ n6072 ;
  assign n6444 = n6401 ^ n6364 ^ n2269 ;
  assign n6445 = n6401 & n6444 ;
  assign n6446 = n6445 ^ n6233 ^ n6060 ;
  assign n6447 = n6401 ^ n6370 ^ n1766 ;
  assign n6448 = n6401 & n6447 ;
  assign n6449 = n6448 ^ n6193 ^ n6027 ;
  assign n6450 = n6401 ^ n6372 ^ n1534 ;
  assign n6451 = n6401 & n6450 ;
  assign n6452 = n6451 ^ n6196 ^ n6007 ;
  assign n6453 = n6401 ^ n6378 ^ n1034 ;
  assign n6454 = n6401 & n6453 ;
  assign n6455 = n6454 ^ n6260 ^ n6015 ;
  assign n6456 = n6401 ^ n6383 ^ n785 ;
  assign n6457 = n6401 & n6456 ;
  assign n6458 = n6457 ^ n6357 ^ n5974 ;
  assign n6459 = n6384 ^ n716 ^ 1'b0 ;
  assign n6460 = n6401 & n6459 ;
  assign n6461 = n6460 ^ n6401 ^ n6292 ;
  assign n6462 = n6401 ^ n6389 ^ n399 ;
  assign n6463 = n6401 & n6462 ;
  assign n6464 = n6463 ^ n6211 ^ n6090 ;
  assign n6465 = n6390 ^ n345 ^ 1'b0 ;
  assign n6466 = n6401 & n6465 ;
  assign n6467 = n6466 ^ n6401 ^ n6295 ;
  assign n6468 = n6401 ^ n6393 ^ n217 ;
  assign n6469 = n6401 & n6468 ;
  assign n6470 = n6469 ^ n6249 ^ n6024 ;
  assign n6471 = n6401 ^ n6394 ^ n179 ;
  assign n6472 = n6401 & n6471 ;
  assign n6473 = n6472 ^ n6259 ^ n6102 ;
  assign n6474 = n6401 ^ n6337 ^ n4534 ;
  assign n6475 = n6401 & n6474 ;
  assign n6476 = n6475 ^ n6234 ^ n6092 ;
  assign n6477 = ( x44 & n6168 ) | ( x44 & n6401 ) | ( n6168 & n6401 ) ;
  assign n6478 = ( ~n6168 & n6367 ) | ( ~n6168 & n6477 ) | ( n6367 & n6477 ) ;
  assign n6479 = ~n6477 & n6478 ;
  assign n6480 = n6401 ^ n6319 ^ n5743 ;
  assign n6481 = n6401 & n6480 ;
  assign n6482 = n6481 ^ n6317 ^ x48 ;
  assign n6483 = n6401 ^ n6331 ^ n5319 ;
  assign n6484 = n6401 & n6483 ;
  assign n6485 = n6484 ^ n6320 ^ n6107 ;
  assign n6486 = n6401 ^ n6335 ^ n4915 ;
  assign n6487 = n6401 & n6486 ;
  assign n6488 = n6487 ^ n6173 ^ n6065 ;
  assign n6489 = n6401 ^ n6336 ^ n4728 ;
  assign n6490 = n6401 & n6489 ;
  assign n6491 = n6490 ^ n6306 ^ n6080 ;
  assign n6492 = n6401 ^ n6339 ^ n4167 ;
  assign n6493 = n6401 & n6492 ;
  assign n6494 = n6493 ^ n6255 ^ n6000 ;
  assign n6495 = n6401 ^ n6341 ^ n3804 ;
  assign n6496 = n6401 & n6495 ;
  assign n6497 = n6496 ^ n6300 ^ n6014 ;
  assign n6498 = n6401 ^ n6343 ^ n3464 ;
  assign n6499 = n6401 & n6498 ;
  assign n6500 = n6499 ^ n6178 ^ n6076 ;
  assign n6501 = n6363 ^ n2404 ^ 1'b0 ;
  assign n6502 = n6401 & n6501 ;
  assign n6503 = n6502 ^ n6401 ^ n6278 ;
  assign n6504 = n6401 ^ n6365 ^ n2139 ;
  assign n6505 = n6401 & n6504 ;
  assign n6506 = n6505 ^ n6187 ^ n6004 ;
  assign n6507 = n6401 ^ n6368 ^ n2009 ;
  assign n6508 = n6401 & n6507 ;
  assign n6509 = n6508 ^ n6190 ^ n6078 ;
  assign n6510 = n6401 ^ n6369 ^ n1885 ;
  assign n6511 = n6401 & n6510 ;
  assign n6512 = n6511 ^ n6245 ^ n6070 ;
  assign n6513 = n6371 ^ n1652 ^ 1'b0 ;
  assign n6514 = n6401 & n6513 ;
  assign n6515 = n6514 ^ n6401 ^ n6283 ;
  assign n6516 = n6401 ^ n6338 ^ n4346 ;
  assign n6517 = n6401 & n6516 ;
  assign n6518 = n6517 ^ n6248 ^ n5997 ;
  assign n6519 = n6401 ^ n6375 ^ n1318 ;
  assign n6520 = n6401 & n6519 ;
  assign n6521 = n6520 ^ n6199 ^ n5983 ;
  assign n6522 = n6401 ^ n6376 ^ n1220 ;
  assign n6523 = n6401 & n6522 ;
  assign n6524 = n6523 ^ n6218 ^ n6010 ;
  assign n6525 = n6401 ^ n6377 ^ n1118 ;
  assign n6526 = n6401 & n6525 ;
  assign n6527 = n6526 ^ n6202 ^ n6106 ;
  assign n6528 = n6401 ^ n6380 ^ n941 ;
  assign n6529 = n6401 & n6528 ;
  assign n6530 = n6529 ^ n6262 ^ n6105 ;
  assign n6531 = n6381 ^ n859 ^ 1'b0 ;
  assign n6532 = n6401 & n6531 ;
  assign n6533 = n6532 ^ n6401 ^ n6282 ;
  assign n6534 = n6401 ^ n6386 ^ n572 ;
  assign n6535 = n6401 & n6534 ;
  assign n6536 = n6535 ^ n6253 ^ n6082 ;
  assign n6537 = n6401 ^ n6387 ^ n514 ;
  assign n6538 = n6401 & n6537 ;
  assign n6539 = n6538 ^ n6205 ^ n6018 ;
  assign n6540 = n6401 ^ n6388 ^ n458 ;
  assign n6541 = n6401 & n6540 ;
  assign n6542 = n6541 ^ n6208 ^ n5976 ;
  assign n6543 = n6401 ^ n6391 ^ n302 ;
  assign n6544 = n6401 & n6543 ;
  assign n6545 = n6544 ^ n6237 ^ n6021 ;
  assign n6546 = n6401 ^ n6395 ^ n144 ;
  assign n6547 = n6401 & n6546 ;
  assign n6548 = n6547 ^ n6303 ^ n6030 ;
  assign n6549 = x42 | x43 ;
  assign n6550 = ~x44 & n6401 ;
  assign n6551 = n6550 ^ x45 ^ 1'b0 ;
  assign n6552 = n6479 | n6551 ;
  assign n6553 = ( ~x44 & n6171 ) | ( ~x44 & n6401 ) | ( n6171 & n6401 ) ;
  assign n6554 = ( x44 & n6171 ) | ( x44 & ~n6549 ) | ( n6171 & ~n6549 ) ;
  assign n6555 = n6553 & n6554 ;
  assign n6556 = n6414 ^ x46 ^ 1'b0 ;
  assign n6557 = n6423 ^ n6312 ^ x47 ;
  assign n6558 = n6552 & ~n6555 ;
  assign n6559 = ( ~n5964 & n6556 ) | ( ~n5964 & n6558 ) | ( n6556 & n6558 ) ;
  assign n6560 = ~n6215 & n6397 ;
  assign n6561 = ( ~n5743 & n6557 ) | ( ~n5743 & n6559 ) | ( n6557 & n6559 ) ;
  assign n6562 = ( ~n5527 & n6482 ) | ( ~n5527 & n6561 ) | ( n6482 & n6561 ) ;
  assign n6563 = ( ~n5319 & n6415 ) | ( ~n5319 & n6562 ) | ( n6415 & n6562 ) ;
  assign n6564 = ( ~n5124 & n6485 ) | ( ~n5124 & n6563 ) | ( n6485 & n6563 ) ;
  assign n6565 = ( n6215 & n6397 ) | ( n6215 & ~n6401 ) | ( n6397 & ~n6401 ) ;
  assign n6566 = ( n136 & n6215 ) | ( n136 & n6397 ) | ( n6215 & n6397 ) ;
  assign n6567 = ( ~n4915 & n6424 ) | ( ~n4915 & n6564 ) | ( n6424 & n6564 ) ;
  assign n6568 = ( ~n4728 & n6488 ) | ( ~n4728 & n6567 ) | ( n6488 & n6567 ) ;
  assign n6569 = ( ~n6215 & n6397 ) | ( ~n6215 & n6401 ) | ( n6397 & n6401 ) ;
  assign n6570 = ( ~n4534 & n6491 ) | ( ~n4534 & n6568 ) | ( n6491 & n6568 ) ;
  assign n6571 = ( ~n4346 & n6476 ) | ( ~n4346 & n6570 ) | ( n6476 & n6570 ) ;
  assign n6572 = ( ~n4167 & n6518 ) | ( ~n4167 & n6571 ) | ( n6518 & n6571 ) ;
  assign n6573 = ( ~n3986 & n6494 ) | ( ~n3986 & n6572 ) | ( n6494 & n6572 ) ;
  assign n6574 = ( ~n3804 & n6425 ) | ( ~n3804 & n6573 ) | ( n6425 & n6573 ) ;
  assign n6575 = ( ~n3631 & n6497 ) | ( ~n3631 & n6574 ) | ( n6497 & n6574 ) ;
  assign n6576 = ( ~n3464 & n6426 ) | ( ~n3464 & n6575 ) | ( n6426 & n6575 ) ;
  assign n6577 = ( ~n3302 & n6500 ) | ( ~n3302 & n6576 ) | ( n6500 & n6576 ) ;
  assign n6578 = ( ~n3141 & n6428 ) | ( ~n3141 & n6577 ) | ( n6428 & n6577 ) ;
  assign n6579 = ( ~n2995 & n6434 ) | ( ~n2995 & n6578 ) | ( n6434 & n6578 ) ;
  assign n6580 = ( ~n2839 & n6437 ) | ( ~n2839 & n6579 ) | ( n6437 & n6579 ) ;
  assign n6581 = ( ~n2690 & n6440 ) | ( ~n2690 & n6580 ) | ( n6440 & n6580 ) ;
  assign n6582 = ( ~n2544 & n6413 ) | ( ~n2544 & n6581 ) | ( n6413 & n6581 ) ;
  assign n6583 = ( ~n2404 & n6443 ) | ( ~n2404 & n6582 ) | ( n6443 & n6582 ) ;
  assign n6584 = ( ~n2269 & n6503 ) | ( ~n2269 & n6583 ) | ( n6503 & n6583 ) ;
  assign n6585 = ( ~n2139 & n6446 ) | ( ~n2139 & n6584 ) | ( n6446 & n6584 ) ;
  assign n6586 = ( ~n2009 & n6506 ) | ( ~n2009 & n6585 ) | ( n6506 & n6585 ) ;
  assign n6587 = ( ~n1885 & n6509 ) | ( ~n1885 & n6586 ) | ( n6509 & n6586 ) ;
  assign n6588 = ( ~n1766 & n6512 ) | ( ~n1766 & n6587 ) | ( n6512 & n6587 ) ;
  assign n6589 = ( ~n1652 & n6449 ) | ( ~n1652 & n6588 ) | ( n6449 & n6588 ) ;
  assign n6590 = ( ~n1534 & n6515 ) | ( ~n1534 & n6589 ) | ( n6515 & n6589 ) ;
  assign n6591 = ( ~n1416 & n6452 ) | ( ~n1416 & n6590 ) | ( n6452 & n6590 ) ;
  assign n6592 = n6575 ^ n3464 ^ 1'b0 ;
  assign n6593 = n6581 ^ n2544 ^ 1'b0 ;
  assign n6594 = ( ~n1318 & n6419 ) | ( ~n1318 & n6591 ) | ( n6419 & n6591 ) ;
  assign n6595 = n6583 ^ n2269 ^ 1'b0 ;
  assign n6596 = ( ~n1220 & n6521 ) | ( ~n1220 & n6594 ) | ( n6521 & n6594 ) ;
  assign n6597 = ( ~n1118 & n6524 ) | ( ~n1118 & n6596 ) | ( n6524 & n6596 ) ;
  assign n6598 = ( ~n1034 & n6527 ) | ( ~n1034 & n6597 ) | ( n6527 & n6597 ) ;
  assign n6599 = n6562 ^ n5319 ^ 1'b0 ;
  assign n6600 = n6573 ^ n3804 ^ 1'b0 ;
  assign n6601 = n6589 ^ n1534 ^ 1'b0 ;
  assign n6602 = n6564 ^ n4915 ^ 1'b0 ;
  assign n6603 = ( n6431 & ~n6560 ) | ( n6431 & n6569 ) | ( ~n6560 & n6569 ) ;
  assign n6604 = ( ~n941 & n6455 ) | ( ~n941 & n6598 ) | ( n6455 & n6598 ) ;
  assign n6605 = ~n6397 & n6566 ;
  assign n6606 = ( ~n6565 & n6566 ) | ( ~n6565 & n6605 ) | ( n6566 & n6605 ) ;
  assign n6607 = ( ~n859 & n6530 ) | ( ~n859 & n6604 ) | ( n6530 & n6604 ) ;
  assign n6608 = n6607 ^ n785 ^ 1'b0 ;
  assign n6609 = ( ~n785 & n6533 ) | ( ~n785 & n6607 ) | ( n6533 & n6607 ) ;
  assign n6610 = n6591 ^ n1318 ^ 1'b0 ;
  assign n6611 = ( ~n716 & n6458 ) | ( ~n716 & n6609 ) | ( n6458 & n6609 ) ;
  assign n6612 = ( ~n640 & n6461 ) | ( ~n640 & n6611 ) | ( n6461 & n6611 ) ;
  assign n6613 = ( ~n572 & n6404 ) | ( ~n572 & n6612 ) | ( n6404 & n6612 ) ;
  assign n6614 = ( ~n514 & n6536 ) | ( ~n514 & n6613 ) | ( n6536 & n6613 ) ;
  assign n6615 = ( ~n458 & n6539 ) | ( ~n458 & n6614 ) | ( n6539 & n6614 ) ;
  assign n6616 = ( ~n399 & n6542 ) | ( ~n399 & n6615 ) | ( n6542 & n6615 ) ;
  assign n6617 = ( ~n345 & n6464 ) | ( ~n345 & n6616 ) | ( n6464 & n6616 ) ;
  assign n6618 = ( ~n302 & n6467 ) | ( ~n302 & n6617 ) | ( n6467 & n6617 ) ;
  assign n6619 = ( ~n261 & n6545 ) | ( ~n261 & n6618 ) | ( n6545 & n6618 ) ;
  assign n6620 = ( ~n217 & n6408 ) | ( ~n217 & n6619 ) | ( n6408 & n6619 ) ;
  assign n6621 = ( ~n179 & n6470 ) | ( ~n179 & n6620 ) | ( n6470 & n6620 ) ;
  assign n6622 = ( ~n144 & n6473 ) | ( ~n144 & n6621 ) | ( n6473 & n6621 ) ;
  assign n6623 = ( ~n134 & n6548 ) | ( ~n134 & n6622 ) | ( n6548 & n6622 ) ;
  assign n6624 = n6431 & n6623 ;
  assign n6625 = ( n6215 & ~n6401 ) | ( n6215 & n6624 ) | ( ~n6401 & n6624 ) ;
  assign n6626 = ( ~x30 & n6603 ) | ( ~x30 & n6623 ) | ( n6603 & n6623 ) ;
  assign n6627 = ~n136 & n6626 ;
  assign n6628 = n6624 | n6627 ;
  assign n6629 = ( n6606 & ~n6625 ) | ( n6606 & n6628 ) | ( ~n6625 & n6628 ) ;
  assign n6630 = n6625 | n6629 ;
  assign n6631 = n6630 ^ n6622 ^ n134 ;
  assign n6632 = n6630 & n6631 ;
  assign n6633 = ( n6479 & ~n6555 ) | ( n6479 & n6630 ) | ( ~n6555 & n6630 ) ;
  assign n6634 = ~n6479 & n6633 ;
  assign n6635 = n6632 ^ n6547 ^ n6329 ;
  assign n6636 = n6599 & n6630 ;
  assign n6637 = n6636 ^ n6630 ^ n6415 ;
  assign n6638 = n6602 & n6630 ;
  assign n6639 = n6638 ^ n6630 ^ n6424 ;
  assign n6640 = n6600 & n6630 ;
  assign n6641 = n6640 ^ n6630 ^ n6425 ;
  assign n6642 = n6592 & n6630 ;
  assign n6643 = n6642 ^ n6630 ^ n6426 ;
  assign n6644 = n6593 & n6630 ;
  assign n6645 = n6644 ^ n6630 ^ n6413 ;
  assign n6646 = n6595 & n6630 ;
  assign n6647 = n6646 ^ n6630 ^ n6503 ;
  assign n6648 = n6630 ^ n6586 ^ n1885 ;
  assign n6649 = n6630 & n6648 ;
  assign n6650 = n6649 ^ n6508 ^ n6191 ;
  assign n6651 = n6601 & n6630 ;
  assign n6652 = n6651 ^ n6630 ^ n6515 ;
  assign n6653 = n6610 & n6630 ;
  assign n6654 = n6653 ^ n6630 ^ n6419 ;
  assign n6655 = n6608 & n6630 ;
  assign n6656 = n6655 ^ n6630 ^ n6533 ;
  assign n6657 = n6630 ^ n6612 ^ n572 ;
  assign n6658 = n6630 & n6657 ;
  assign n6659 = n6658 ^ n6403 ^ n6241 ;
  assign n6660 = n6630 ^ n6563 ^ n5124 ;
  assign n6661 = n6630 & n6660 ;
  assign n6662 = n6661 ^ n6484 ^ n6328 ;
  assign n6663 = n6630 ^ n6567 ^ n4728 ;
  assign n6664 = n6630 & n6663 ;
  assign n6665 = n6664 ^ n6487 ^ n6174 ;
  assign n6666 = n6630 ^ n6576 ^ n3302 ;
  assign n6667 = n6630 & n6666 ;
  assign n6668 = n6667 ^ n6499 ^ n6179 ;
  assign n6669 = n6630 ^ n6578 ^ n2995 ;
  assign n6670 = n6630 & n6669 ;
  assign n6671 = n6670 ^ n6433 ^ n6256 ;
  assign n6672 = n6630 ^ n6582 ^ n2404 ;
  assign n6673 = n6630 & n6672 ;
  assign n6674 = n6673 ^ n6442 ^ n6185 ;
  assign n6675 = n6630 ^ n6584 ^ n2139 ;
  assign n6676 = n6630 & n6675 ;
  assign n6677 = n6676 ^ n6445 ^ n6244 ;
  assign n6678 = n6630 ^ n6585 ^ n2009 ;
  assign n6679 = n6630 & n6678 ;
  assign n6680 = n6679 ^ n6505 ^ n6188 ;
  assign n6681 = n6630 ^ n6588 ^ n1652 ;
  assign n6682 = n6630 & n6681 ;
  assign n6683 = n6682 ^ n6448 ^ n6194 ;
  assign n6684 = n6630 ^ n6590 ^ n1416 ;
  assign n6685 = n6630 & n6684 ;
  assign n6686 = n6685 ^ n6451 ^ n6197 ;
  assign n6687 = n6630 ^ n6594 ^ n1220 ;
  assign n6688 = n6630 & n6687 ;
  assign n6689 = n6688 ^ n6520 ^ n6200 ;
  assign n6690 = n6630 ^ n6598 ^ n941 ;
  assign n6691 = n6630 & n6690 ;
  assign n6692 = n6691 ^ n6454 ^ n6263 ;
  assign n6693 = n6630 ^ n6604 ^ n859 ;
  assign n6694 = n6630 & n6693 ;
  assign n6695 = n6694 ^ n6529 ^ n6264 ;
  assign n6696 = n6630 ^ n6615 ^ n399 ;
  assign n6697 = n6630 & n6696 ;
  assign n6698 = n6697 ^ n6541 ^ n6209 ;
  assign n6699 = n6630 ^ n6616 ^ n345 ;
  assign n6700 = n6630 & n6699 ;
  assign n6701 = n6700 ^ n6463 ^ n6212 ;
  assign n6702 = n6630 ^ n6614 ^ n458 ;
  assign n6703 = n6630 ^ n6609 ^ n716 ;
  assign n6704 = n6630 ^ n6577 ^ n3141 ;
  assign n6705 = n6630 ^ n6574 ^ n3631 ;
  assign n6706 = n6630 ^ n6570 ^ n4346 ;
  assign n6707 = n6630 ^ n6620 ^ n179 ;
  assign n6708 = n6630 ^ n6618 ^ n261 ;
  assign n6709 = n6630 ^ n6561 ^ n5527 ;
  assign n6710 = n6630 & n6709 ;
  assign n6711 = n6619 ^ n217 ^ 1'b0 ;
  assign n6712 = n6630 ^ n6597 ^ n1034 ;
  assign n6713 = n6630 ^ n6568 ^ n4534 ;
  assign n6714 = n6630 ^ n6596 ^ n1118 ;
  assign n6715 = n6630 ^ n6572 ^ n3986 ;
  assign n6716 = n6617 ^ n302 ^ 1'b0 ;
  assign n6717 = n6630 & n6716 ;
  assign n6718 = n6630 ^ n6579 ^ n2839 ;
  assign n6719 = n6630 ^ n6571 ^ n4167 ;
  assign n6720 = n6630 ^ n6580 ^ n2690 ;
  assign n6721 = n6630 ^ n6613 ^ n514 ;
  assign n6722 = n6630 ^ n6621 ^ n144 ;
  assign n6723 = n6630 ^ n6587 ^ n1766 ;
  assign n6724 = n6630 ^ n6559 ^ n5743 ;
  assign n6725 = n6634 ^ n6550 ^ x45 ;
  assign n6726 = n6710 ^ n6481 ^ n6323 ;
  assign n6727 = n6630 & n6721 ;
  assign n6728 = n6727 ^ n6535 ^ n6258 ;
  assign n6729 = n6630 & n6708 ;
  assign n6730 = n6729 ^ n6544 ^ n6240 ;
  assign n6731 = n6630 & n6705 ;
  assign n6732 = n6731 ^ n6496 ^ n6302 ;
  assign n6733 = n6630 & n6713 ;
  assign n6734 = n5964 & n6558 ;
  assign n6735 = n6733 ^ n6490 ^ n6307 ;
  assign n6736 = ~n6549 & n6630 ;
  assign n6737 = n6606 & ~n6736 ;
  assign n6738 = n6630 & n6714 ;
  assign n6739 = n6738 ^ n6523 ^ n6230 ;
  assign n6740 = n6630 & n6720 ;
  assign n6741 = n6740 ^ n6439 ^ n6242 ;
  assign n6742 = n6630 & n6719 ;
  assign n6743 = n6742 ^ n6517 ^ n6254 ;
  assign n6744 = n6630 & n6712 ;
  assign n6745 = n6744 ^ n6526 ^ n6203 ;
  assign n6746 = ( n6401 & ~n6628 ) | ( n6401 & n6736 ) | ( ~n6628 & n6736 ) ;
  assign n6747 = n6630 & n6718 ;
  assign n6748 = n6747 ^ n6436 ^ n6239 ;
  assign n6749 = n6630 & n6723 ;
  assign n6750 = n6749 ^ n6511 ^ n6266 ;
  assign n6751 = ( ~n5964 & n6630 ) | ( ~n5964 & n6734 ) | ( n6630 & n6734 ) ;
  assign n6752 = ( ~n6558 & n6734 ) | ( ~n6558 & n6751 ) | ( n6734 & n6751 ) ;
  assign n6753 = n6752 ^ n6414 ^ x46 ;
  assign n6754 = n6630 & n6724 ;
  assign n6755 = n6630 & n6707 ;
  assign n6756 = ( n6736 & ~n6737 ) | ( n6736 & n6746 ) | ( ~n6737 & n6746 ) ;
  assign n6757 = n6630 & n6702 ;
  assign n6758 = n6757 ^ n6538 ^ n6206 ;
  assign n6759 = n6630 & n6703 ;
  assign n6760 = n6630 & n6706 ;
  assign n6761 = n6759 ^ n6457 ^ n6358 ;
  assign n6762 = n6760 ^ n6475 ^ n6243 ;
  assign n6763 = n6755 ^ n6469 ^ n6250 ;
  assign n6764 = n6630 & n6722 ;
  assign n6765 = n6630 & n6715 ;
  assign n6766 = n6765 ^ n6493 ^ n6257 ;
  assign n6767 = n6611 ^ n640 ^ 1'b0 ;
  assign n6768 = n6630 & n6704 ;
  assign n6769 = n6768 ^ n6427 ^ n6182 ;
  assign n6770 = n6717 ^ n6630 ^ n6467 ;
  assign n6771 = n6630 & n6767 ;
  assign n6772 = n6771 ^ n6630 ^ n6461 ;
  assign n6773 = n6630 & n6711 ;
  assign n6774 = n6764 ^ n6472 ^ n6261 ;
  assign n6775 = n6754 ^ n6423 ^ n6314 ;
  assign n6776 = n6773 ^ n6630 ^ n6408 ;
  assign n6777 = n6756 ^ x44 ^ 1'b0 ;
  assign n6778 = x40 | x41 ;
  assign n6779 = ( x42 & ~n6400 ) | ( x42 & n6778 ) | ( ~n6400 & n6778 ) ;
  assign n6780 = ( x42 & n6401 ) | ( x42 & ~n6778 ) | ( n6401 & ~n6778 ) ;
  assign n6781 = ( ~x42 & n6401 ) | ( ~x42 & n6630 ) | ( n6401 & n6630 ) ;
  assign n6782 = n6780 & n6781 ;
  assign n6783 = x42 & n6630 ;
  assign n6784 = ( ~n6401 & n6779 ) | ( ~n6401 & n6783 ) | ( n6779 & n6783 ) ;
  assign n6785 = ~n6783 & n6784 ;
  assign n6786 = ( ~n6431 & n6624 ) | ( ~n6431 & n6630 ) | ( n6624 & n6630 ) ;
  assign n6787 = n6623 & ~n6624 ;
  assign n6788 = ( n136 & n6431 ) | ( n136 & n6623 ) | ( n6431 & n6623 ) ;
  assign n6789 = n6783 ^ n6630 ^ x43 ;
  assign n6790 = ( n6623 & n6624 ) | ( n6623 & ~n6630 ) | ( n6624 & ~n6630 ) ;
  assign n6791 = n6785 | n6789 ;
  assign n6792 = ~n6782 & n6791 ;
  assign n6793 = n6431 & ~n6630 ;
  assign n6794 = ( ~n6171 & n6777 ) | ( ~n6171 & n6792 ) | ( n6777 & n6792 ) ;
  assign n6795 = ( ~n5964 & n6725 ) | ( ~n5964 & n6794 ) | ( n6725 & n6794 ) ;
  assign n6796 = ( ~n5743 & n6753 ) | ( ~n5743 & n6795 ) | ( n6753 & n6795 ) ;
  assign n6797 = ( ~n5527 & n6775 ) | ( ~n5527 & n6796 ) | ( n6775 & n6796 ) ;
  assign n6798 = ( ~n5319 & n6726 ) | ( ~n5319 & n6797 ) | ( n6726 & n6797 ) ;
  assign n6799 = n6782 | n6785 ;
  assign n6800 = ( ~n5124 & n6637 ) | ( ~n5124 & n6798 ) | ( n6637 & n6798 ) ;
  assign n6801 = ( ~n4915 & n6662 ) | ( ~n4915 & n6800 ) | ( n6662 & n6800 ) ;
  assign n6802 = ( ~n4728 & n6639 ) | ( ~n4728 & n6801 ) | ( n6639 & n6801 ) ;
  assign n6803 = ( ~n4534 & n6665 ) | ( ~n4534 & n6802 ) | ( n6665 & n6802 ) ;
  assign n6804 = ( ~n4346 & n6735 ) | ( ~n4346 & n6803 ) | ( n6735 & n6803 ) ;
  assign n6805 = ( n6624 & n6786 ) | ( n6624 & ~n6787 ) | ( n6786 & ~n6787 ) ;
  assign n6806 = ( ~n4167 & n6762 ) | ( ~n4167 & n6804 ) | ( n6762 & n6804 ) ;
  assign n6807 = ( ~n3986 & n6743 ) | ( ~n3986 & n6806 ) | ( n6743 & n6806 ) ;
  assign n6808 = ( ~n3804 & n6766 ) | ( ~n3804 & n6807 ) | ( n6766 & n6807 ) ;
  assign n6809 = ( ~n3631 & n6641 ) | ( ~n3631 & n6808 ) | ( n6641 & n6808 ) ;
  assign n6810 = ( ~n3464 & n6732 ) | ( ~n3464 & n6809 ) | ( n6732 & n6809 ) ;
  assign n6811 = ( ~n3302 & n6643 ) | ( ~n3302 & n6810 ) | ( n6643 & n6810 ) ;
  assign n6812 = ( ~n3141 & n6668 ) | ( ~n3141 & n6811 ) | ( n6668 & n6811 ) ;
  assign n6813 = ( ~n2995 & n6769 ) | ( ~n2995 & n6812 ) | ( n6769 & n6812 ) ;
  assign n6814 = ( ~n2839 & n6671 ) | ( ~n2839 & n6813 ) | ( n6671 & n6813 ) ;
  assign n6815 = ( ~n2690 & n6748 ) | ( ~n2690 & n6814 ) | ( n6748 & n6814 ) ;
  assign n6816 = ( ~n2544 & n6741 ) | ( ~n2544 & n6815 ) | ( n6741 & n6815 ) ;
  assign n6817 = n6788 & ~n6790 ;
  assign n6818 = n6793 | n6817 ;
  assign n6819 = ( n6627 & n6805 ) | ( n6627 & ~n6818 ) | ( n6805 & ~n6818 ) ;
  assign n6820 = ( ~n2404 & n6645 ) | ( ~n2404 & n6816 ) | ( n6645 & n6816 ) ;
  assign n6821 = ( ~n2269 & n6674 ) | ( ~n2269 & n6820 ) | ( n6674 & n6820 ) ;
  assign n6822 = ( x35 & x36 ) | ( x35 & ~n6817 ) | ( x36 & ~n6817 ) ;
  assign n6823 = ( ~n2139 & n6647 ) | ( ~n2139 & n6821 ) | ( n6647 & n6821 ) ;
  assign n6824 = ( ~n2009 & n6677 ) | ( ~n2009 & n6823 ) | ( n6677 & n6823 ) ;
  assign n6825 = ( x37 & ~n6817 ) | ( x37 & n6822 ) | ( ~n6817 & n6822 ) ;
  assign n6826 = ( ~n1885 & n6680 ) | ( ~n1885 & n6824 ) | ( n6680 & n6824 ) ;
  assign n6827 = ( ~n1766 & n6650 ) | ( ~n1766 & n6826 ) | ( n6650 & n6826 ) ;
  assign n6828 = ( ~n1652 & n6750 ) | ( ~n1652 & n6827 ) | ( n6750 & n6827 ) ;
  assign n6829 = ( ~n1534 & n6683 ) | ( ~n1534 & n6828 ) | ( n6683 & n6828 ) ;
  assign n6830 = ( ~n1416 & n6652 ) | ( ~n1416 & n6829 ) | ( n6652 & n6829 ) ;
  assign n6831 = ( ~n1318 & n6686 ) | ( ~n1318 & n6830 ) | ( n6686 & n6830 ) ;
  assign n6832 = ( ~n1220 & n6654 ) | ( ~n1220 & n6831 ) | ( n6654 & n6831 ) ;
  assign n6833 = ( ~n1118 & n6689 ) | ( ~n1118 & n6832 ) | ( n6689 & n6832 ) ;
  assign n6834 = ( ~n1034 & n6739 ) | ( ~n1034 & n6833 ) | ( n6739 & n6833 ) ;
  assign n6835 = ( ~n941 & n6745 ) | ( ~n941 & n6834 ) | ( n6745 & n6834 ) ;
  assign n6836 = ( ~n859 & n6692 ) | ( ~n859 & n6835 ) | ( n6692 & n6835 ) ;
  assign n6837 = ( ~n785 & n6695 ) | ( ~n785 & n6836 ) | ( n6695 & n6836 ) ;
  assign n6838 = ( ~n716 & n6656 ) | ( ~n716 & n6837 ) | ( n6656 & n6837 ) ;
  assign n6839 = ( ~n640 & n6761 ) | ( ~n640 & n6838 ) | ( n6761 & n6838 ) ;
  assign n6840 = ( ~n572 & n6772 ) | ( ~n572 & n6839 ) | ( n6772 & n6839 ) ;
  assign n6841 = ( ~n514 & n6659 ) | ( ~n514 & n6840 ) | ( n6659 & n6840 ) ;
  assign n6842 = ( ~n458 & n6728 ) | ( ~n458 & n6841 ) | ( n6728 & n6841 ) ;
  assign n6843 = ( ~n399 & n6758 ) | ( ~n399 & n6842 ) | ( n6758 & n6842 ) ;
  assign n6844 = ( ~n345 & n6698 ) | ( ~n345 & n6843 ) | ( n6698 & n6843 ) ;
  assign n6845 = ( ~n302 & n6701 ) | ( ~n302 & n6844 ) | ( n6701 & n6844 ) ;
  assign n6846 = ( ~n261 & n6770 ) | ( ~n261 & n6845 ) | ( n6770 & n6845 ) ;
  assign n6847 = ( ~n217 & n6730 ) | ( ~n217 & n6846 ) | ( n6730 & n6846 ) ;
  assign n6848 = ( ~n179 & n6776 ) | ( ~n179 & n6847 ) | ( n6776 & n6847 ) ;
  assign n6849 = ( ~n144 & n6763 ) | ( ~n144 & n6848 ) | ( n6763 & n6848 ) ;
  assign n6850 = ( ~n134 & n6774 ) | ( ~n134 & n6849 ) | ( n6774 & n6849 ) ;
  assign n6851 = ( ~n136 & n6635 ) | ( ~n136 & n6850 ) | ( n6635 & n6850 ) ;
  assign n6852 = n6805 | n6851 ;
  assign n6853 = n6635 & n6850 ;
  assign n6854 = ( n6818 & n6825 ) | ( n6818 & ~n6853 ) | ( n6825 & ~n6853 ) ;
  assign n6855 = ~n6818 & n6854 ;
  assign n6856 = ~n136 & n6852 ;
  assign n6857 = n6853 | n6856 ;
  assign n6858 = n6818 | n6857 ;
  assign n6859 = n6799 & n6858 ;
  assign n6860 = n6858 ^ n6794 ^ n5964 ;
  assign n6861 = n6858 & n6860 ;
  assign n6862 = n6858 ^ n6800 ^ n4915 ;
  assign n6863 = n6859 ^ n6858 ^ n6789 ;
  assign n6864 = n6858 & n6862 ;
  assign n6865 = ~n6778 & n6858 ;
  assign n6866 = n6858 ^ n6809 ^ n3464 ;
  assign n6867 = n6858 ^ n6796 ^ n5527 ;
  assign n6868 = n6858 ^ n6827 ^ n1652 ;
  assign n6869 = n6861 ^ n6634 ^ n6551 ;
  assign n6870 = n6858 ^ n6849 ^ n134 ;
  assign n6871 = n6858 ^ n6807 ^ n3804 ;
  assign n6872 = n6858 & n6867 ;
  assign n6873 = n6858 & n6870 ;
  assign n6874 = n6858 & n6871 ;
  assign n6875 = n6873 ^ n6764 ^ n6473 ;
  assign n6876 = n6858 ^ n6797 ^ n5319 ;
  assign n6877 = n6858 & n6876 ;
  assign n6878 = n6877 ^ n6710 ^ n6482 ;
  assign n6879 = n6858 & n6866 ;
  assign n6880 = n6857 & ~n6865 ;
  assign n6881 = ( n6819 & n6865 ) | ( n6819 & ~n6880 ) | ( n6865 & ~n6880 ) ;
  assign n6882 = n6858 & n6868 ;
  assign n6883 = n6874 ^ n6765 ^ n6494 ;
  assign n6884 = n6879 ^ n6731 ^ n6497 ;
  assign n6885 = n6882 ^ n6749 ^ n6512 ;
  assign n6886 = n6864 ^ n6661 ^ n6485 ;
  assign n6887 = n6872 ^ n6754 ^ n6557 ;
  assign n6888 = n6858 ^ n6804 ^ n4167 ;
  assign n6889 = n6858 & n6888 ;
  assign n6890 = n6889 ^ n6760 ^ n6476 ;
  assign n6891 = n6858 ^ n6812 ^ n2995 ;
  assign n6892 = n6858 & n6891 ;
  assign n6893 = n6892 ^ n6768 ^ n6428 ;
  assign n6894 = n6858 ^ n6813 ^ n2839 ;
  assign n6895 = n6858 & n6894 ;
  assign n6896 = n6858 ^ n6814 ^ n2690 ;
  assign n6897 = n6858 & n6896 ;
  assign n6898 = n6897 ^ n6747 ^ n6437 ;
  assign n6899 = n6858 ^ n6815 ^ n2544 ;
  assign n6900 = n6858 & n6899 ;
  assign n6901 = n6900 ^ n6740 ^ n6440 ;
  assign n6902 = n6821 ^ n2139 ^ 1'b0 ;
  assign n6903 = n6858 & n6902 ;
  assign n6904 = n6903 ^ n6858 ^ n6647 ;
  assign n6905 = n6858 ^ n6823 ^ n2009 ;
  assign n6906 = n6895 ^ n6670 ^ n6434 ;
  assign n6907 = n6858 & n6905 ;
  assign n6908 = n6907 ^ n6676 ^ n6446 ;
  assign n6909 = n6858 ^ n6824 ^ n1885 ;
  assign n6910 = n6858 & n6909 ;
  assign n6911 = n6910 ^ n6679 ^ n6506 ;
  assign n6912 = n6858 ^ n6828 ^ n1534 ;
  assign n6913 = n6858 & n6912 ;
  assign n6914 = n6913 ^ n6682 ^ n6449 ;
  assign n6915 = n6858 ^ n6830 ^ n1318 ;
  assign n6916 = n6858 & n6915 ;
  assign n6917 = n6916 ^ n6685 ^ n6452 ;
  assign n6918 = n6858 ^ n6832 ^ n1118 ;
  assign n6919 = n6858 & n6918 ;
  assign n6920 = n6919 ^ n6688 ^ n6521 ;
  assign n6921 = n6858 ^ n6838 ^ n640 ;
  assign n6922 = n6858 & n6921 ;
  assign n6923 = n6922 ^ n6759 ^ n6458 ;
  assign n6924 = n6858 ^ n6841 ^ n458 ;
  assign n6925 = n6858 & n6924 ;
  assign n6926 = n6925 ^ n6727 ^ n6536 ;
  assign n6927 = n6858 ^ n6842 ^ n399 ;
  assign n6928 = n6858 & n6927 ;
  assign n6929 = n6928 ^ n6757 ^ n6539 ;
  assign n6930 = n6858 ^ n6843 ^ n345 ;
  assign n6931 = n6858 & n6930 ;
  assign n6932 = n6931 ^ n6697 ^ n6542 ;
  assign n6933 = n6858 ^ n6844 ^ n302 ;
  assign n6934 = n6858 & n6933 ;
  assign n6935 = n6934 ^ n6700 ^ n6464 ;
  assign n6936 = n6858 ^ n6795 ^ n5743 ;
  assign n6937 = n6858 & n6936 ;
  assign n6938 = n6937 ^ n6752 ^ n6556 ;
  assign n6939 = n6858 ^ n6802 ^ n4534 ;
  assign n6940 = n6858 & n6939 ;
  assign n6941 = n6940 ^ n6664 ^ n6488 ;
  assign n6942 = n6858 ^ n6806 ^ n3986 ;
  assign n6943 = n6858 & n6942 ;
  assign n6944 = n6943 ^ n6742 ^ n6518 ;
  assign n6945 = n6808 ^ n3631 ^ 1'b0 ;
  assign n6946 = n6858 & n6945 ;
  assign n6947 = n6946 ^ n6858 ^ n6641 ;
  assign n6948 = n6810 ^ n3302 ^ 1'b0 ;
  assign n6949 = n6858 & n6948 ;
  assign n6950 = n6949 ^ n6858 ^ n6643 ;
  assign n6951 = n6858 ^ n6811 ^ n3141 ;
  assign n6952 = n6858 & n6951 ;
  assign n6953 = n6952 ^ n6667 ^ n6500 ;
  assign n6954 = n6816 ^ n2404 ^ 1'b0 ;
  assign n6955 = n6858 & n6954 ;
  assign n6956 = n6955 ^ n6858 ^ n6645 ;
  assign n6957 = n6858 ^ n6820 ^ n2269 ;
  assign n6958 = n6858 & n6957 ;
  assign n6959 = n6958 ^ n6673 ^ n6443 ;
  assign n6960 = n6831 ^ n1220 ^ 1'b0 ;
  assign n6961 = n6858 & n6960 ;
  assign n6962 = n6961 ^ n6858 ^ n6654 ;
  assign n6963 = n6858 ^ n6833 ^ n1034 ;
  assign n6964 = n6858 & n6963 ;
  assign n6965 = n6964 ^ n6738 ^ n6524 ;
  assign n6966 = n6858 ^ n6840 ^ n514 ;
  assign n6967 = n6858 & n6966 ;
  assign n6968 = n6967 ^ n6658 ^ n6404 ;
  assign n6969 = n6858 ^ n6846 ^ n217 ;
  assign n6970 = n6858 & n6969 ;
  assign n6971 = n6970 ^ n6729 ^ n6545 ;
  assign n6972 = n6847 ^ n179 ^ 1'b0 ;
  assign n6973 = n6858 & n6972 ;
  assign n6974 = n6973 ^ n6858 ^ n6776 ;
  assign n6975 = n6858 ^ n6848 ^ n144 ;
  assign n6976 = n6858 & n6975 ;
  assign n6977 = n6976 ^ n6755 ^ n6470 ;
  assign n6978 = x37 | x38 ;
  assign n6979 = x40 & n6858 ;
  assign n6980 = ( x40 & ~n6628 ) | ( x40 & n6978 ) | ( ~n6628 & n6978 ) ;
  assign n6981 = ( ~n6630 & n6979 ) | ( ~n6630 & n6980 ) | ( n6979 & n6980 ) ;
  assign n6982 = n6979 ^ n6858 ^ x41 ;
  assign n6983 = ~n6979 & n6981 ;
  assign n6984 = n6801 ^ n4728 ^ 1'b0 ;
  assign n6985 = n6858 & n6984 ;
  assign n6986 = x40 | n6978 ;
  assign n6987 = ( n6635 & ~n6850 ) | ( n6635 & n6858 ) | ( ~n6850 & n6858 ) ;
  assign n6988 = n6635 & ~n6850 ;
  assign n6989 = ( n6875 & n6987 ) | ( n6875 & ~n6988 ) | ( n6987 & ~n6988 ) ;
  assign n6990 = n6858 ^ n6836 ^ n785 ;
  assign n6991 = n6985 ^ n6858 ^ n6639 ;
  assign n6992 = n6839 ^ n572 ^ 1'b0 ;
  assign n6993 = n6858 & n6992 ;
  assign n6994 = n6993 ^ n6858 ^ n6772 ;
  assign n6995 = n6829 ^ n1416 ^ 1'b0 ;
  assign n6996 = n6858 & n6995 ;
  assign n6997 = n6996 ^ n6858 ^ n6652 ;
  assign n6998 = n6845 ^ n261 ^ 1'b0 ;
  assign n6999 = n6858 & n6998 ;
  assign n7000 = n6999 ^ n6858 ^ n6770 ;
  assign n7001 = n6798 ^ n5124 ^ 1'b0 ;
  assign n7002 = n6858 & n6990 ;
  assign n7003 = n6881 ^ x42 ^ 1'b0 ;
  assign n7004 = n6858 ^ n6792 ^ n6171 ;
  assign n7005 = n6858 ^ n6803 ^ n4346 ;
  assign n7006 = n6858 ^ n6826 ^ n1766 ;
  assign n7007 = n6858 & n7006 ;
  assign n7008 = ( n6630 & n6979 ) | ( n6630 & ~n6986 ) | ( n6979 & ~n6986 ) ;
  assign n7009 = n7002 ^ n6694 ^ n6530 ;
  assign n7010 = n7007 ^ n6649 ^ n6509 ;
  assign n7011 = n6858 & n7001 ;
  assign n7012 = n6858 & n7005 ;
  assign n7013 = n7011 ^ n6858 ^ n6637 ;
  assign n7014 = n6858 ^ n6834 ^ n941 ;
  assign n7015 = n6858 & n7004 ;
  assign n7016 = n6858 & n7014 ;
  assign n7017 = n7015 ^ n6756 ^ x44 ;
  assign n7018 = n7016 ^ n6744 ^ n6527 ;
  assign n7019 = n6858 ^ n6835 ^ n859 ;
  assign n7020 = ( n6850 & n6851 ) | ( n6850 & n6858 ) | ( n6851 & n6858 ) ;
  assign n7021 = n6635 & ~n7020 ;
  assign n7022 = n7021 ^ n7020 ^ n6851 ;
  assign n7023 = n6858 & n7019 ;
  assign n7024 = n6837 ^ n716 ^ 1'b0 ;
  assign n7025 = n6858 & n7024 ;
  assign n7026 = n7012 ^ n6733 ^ n6491 ;
  assign n7027 = n7025 ^ n6858 ^ n6656 ;
  assign n7028 = n7023 ^ n6691 ^ n6455 ;
  assign n7029 = n6635 & ~n6858 ;
  assign n7030 = n6983 | n7008 ;
  assign n7031 = n6982 | n6983 ;
  assign n7032 = ~n7008 & n7031 ;
  assign n7033 = ( ~n6401 & n7003 ) | ( ~n6401 & n7032 ) | ( n7003 & n7032 ) ;
  assign n7034 = ( ~n6171 & n6863 ) | ( ~n6171 & n7033 ) | ( n6863 & n7033 ) ;
  assign n7035 = ( ~n5964 & n7017 ) | ( ~n5964 & n7034 ) | ( n7017 & n7034 ) ;
  assign n7036 = ( ~n5743 & n6869 ) | ( ~n5743 & n7035 ) | ( n6869 & n7035 ) ;
  assign n7037 = ( ~n5527 & n6938 ) | ( ~n5527 & n7036 ) | ( n6938 & n7036 ) ;
  assign n7038 = ( ~n5319 & n6887 ) | ( ~n5319 & n7037 ) | ( n6887 & n7037 ) ;
  assign n7039 = ( ~n5124 & n6878 ) | ( ~n5124 & n7038 ) | ( n6878 & n7038 ) ;
  assign n7040 = ( ~n4915 & n7013 ) | ( ~n4915 & n7039 ) | ( n7013 & n7039 ) ;
  assign n7041 = ( ~n4728 & n6886 ) | ( ~n4728 & n7040 ) | ( n6886 & n7040 ) ;
  assign n7042 = ( ~n4534 & n6991 ) | ( ~n4534 & n7041 ) | ( n6991 & n7041 ) ;
  assign n7043 = ( ~n4346 & n6941 ) | ( ~n4346 & n7042 ) | ( n6941 & n7042 ) ;
  assign n7044 = ( ~n4167 & n7026 ) | ( ~n4167 & n7043 ) | ( n7026 & n7043 ) ;
  assign n7045 = ( ~n3986 & n6890 ) | ( ~n3986 & n7044 ) | ( n6890 & n7044 ) ;
  assign n7046 = ( ~n3804 & n6944 ) | ( ~n3804 & n7045 ) | ( n6944 & n7045 ) ;
  assign n7047 = ( ~n3631 & n6883 ) | ( ~n3631 & n7046 ) | ( n6883 & n7046 ) ;
  assign n7048 = ( ~n3464 & n6947 ) | ( ~n3464 & n7047 ) | ( n6947 & n7047 ) ;
  assign n7049 = ( ~n3302 & n6884 ) | ( ~n3302 & n7048 ) | ( n6884 & n7048 ) ;
  assign n7050 = ( ~n3141 & n6950 ) | ( ~n3141 & n7049 ) | ( n6950 & n7049 ) ;
  assign n7051 = ( ~n2995 & n6953 ) | ( ~n2995 & n7050 ) | ( n6953 & n7050 ) ;
  assign n7052 = ( ~n2839 & n6893 ) | ( ~n2839 & n7051 ) | ( n6893 & n7051 ) ;
  assign n7053 = ( ~n2690 & n6906 ) | ( ~n2690 & n7052 ) | ( n6906 & n7052 ) ;
  assign n7054 = ( ~n2544 & n6898 ) | ( ~n2544 & n7053 ) | ( n6898 & n7053 ) ;
  assign n7055 = ( ~n2404 & n6901 ) | ( ~n2404 & n7054 ) | ( n6901 & n7054 ) ;
  assign n7056 = ( ~n2269 & n6956 ) | ( ~n2269 & n7055 ) | ( n6956 & n7055 ) ;
  assign n7057 = ( ~n2139 & n6959 ) | ( ~n2139 & n7056 ) | ( n6959 & n7056 ) ;
  assign n7058 = ( ~n2009 & n6904 ) | ( ~n2009 & n7057 ) | ( n6904 & n7057 ) ;
  assign n7059 = ( ~n1885 & n6908 ) | ( ~n1885 & n7058 ) | ( n6908 & n7058 ) ;
  assign n7060 = ( ~n1766 & n6911 ) | ( ~n1766 & n7059 ) | ( n6911 & n7059 ) ;
  assign n7061 = ( ~n1652 & n7010 ) | ( ~n1652 & n7060 ) | ( n7010 & n7060 ) ;
  assign n7062 = ( ~n1534 & n6885 ) | ( ~n1534 & n7061 ) | ( n6885 & n7061 ) ;
  assign n7063 = ( ~n1416 & n6914 ) | ( ~n1416 & n7062 ) | ( n6914 & n7062 ) ;
  assign n7064 = ( ~n1318 & n6997 ) | ( ~n1318 & n7063 ) | ( n6997 & n7063 ) ;
  assign n7065 = ( ~n1220 & n6917 ) | ( ~n1220 & n7064 ) | ( n6917 & n7064 ) ;
  assign n7066 = ( ~n1118 & n6962 ) | ( ~n1118 & n7065 ) | ( n6962 & n7065 ) ;
  assign n7067 = ( ~n1034 & n6920 ) | ( ~n1034 & n7066 ) | ( n6920 & n7066 ) ;
  assign n7068 = ( ~n941 & n6965 ) | ( ~n941 & n7067 ) | ( n6965 & n7067 ) ;
  assign n7069 = ( ~n859 & n7018 ) | ( ~n859 & n7068 ) | ( n7018 & n7068 ) ;
  assign n7070 = ( ~n785 & n7028 ) | ( ~n785 & n7069 ) | ( n7028 & n7069 ) ;
  assign n7071 = ( ~n716 & n7009 ) | ( ~n716 & n7070 ) | ( n7009 & n7070 ) ;
  assign n7072 = ( ~n640 & n7027 ) | ( ~n640 & n7071 ) | ( n7027 & n7071 ) ;
  assign n7073 = ( ~n572 & n6923 ) | ( ~n572 & n7072 ) | ( n6923 & n7072 ) ;
  assign n7074 = ( ~n514 & n6994 ) | ( ~n514 & n7073 ) | ( n6994 & n7073 ) ;
  assign n7075 = ( ~n458 & n6968 ) | ( ~n458 & n7074 ) | ( n6968 & n7074 ) ;
  assign n7076 = ( ~n399 & n6926 ) | ( ~n399 & n7075 ) | ( n6926 & n7075 ) ;
  assign n7077 = ( ~n345 & n6929 ) | ( ~n345 & n7076 ) | ( n6929 & n7076 ) ;
  assign n7078 = ( ~n302 & n6932 ) | ( ~n302 & n7077 ) | ( n6932 & n7077 ) ;
  assign n7079 = ( ~n261 & n6935 ) | ( ~n261 & n7078 ) | ( n6935 & n7078 ) ;
  assign n7080 = ( ~n217 & n7000 ) | ( ~n217 & n7079 ) | ( n7000 & n7079 ) ;
  assign n7081 = ( ~n179 & n6971 ) | ( ~n179 & n7080 ) | ( n6971 & n7080 ) ;
  assign n7082 = ( ~n144 & n6974 ) | ( ~n144 & n7081 ) | ( n6974 & n7081 ) ;
  assign n7083 = ( ~n134 & n6977 ) | ( ~n134 & n7082 ) | ( n6977 & n7082 ) ;
  assign n7084 = ( ~x30 & n6989 ) | ( ~x30 & n7083 ) | ( n6989 & n7083 ) ;
  assign n7085 = n6875 & n7083 ;
  assign n7086 = ~n136 & n7084 ;
  assign n7087 = n7022 | n7085 ;
  assign n7088 = n7086 | n7087 ;
  assign n7089 = n7029 | n7088 ;
  assign n7090 = n7089 ^ n7082 ^ n134 ;
  assign n7091 = n7089 & n7090 ;
  assign n7092 = n7091 ^ n6976 ^ n6763 ;
  assign n7093 = n7030 & n7089 ;
  assign n7094 = n7093 ^ n7089 ^ n6982 ;
  assign n7095 = n7089 ^ n7061 ^ n1534 ;
  assign n7096 = n7089 & n7095 ;
  assign n7097 = n7096 ^ n6882 ^ n6750 ;
  assign n7098 = n7089 ^ n7072 ^ n572 ;
  assign n7099 = n7089 & n7098 ;
  assign n7100 = n7099 ^ n6922 ^ n6761 ;
  assign n7101 = n7089 ^ n7080 ^ n179 ;
  assign n7102 = n7089 & n7101 ;
  assign n7103 = n7102 ^ n6970 ^ n6730 ;
  assign n7104 = n7089 ^ n7052 ^ n2690 ;
  assign n7105 = n7089 & n7104 ;
  assign n7106 = n7105 ^ n6895 ^ n6671 ;
  assign n7107 = n7089 ^ n7059 ^ n1766 ;
  assign n7108 = n7089 & n7107 ;
  assign n7109 = n7108 ^ n6910 ^ n6680 ;
  assign n7110 = n7063 ^ n1318 ^ 1'b0 ;
  assign n7111 = n7089 & n7110 ;
  assign n7112 = n7111 ^ n7089 ^ n6997 ;
  assign n7113 = n7089 ^ n7064 ^ n1220 ;
  assign n7114 = n7089 & n7113 ;
  assign n7115 = n7114 ^ n6916 ^ n6686 ;
  assign n7116 = n7089 ^ n7069 ^ n785 ;
  assign n7117 = n7089 & n7116 ;
  assign n7118 = n7117 ^ n7023 ^ n6692 ;
  assign n7119 = n7089 ^ n7070 ^ n716 ;
  assign n7120 = n7089 & n7119 ;
  assign n7121 = n7120 ^ n7002 ^ n6695 ;
  assign n7122 = n7071 ^ n640 ^ 1'b0 ;
  assign n7123 = n7089 & n7122 ;
  assign n7124 = n7123 ^ n7089 ^ n7027 ;
  assign n7125 = n7073 ^ n514 ^ 1'b0 ;
  assign n7126 = n7089 & n7125 ;
  assign n7127 = n7126 ^ n7089 ^ n6994 ;
  assign n7128 = n7089 ^ n7074 ^ n458 ;
  assign n7129 = n7089 & n7128 ;
  assign n7130 = n7129 ^ n6967 ^ n6659 ;
  assign n7131 = n7089 ^ n7075 ^ n399 ;
  assign n7132 = n7089 & n7131 ;
  assign n7133 = n7132 ^ n6925 ^ n6728 ;
  assign n7134 = n7089 ^ n7076 ^ n345 ;
  assign n7135 = n7089 & n7134 ;
  assign n7136 = n7135 ^ n6928 ^ n6758 ;
  assign n7137 = n7089 ^ n7077 ^ n302 ;
  assign n7138 = n7089 & n7137 ;
  assign n7139 = n7138 ^ n6931 ^ n6698 ;
  assign n7140 = n7089 ^ n7078 ^ n261 ;
  assign n7141 = n7089 & n7140 ;
  assign n7142 = n7141 ^ n6934 ^ n6701 ;
  assign n7143 = n7081 ^ n144 ^ 1'b0 ;
  assign n7144 = n7089 & n7143 ;
  assign n7145 = n7144 ^ n7089 ^ n6974 ;
  assign n7146 = n7089 ^ n7068 ^ n859 ;
  assign n7147 = n7089 ^ n7037 ^ n5319 ;
  assign n7148 = n7049 ^ n3141 ^ 1'b0 ;
  assign n7149 = n7089 & n7147 ;
  assign n7150 = n7089 ^ n7035 ^ n5743 ;
  assign n7151 = n7089 ^ n7034 ^ n5964 ;
  assign n7152 = n7089 ^ n7056 ^ n2139 ;
  assign n7153 = n7089 ^ n7053 ^ n2544 ;
  assign n7154 = n7089 ^ n7046 ^ n3631 ;
  assign n7155 = n7089 ^ n7058 ^ n1885 ;
  assign n7156 = n7089 ^ n7062 ^ n1416 ;
  assign n7157 = n7089 ^ n7045 ^ n3804 ;
  assign n7158 = n7089 ^ n7044 ^ n3986 ;
  assign n7159 = n7089 ^ n7067 ^ n941 ;
  assign n7160 = n7089 ^ n7066 ^ n1034 ;
  assign n7161 = n7149 ^ n6872 ^ n6775 ;
  assign n7162 = n7089 & n7150 ;
  assign n7163 = ( x37 & n6856 ) | ( x37 & n7089 ) | ( n6856 & n7089 ) ;
  assign n7164 = ( n6855 & ~n6856 ) | ( n6855 & n7163 ) | ( ~n6856 & n7163 ) ;
  assign n7165 = n7089 ^ n7042 ^ n4346 ;
  assign n7166 = n7089 ^ n7054 ^ n2404 ;
  assign n7167 = n7089 ^ n7050 ^ n2995 ;
  assign n7168 = n7089 ^ n7051 ^ n2839 ;
  assign n7169 = n7089 ^ n7048 ^ n3302 ;
  assign n7170 = n7089 ^ n7038 ^ n5124 ;
  assign n7171 = n7089 ^ n7043 ^ n4167 ;
  assign n7172 = n7089 ^ n7040 ^ n4728 ;
  assign n7173 = n7089 & n7155 ;
  assign n7174 = n7089 ^ n7060 ^ n1652 ;
  assign n7175 = n7162 ^ n6861 ^ n6725 ;
  assign n7176 = ~n7163 & n7164 ;
  assign n7177 = n7089 & n7151 ;
  assign n7178 = n7089 & n7166 ;
  assign n7179 = n7178 ^ n6900 ^ n6741 ;
  assign n7180 = n7089 & n7167 ;
  assign n7181 = n7180 ^ n6952 ^ n6668 ;
  assign n7182 = n7177 ^ n7015 ^ n6777 ;
  assign n7183 = n7089 & n7158 ;
  assign n7184 = n7183 ^ n6889 ^ n6762 ;
  assign n7185 = n7089 & n7174 ;
  assign n7186 = n7185 ^ n7007 ^ n6650 ;
  assign n7187 = n7089 & n7156 ;
  assign n7188 = n7187 ^ n6913 ^ n6683 ;
  assign n7189 = n7089 & n7168 ;
  assign n7190 = n7189 ^ n6892 ^ n6769 ;
  assign n7191 = n7089 & n7165 ;
  assign n7192 = n7191 ^ n6940 ^ n6665 ;
  assign n7193 = n7089 & n7171 ;
  assign n7194 = n7089 & n7157 ;
  assign n7195 = n7193 ^ n7012 ^ n6735 ;
  assign n7196 = n7194 ^ n6943 ^ n6743 ;
  assign n7197 = n7089 & n7172 ;
  assign n7198 = n7089 & n7169 ;
  assign n7199 = n7198 ^ n6879 ^ n6732 ;
  assign n7200 = n7089 ^ n7036 ^ n5527 ;
  assign n7201 = n7197 ^ n6864 ^ n6662 ;
  assign n7202 = n7089 & n7159 ;
  assign n7203 = n7089 & n7152 ;
  assign n7204 = n7203 ^ n6958 ^ n6674 ;
  assign n7205 = n7202 ^ n6964 ^ n6739 ;
  assign n7206 = n7089 & n7170 ;
  assign n7207 = n7206 ^ n6877 ^ n6726 ;
  assign n7208 = n7089 & n7154 ;
  assign n7209 = n7208 ^ n6874 ^ n6766 ;
  assign n7210 = n7089 & n7200 ;
  assign n7211 = n7210 ^ n6937 ^ n6753 ;
  assign n7212 = n7089 & n7148 ;
  assign n7213 = n7212 ^ n7089 ^ n6950 ;
  assign n7214 = n7089 & n7146 ;
  assign n7215 = n7089 & n7160 ;
  assign n7216 = n7089 & n7153 ;
  assign n7217 = n7214 ^ n7016 ^ n6745 ;
  assign n7218 = n7216 ^ n6897 ^ n6748 ;
  assign n7219 = n7215 ^ n6919 ^ n6689 ;
  assign n7220 = ~x37 & n7089 ;
  assign n7221 = n7065 ^ n1118 ^ 1'b0 ;
  assign n7222 = n7079 ^ n217 ^ 1'b0 ;
  assign n7223 = n7220 ^ x38 ^ 1'b0 ;
  assign n7224 = n7176 | n7223 ;
  assign n7225 = n7089 & n7222 ;
  assign n7226 = n7225 ^ n7089 ^ n7000 ;
  assign n7227 = n7089 & n7221 ;
  assign n7228 = n6858 & ~n7088 ;
  assign n7229 = n7041 ^ n4534 ^ 1'b0 ;
  assign n7230 = n6978 & n7089 ;
  assign n7231 = n7089 & n7229 ;
  assign n7232 = ( n7089 & n7228 ) | ( n7089 & ~n7230 ) | ( n7228 & ~n7230 ) ;
  assign n7233 = ( ~x37 & n6858 ) | ( ~x37 & n7089 ) | ( n6858 & n7089 ) ;
  assign n7234 = n7173 ^ n6907 ^ n6677 ;
  assign n7235 = n7231 ^ n7089 ^ n6991 ;
  assign n7236 = ( x33 & x34 ) | ( x33 & ~n7029 ) | ( x34 & ~n7029 ) ;
  assign n7237 = n7047 ^ n3464 ^ 1'b0 ;
  assign n7238 = x35 | x36 ;
  assign n7239 = n7227 ^ n7089 ^ n6962 ;
  assign n7240 = ( x37 & n6858 ) | ( x37 & ~n7238 ) | ( n6858 & ~n7238 ) ;
  assign n7241 = ( x35 & ~n7029 ) | ( x35 & n7236 ) | ( ~n7029 & n7236 ) ;
  assign n7242 = n7089 & n7237 ;
  assign n7243 = n7089 ^ n7032 ^ n6401 ;
  assign n7244 = n7233 & n7240 ;
  assign n7245 = n7224 & ~n7244 ;
  assign n7246 = n7029 | n7085 ;
  assign n7247 = n7242 ^ n7089 ^ n6947 ;
  assign n7248 = n7039 ^ n4915 ^ 1'b0 ;
  assign n7249 = n7089 & n7248 ;
  assign n7250 = ( ~n7022 & n7241 ) | ( ~n7022 & n7246 ) | ( n7241 & n7246 ) ;
  assign n7251 = ~n7246 & n7250 ;
  assign n7252 = n7232 ^ x40 ^ 1'b0 ;
  assign n7253 = ( ~n6630 & n7245 ) | ( ~n6630 & n7252 ) | ( n7245 & n7252 ) ;
  assign n7254 = n7249 ^ n7089 ^ n7013 ;
  assign n7255 = ( n136 & n6875 ) | ( n136 & n7083 ) | ( n6875 & n7083 ) ;
  assign n7256 = n7089 & n7243 ;
  assign n7257 = ( n6875 & n7022 ) | ( n6875 & ~n7029 ) | ( n7022 & ~n7029 ) ;
  assign n7258 = ( ~n6875 & n7083 ) | ( ~n6875 & n7089 ) | ( n7083 & n7089 ) ;
  assign n7259 = n7055 ^ n2269 ^ 1'b0 ;
  assign n7260 = n7256 ^ n6881 ^ x42 ;
  assign n7261 = ( n7083 & n7085 ) | ( n7083 & ~n7089 ) | ( n7085 & ~n7089 ) ;
  assign n7262 = n7255 & ~n7261 ;
  assign n7263 = ~n6875 & n7083 ;
  assign n7264 = n7057 ^ n2009 ^ 1'b0 ;
  assign n7265 = n7089 & n7264 ;
  assign n7266 = ~n7088 & n7257 ;
  assign n7267 = n7033 ^ n6171 ^ 1'b0 ;
  assign n7268 = n7089 & n7267 ;
  assign n7269 = ( ~n6401 & n7094 ) | ( ~n6401 & n7253 ) | ( n7094 & n7253 ) ;
  assign n7270 = n7268 ^ n7089 ^ n6863 ;
  assign n7271 = ( n7092 & n7258 ) | ( n7092 & ~n7263 ) | ( n7258 & ~n7263 ) ;
  assign n7272 = n7089 & n7259 ;
  assign n7273 = n7272 ^ n7089 ^ n6956 ;
  assign n7274 = n7265 ^ n7089 ^ n6904 ;
  assign n7275 = ( ~n6171 & n7260 ) | ( ~n6171 & n7269 ) | ( n7260 & n7269 ) ;
  assign n7276 = ( ~n5964 & n7270 ) | ( ~n5964 & n7275 ) | ( n7270 & n7275 ) ;
  assign n7277 = n7275 ^ n5964 ^ 1'b0 ;
  assign n7278 = ( ~n5743 & n7182 ) | ( ~n5743 & n7276 ) | ( n7182 & n7276 ) ;
  assign n7279 = ( ~n5527 & n7175 ) | ( ~n5527 & n7278 ) | ( n7175 & n7278 ) ;
  assign n7280 = ( ~n5319 & n7211 ) | ( ~n5319 & n7279 ) | ( n7211 & n7279 ) ;
  assign n7281 = ( ~n5124 & n7161 ) | ( ~n5124 & n7280 ) | ( n7161 & n7280 ) ;
  assign n7282 = ( ~n4915 & n7207 ) | ( ~n4915 & n7281 ) | ( n7207 & n7281 ) ;
  assign n7283 = ( ~n4728 & n7254 ) | ( ~n4728 & n7282 ) | ( n7254 & n7282 ) ;
  assign n7284 = ( ~n4534 & n7201 ) | ( ~n4534 & n7283 ) | ( n7201 & n7283 ) ;
  assign n7285 = ( ~n4346 & n7235 ) | ( ~n4346 & n7284 ) | ( n7235 & n7284 ) ;
  assign n7286 = ( ~n4167 & n7192 ) | ( ~n4167 & n7285 ) | ( n7192 & n7285 ) ;
  assign n7287 = ( ~n3986 & n7195 ) | ( ~n3986 & n7286 ) | ( n7195 & n7286 ) ;
  assign n7288 = ( ~n3804 & n7184 ) | ( ~n3804 & n7287 ) | ( n7184 & n7287 ) ;
  assign n7289 = ( ~n3631 & n7196 ) | ( ~n3631 & n7288 ) | ( n7196 & n7288 ) ;
  assign n7290 = ( ~n3464 & n7209 ) | ( ~n3464 & n7289 ) | ( n7209 & n7289 ) ;
  assign n7291 = ( ~n3302 & n7247 ) | ( ~n3302 & n7290 ) | ( n7247 & n7290 ) ;
  assign n7292 = ( ~n3141 & n7199 ) | ( ~n3141 & n7291 ) | ( n7199 & n7291 ) ;
  assign n7293 = ( ~n2995 & n7213 ) | ( ~n2995 & n7292 ) | ( n7213 & n7292 ) ;
  assign n7294 = ( ~n2839 & n7181 ) | ( ~n2839 & n7293 ) | ( n7181 & n7293 ) ;
  assign n7295 = ( ~n2690 & n7190 ) | ( ~n2690 & n7294 ) | ( n7190 & n7294 ) ;
  assign n7296 = ( ~n2544 & n7106 ) | ( ~n2544 & n7295 ) | ( n7106 & n7295 ) ;
  assign n7297 = ( ~n2404 & n7218 ) | ( ~n2404 & n7296 ) | ( n7218 & n7296 ) ;
  assign n7298 = ( ~n2269 & n7179 ) | ( ~n2269 & n7297 ) | ( n7179 & n7297 ) ;
  assign n7299 = ( ~n2139 & n7273 ) | ( ~n2139 & n7298 ) | ( n7273 & n7298 ) ;
  assign n7300 = ( ~n2009 & n7204 ) | ( ~n2009 & n7299 ) | ( n7204 & n7299 ) ;
  assign n7301 = ( ~n1885 & n7274 ) | ( ~n1885 & n7300 ) | ( n7274 & n7300 ) ;
  assign n7302 = ( ~n1766 & n7234 ) | ( ~n1766 & n7301 ) | ( n7234 & n7301 ) ;
  assign n7303 = ( ~n1652 & n7109 ) | ( ~n1652 & n7302 ) | ( n7109 & n7302 ) ;
  assign n7304 = ( ~n1534 & n7186 ) | ( ~n1534 & n7303 ) | ( n7186 & n7303 ) ;
  assign n7305 = ( ~n1416 & n7097 ) | ( ~n1416 & n7304 ) | ( n7097 & n7304 ) ;
  assign n7306 = ( ~n1318 & n7188 ) | ( ~n1318 & n7305 ) | ( n7188 & n7305 ) ;
  assign n7307 = ( ~n1220 & n7112 ) | ( ~n1220 & n7306 ) | ( n7112 & n7306 ) ;
  assign n7308 = ( ~n1118 & n7115 ) | ( ~n1118 & n7307 ) | ( n7115 & n7307 ) ;
  assign n7309 = ( ~n1034 & n7239 ) | ( ~n1034 & n7308 ) | ( n7239 & n7308 ) ;
  assign n7310 = ( ~n941 & n7219 ) | ( ~n941 & n7309 ) | ( n7219 & n7309 ) ;
  assign n7311 = ( ~n859 & n7205 ) | ( ~n859 & n7310 ) | ( n7205 & n7310 ) ;
  assign n7312 = ( ~n785 & n7217 ) | ( ~n785 & n7311 ) | ( n7217 & n7311 ) ;
  assign n7313 = ( ~n716 & n7118 ) | ( ~n716 & n7312 ) | ( n7118 & n7312 ) ;
  assign n7314 = ( ~n640 & n7121 ) | ( ~n640 & n7313 ) | ( n7121 & n7313 ) ;
  assign n7315 = n7314 ^ n572 ^ 1'b0 ;
  assign n7316 = ( ~n572 & n7124 ) | ( ~n572 & n7314 ) | ( n7124 & n7314 ) ;
  assign n7317 = ( ~n514 & n7100 ) | ( ~n514 & n7316 ) | ( n7100 & n7316 ) ;
  assign n7318 = n7317 ^ n458 ^ 1'b0 ;
  assign n7319 = ( ~n458 & n7127 ) | ( ~n458 & n7317 ) | ( n7127 & n7317 ) ;
  assign n7320 = n7298 ^ n2139 ^ 1'b0 ;
  assign n7321 = n7300 ^ n1885 ^ 1'b0 ;
  assign n7322 = n7306 ^ n1220 ^ 1'b0 ;
  assign n7323 = n7308 ^ n1034 ^ 1'b0 ;
  assign n7324 = ( ~n399 & n7130 ) | ( ~n399 & n7319 ) | ( n7130 & n7319 ) ;
  assign n7325 = ( ~n345 & n7133 ) | ( ~n345 & n7324 ) | ( n7133 & n7324 ) ;
  assign n7326 = ( ~n302 & n7136 ) | ( ~n302 & n7325 ) | ( n7136 & n7325 ) ;
  assign n7327 = ( ~n261 & n7139 ) | ( ~n261 & n7326 ) | ( n7139 & n7326 ) ;
  assign n7328 = ( ~n217 & n7142 ) | ( ~n217 & n7327 ) | ( n7142 & n7327 ) ;
  assign n7329 = ( ~n179 & n7226 ) | ( ~n179 & n7328 ) | ( n7226 & n7328 ) ;
  assign n7330 = ( ~n144 & n7103 ) | ( ~n144 & n7329 ) | ( n7103 & n7329 ) ;
  assign n7331 = ( ~n134 & n7145 ) | ( ~n134 & n7330 ) | ( n7145 & n7330 ) ;
  assign n7332 = n7092 & n7331 ;
  assign n7333 = ( ~x30 & n7271 ) | ( ~x30 & n7331 ) | ( n7271 & n7331 ) ;
  assign n7334 = ~n136 & n7333 ;
  assign n7335 = n7332 | n7334 ;
  assign n7336 = n7262 | n7335 ;
  assign n7337 = n7266 | n7336 ;
  assign n7338 = ( n7176 & ~n7244 ) | ( n7176 & n7337 ) | ( ~n7244 & n7337 ) ;
  assign n7339 = ~n7176 & n7338 ;
  assign n7340 = n7277 & n7337 ;
  assign n7341 = n7340 ^ n7337 ^ n7270 ;
  assign n7342 = n7337 ^ n7279 ^ n5319 ;
  assign n7343 = n7337 & n7342 ;
  assign n7344 = n7343 ^ n7210 ^ n6938 ;
  assign n7345 = n7337 ^ n7281 ^ n4915 ;
  assign n7346 = n7337 & n7345 ;
  assign n7347 = n7346 ^ n7206 ^ n6878 ;
  assign n7348 = n7320 & n7337 ;
  assign n7349 = n7348 ^ n7337 ^ n7273 ;
  assign n7350 = n7321 & n7337 ;
  assign n7351 = n7350 ^ n7337 ^ n7274 ;
  assign n7352 = n7322 & n7337 ;
  assign n7353 = n7352 ^ n7337 ^ n7112 ;
  assign n7354 = n7323 & n7337 ;
  assign n7355 = n7354 ^ n7337 ^ n7239 ;
  assign n7356 = n7315 & n7337 ;
  assign n7357 = n7356 ^ n7337 ^ n7124 ;
  assign n7358 = n7337 ^ n7316 ^ n514 ;
  assign n7359 = n7337 & n7358 ;
  assign n7360 = n7359 ^ n7099 ^ n6923 ;
  assign n7361 = n7318 & n7337 ;
  assign n7362 = n7361 ^ n7337 ^ n7127 ;
  assign n7363 = n7337 ^ n7324 ^ n345 ;
  assign n7364 = n7337 & n7363 ;
  assign n7365 = n7364 ^ n7132 ^ n6926 ;
  assign n7366 = n7337 ^ n7327 ^ n217 ;
  assign n7367 = n7337 & n7366 ;
  assign n7368 = n7367 ^ n7141 ^ n6935 ;
  assign n7369 = n7328 ^ n179 ^ 1'b0 ;
  assign n7370 = n7337 & n7369 ;
  assign n7371 = n7370 ^ n7337 ^ n7226 ;
  assign n7372 = n7337 ^ n7329 ^ n144 ;
  assign n7373 = ~n7238 & n7337 ;
  assign n7374 = ( n7262 & n7266 ) | ( n7262 & ~n7373 ) | ( n7266 & ~n7373 ) ;
  assign n7375 = n7089 & ~n7335 ;
  assign n7376 = n7373 | n7375 ;
  assign n7377 = ( n7373 & ~n7374 ) | ( n7373 & n7376 ) | ( ~n7374 & n7376 ) ;
  assign n7378 = ( x35 & n7086 ) | ( x35 & n7337 ) | ( n7086 & n7337 ) ;
  assign n7379 = ( ~n7086 & n7251 ) | ( ~n7086 & n7378 ) | ( n7251 & n7378 ) ;
  assign n7380 = ~n7378 & n7379 ;
  assign n7381 = n7337 ^ n7280 ^ n5124 ;
  assign n7382 = n7337 & n7381 ;
  assign n7383 = n7382 ^ n7149 ^ n6887 ;
  assign n7384 = n7337 ^ n7283 ^ n4534 ;
  assign n7385 = n7337 & n7384 ;
  assign n7386 = n7385 ^ n7197 ^ n6886 ;
  assign n7387 = n7284 ^ n4346 ^ 1'b0 ;
  assign n7388 = n7337 & n7387 ;
  assign n7389 = n7337 ^ n7285 ^ n4167 ;
  assign n7390 = n7337 & n7389 ;
  assign n7391 = n7337 ^ n7287 ^ n3804 ;
  assign n7392 = n7337 & n7391 ;
  assign n7393 = n7392 ^ n7183 ^ n6890 ;
  assign n7394 = n7337 ^ n7291 ^ n3141 ;
  assign n7395 = n7337 & n7394 ;
  assign n7396 = n7395 ^ n7198 ^ n6884 ;
  assign n7397 = n7337 ^ n7293 ^ n2839 ;
  assign n7398 = n7337 & n7397 ;
  assign n7399 = n7390 ^ n7191 ^ n6941 ;
  assign n7400 = n7398 ^ n7180 ^ n6953 ;
  assign n7401 = n7337 ^ n7294 ^ n2690 ;
  assign n7402 = n7337 & n7401 ;
  assign n7403 = n7402 ^ n7189 ^ n6893 ;
  assign n7404 = n7337 ^ n7296 ^ n2404 ;
  assign n7405 = n7337 & n7404 ;
  assign n7406 = n7405 ^ n7216 ^ n6898 ;
  assign n7407 = n7337 ^ n7297 ^ n2269 ;
  assign n7408 = n7337 & n7407 ;
  assign n7409 = n7408 ^ n7178 ^ n6901 ;
  assign n7410 = n7337 ^ n7299 ^ n2009 ;
  assign n7411 = n7337 & n7410 ;
  assign n7412 = n7411 ^ n7203 ^ n6959 ;
  assign n7413 = n7337 ^ n7302 ^ n1652 ;
  assign n7414 = n7337 & n7413 ;
  assign n7415 = n7414 ^ n7108 ^ n6911 ;
  assign n7416 = n7337 ^ n7303 ^ n1534 ;
  assign n7417 = n7337 & n7416 ;
  assign n7418 = n7417 ^ n7185 ^ n7010 ;
  assign n7419 = n7337 ^ n7304 ^ n1416 ;
  assign n7420 = n7337 & n7419 ;
  assign n7421 = n7420 ^ n7096 ^ n6885 ;
  assign n7422 = n7337 ^ n7305 ^ n1318 ;
  assign n7423 = n7337 & n7422 ;
  assign n7424 = n7423 ^ n7187 ^ n6914 ;
  assign n7425 = n7337 ^ n7307 ^ n1118 ;
  assign n7426 = n7337 & n7425 ;
  assign n7427 = n7426 ^ n7114 ^ n6917 ;
  assign n7428 = n7337 ^ n7309 ^ n941 ;
  assign n7429 = n7337 & n7428 ;
  assign n7430 = n7429 ^ n7215 ^ n6920 ;
  assign n7431 = n7337 ^ n7311 ^ n785 ;
  assign n7432 = n7337 & n7431 ;
  assign n7433 = n7432 ^ n7214 ^ n7018 ;
  assign n7434 = n7337 ^ n7313 ^ n640 ;
  assign n7435 = n7337 & n7434 ;
  assign n7436 = n7435 ^ n7120 ^ n7009 ;
  assign n7437 = n7337 ^ n7319 ^ n399 ;
  assign n7438 = n7337 & n7437 ;
  assign n7439 = n7438 ^ n7129 ^ n6968 ;
  assign n7440 = n7337 ^ n7325 ^ n302 ;
  assign n7441 = n7337 & n7440 ;
  assign n7442 = n7441 ^ n7135 ^ n6929 ;
  assign n7443 = n7337 ^ n7326 ^ n261 ;
  assign n7444 = n7337 & n7443 ;
  assign n7445 = n7444 ^ n7138 ^ n6932 ;
  assign n7446 = n7337 & n7372 ;
  assign n7447 = n7446 ^ n7102 ^ n6971 ;
  assign n7448 = n7388 ^ n7337 ^ n7235 ;
  assign n7449 = n7330 ^ n134 ^ 1'b0 ;
  assign n7450 = n7337 ^ n7269 ^ n6171 ;
  assign n7451 = n7337 ^ n7289 ^ n3464 ;
  assign n7452 = n7253 ^ n6401 ^ 1'b0 ;
  assign n7453 = n7337 ^ n7301 ^ n1766 ;
  assign n7454 = n7337 ^ n7312 ^ n716 ;
  assign n7455 = n7339 ^ n7220 ^ x38 ;
  assign n7456 = n7337 ^ n7286 ^ n3986 ;
  assign n7457 = n7337 ^ n7295 ^ n2544 ;
  assign n7458 = n7337 & n7453 ;
  assign n7459 = n7292 ^ n2995 ^ 1'b0 ;
  assign n7460 = n7337 & n7450 ;
  assign n7461 = n7337 & n7459 ;
  assign n7462 = n7460 ^ n7256 ^ n7003 ;
  assign n7463 = n7461 ^ n7337 ^ n7213 ;
  assign n7464 = ~x35 & n7337 ;
  assign n7465 = n7458 ^ n7173 ^ n6908 ;
  assign n7466 = n7464 ^ x36 ^ 1'b0 ;
  assign n7467 = n7380 | n7466 ;
  assign n7468 = n7337 & n7454 ;
  assign n7469 = n7337 ^ n7310 ^ n859 ;
  assign n7470 = n7337 & n7469 ;
  assign n7471 = n7337 ^ n7278 ^ n5527 ;
  assign n7472 = n7290 ^ n3302 ^ 1'b0 ;
  assign n7473 = n7337 ^ n7288 ^ n3631 ;
  assign n7474 = n7337 & n7451 ;
  assign n7475 = n7474 ^ n7208 ^ n6883 ;
  assign n7476 = n7337 & n7472 ;
  assign n7477 = n7377 ^ x37 ^ 1'b0 ;
  assign n7478 = n7337 & n7457 ;
  assign n7479 = n7282 ^ n4728 ^ 1'b0 ;
  assign n7480 = n7337 ^ n7245 ^ n6630 ;
  assign n7481 = n7468 ^ n7117 ^ n7028 ;
  assign n7482 = n7337 ^ n7276 ^ n5743 ;
  assign n7483 = n7478 ^ n7105 ^ n6906 ;
  assign n7484 = ( ~x35 & n7089 ) | ( ~x35 & n7337 ) | ( n7089 & n7337 ) ;
  assign n7485 = ( n7331 & n7332 ) | ( n7331 & ~n7337 ) | ( n7332 & ~n7337 ) ;
  assign n7486 = n7337 & n7452 ;
  assign n7487 = n7476 ^ n7337 ^ n7247 ;
  assign n7488 = ( n136 & n7092 ) | ( n136 & n7331 ) | ( n7092 & n7331 ) ;
  assign n7489 = n7486 ^ n7337 ^ n7094 ;
  assign n7490 = n7337 & n7449 ;
  assign n7491 = n7337 & n7480 ;
  assign n7492 = x33 | x34 ;
  assign n7493 = ( x35 & n7089 ) | ( x35 & ~n7492 ) | ( n7089 & ~n7492 ) ;
  assign n7494 = n7484 & n7493 ;
  assign n7495 = n7491 ^ n7232 ^ x40 ;
  assign n7496 = n7467 & ~n7494 ;
  assign n7497 = ( ~n6858 & n7477 ) | ( ~n6858 & n7496 ) | ( n7477 & n7496 ) ;
  assign n7498 = n7490 ^ n7337 ^ n7145 ;
  assign n7499 = n7337 & n7456 ;
  assign n7500 = ( ~n6630 & n7455 ) | ( ~n6630 & n7497 ) | ( n7455 & n7497 ) ;
  assign n7501 = n7499 ^ n7193 ^ n7026 ;
  assign n7502 = n7337 & n7471 ;
  assign n7503 = ( ~n6401 & n7495 ) | ( ~n6401 & n7500 ) | ( n7495 & n7500 ) ;
  assign n7504 = n7502 ^ n7162 ^ n6869 ;
  assign n7505 = n7092 & ~n7331 ;
  assign n7506 = n7337 & n7473 ;
  assign n7507 = ( n7092 & ~n7331 ) | ( n7092 & n7337 ) | ( ~n7331 & n7337 ) ;
  assign n7508 = ( n7498 & ~n7505 ) | ( n7498 & n7507 ) | ( ~n7505 & n7507 ) ;
  assign n7509 = n7337 & n7479 ;
  assign n7510 = ( ~n6171 & n7489 ) | ( ~n6171 & n7503 ) | ( n7489 & n7503 ) ;
  assign n7511 = n7506 ^ n7194 ^ n6944 ;
  assign n7512 = ( ~n5964 & n7462 ) | ( ~n5964 & n7510 ) | ( n7462 & n7510 ) ;
  assign n7513 = n7337 & n7482 ;
  assign n7514 = n7513 ^ n7177 ^ n7017 ;
  assign n7515 = n7470 ^ n7202 ^ n6965 ;
  assign n7516 = ~n7485 & n7488 ;
  assign n7517 = ( ~n5743 & n7341 ) | ( ~n5743 & n7512 ) | ( n7341 & n7512 ) ;
  assign n7518 = n7509 ^ n7337 ^ n7254 ;
  assign n7519 = n7092 & ~n7337 ;
  assign n7520 = ( ~n5527 & n7514 ) | ( ~n5527 & n7517 ) | ( n7514 & n7517 ) ;
  assign n7521 = ( ~n5319 & n7504 ) | ( ~n5319 & n7520 ) | ( n7504 & n7520 ) ;
  assign n7522 = ( ~n5124 & n7344 ) | ( ~n5124 & n7521 ) | ( n7344 & n7521 ) ;
  assign n7523 = ( ~n4915 & n7383 ) | ( ~n4915 & n7522 ) | ( n7383 & n7522 ) ;
  assign n7524 = ( ~n4728 & n7347 ) | ( ~n4728 & n7523 ) | ( n7347 & n7523 ) ;
  assign n7525 = ( ~n4534 & n7518 ) | ( ~n4534 & n7524 ) | ( n7518 & n7524 ) ;
  assign n7526 = ( ~n4346 & n7386 ) | ( ~n4346 & n7525 ) | ( n7386 & n7525 ) ;
  assign n7527 = ( ~n4167 & n7448 ) | ( ~n4167 & n7526 ) | ( n7448 & n7526 ) ;
  assign n7528 = ( ~n3986 & n7399 ) | ( ~n3986 & n7527 ) | ( n7399 & n7527 ) ;
  assign n7529 = ( ~n3804 & n7501 ) | ( ~n3804 & n7528 ) | ( n7501 & n7528 ) ;
  assign n7530 = ( ~n3631 & n7393 ) | ( ~n3631 & n7529 ) | ( n7393 & n7529 ) ;
  assign n7531 = ( ~n3464 & n7511 ) | ( ~n3464 & n7530 ) | ( n7511 & n7530 ) ;
  assign n7532 = ( ~n3302 & n7475 ) | ( ~n3302 & n7531 ) | ( n7475 & n7531 ) ;
  assign n7533 = ( ~n3141 & n7487 ) | ( ~n3141 & n7532 ) | ( n7487 & n7532 ) ;
  assign n7534 = ( ~n2995 & n7396 ) | ( ~n2995 & n7533 ) | ( n7396 & n7533 ) ;
  assign n7535 = ( ~n2839 & n7463 ) | ( ~n2839 & n7534 ) | ( n7463 & n7534 ) ;
  assign n7536 = ( ~n2690 & n7400 ) | ( ~n2690 & n7535 ) | ( n7400 & n7535 ) ;
  assign n7537 = ( ~n2544 & n7403 ) | ( ~n2544 & n7536 ) | ( n7403 & n7536 ) ;
  assign n7538 = ( ~n2404 & n7483 ) | ( ~n2404 & n7537 ) | ( n7483 & n7537 ) ;
  assign n7539 = ( ~n2269 & n7406 ) | ( ~n2269 & n7538 ) | ( n7406 & n7538 ) ;
  assign n7540 = ( ~n2139 & n7409 ) | ( ~n2139 & n7539 ) | ( n7409 & n7539 ) ;
  assign n7541 = ( ~n2009 & n7349 ) | ( ~n2009 & n7540 ) | ( n7349 & n7540 ) ;
  assign n7542 = ( ~n1885 & n7412 ) | ( ~n1885 & n7541 ) | ( n7412 & n7541 ) ;
  assign n7543 = ( ~n1766 & n7351 ) | ( ~n1766 & n7542 ) | ( n7351 & n7542 ) ;
  assign n7544 = ( ~n1652 & n7465 ) | ( ~n1652 & n7543 ) | ( n7465 & n7543 ) ;
  assign n7545 = ( ~n1534 & n7415 ) | ( ~n1534 & n7544 ) | ( n7415 & n7544 ) ;
  assign n7546 = ( ~n1416 & n7418 ) | ( ~n1416 & n7545 ) | ( n7418 & n7545 ) ;
  assign n7547 = ( ~n1318 & n7421 ) | ( ~n1318 & n7546 ) | ( n7421 & n7546 ) ;
  assign n7548 = ( ~n1220 & n7424 ) | ( ~n1220 & n7547 ) | ( n7424 & n7547 ) ;
  assign n7549 = ( ~n1118 & n7353 ) | ( ~n1118 & n7548 ) | ( n7353 & n7548 ) ;
  assign n7550 = ( ~n1034 & n7427 ) | ( ~n1034 & n7549 ) | ( n7427 & n7549 ) ;
  assign n7551 = ( ~n941 & n7355 ) | ( ~n941 & n7550 ) | ( n7355 & n7550 ) ;
  assign n7552 = ( ~n859 & n7430 ) | ( ~n859 & n7551 ) | ( n7430 & n7551 ) ;
  assign n7553 = ( ~n785 & n7515 ) | ( ~n785 & n7552 ) | ( n7515 & n7552 ) ;
  assign n7554 = ( ~n716 & n7433 ) | ( ~n716 & n7553 ) | ( n7433 & n7553 ) ;
  assign n7555 = ( ~n640 & n7481 ) | ( ~n640 & n7554 ) | ( n7481 & n7554 ) ;
  assign n7556 = ( ~n572 & n7436 ) | ( ~n572 & n7555 ) | ( n7436 & n7555 ) ;
  assign n7557 = ( ~n514 & n7357 ) | ( ~n514 & n7556 ) | ( n7357 & n7556 ) ;
  assign n7558 = ( ~n458 & n7360 ) | ( ~n458 & n7557 ) | ( n7360 & n7557 ) ;
  assign n7559 = n7556 ^ n514 ^ 1'b0 ;
  assign n7560 = ( ~n399 & n7362 ) | ( ~n399 & n7558 ) | ( n7362 & n7558 ) ;
  assign n7561 = ( ~n345 & n7439 ) | ( ~n345 & n7560 ) | ( n7439 & n7560 ) ;
  assign n7562 = ( ~n302 & n7365 ) | ( ~n302 & n7561 ) | ( n7365 & n7561 ) ;
  assign n7563 = ( ~n261 & n7442 ) | ( ~n261 & n7562 ) | ( n7442 & n7562 ) ;
  assign n7564 = ( ~n217 & n7445 ) | ( ~n217 & n7563 ) | ( n7445 & n7563 ) ;
  assign n7565 = ( ~n179 & n7368 ) | ( ~n179 & n7564 ) | ( n7368 & n7564 ) ;
  assign n7566 = ( ~n144 & n7371 ) | ( ~n144 & n7565 ) | ( n7371 & n7565 ) ;
  assign n7567 = ( ~n134 & n7447 ) | ( ~n134 & n7566 ) | ( n7447 & n7566 ) ;
  assign n7568 = ( ~x30 & n7508 ) | ( ~x30 & n7567 ) | ( n7508 & n7567 ) ;
  assign n7569 = ~n136 & n7568 ;
  assign n7570 = ~n7498 & n7567 ;
  assign n7571 = ( n7567 & n7569 ) | ( n7567 & ~n7570 ) | ( n7569 & ~n7570 ) ;
  assign n7572 = ( n7498 & n7516 ) | ( n7498 & ~n7519 ) | ( n7516 & ~n7519 ) ;
  assign n7573 = n7565 ^ n144 ^ 1'b0 ;
  assign n7574 = n7516 | n7571 ;
  assign n7575 = n7519 | n7574 ;
  assign n7576 = n7575 ^ n7564 ^ n179 ;
  assign n7577 = n7573 & n7575 ;
  assign n7578 = n7575 & n7576 ;
  assign n7579 = ( n7380 & ~n7494 ) | ( n7380 & n7575 ) | ( ~n7494 & n7575 ) ;
  assign n7580 = ~n7380 & n7579 ;
  assign n7581 = n7575 ^ n7555 ^ n572 ;
  assign n7582 = n7559 & n7575 ;
  assign n7583 = n7582 ^ n7575 ^ n7357 ;
  assign n7584 = n7577 ^ n7575 ^ n7371 ;
  assign n7585 = n7575 ^ n7563 ^ n217 ;
  assign n7586 = n7575 ^ n7562 ^ n261 ;
  assign n7587 = n7575 ^ n7561 ^ n302 ;
  assign n7588 = n7575 & n7587 ;
  assign n7589 = n7575 & n7585 ;
  assign n7590 = n7575 & n7586 ;
  assign n7591 = n7575 ^ n7560 ^ n345 ;
  assign n7592 = n7575 & n7591 ;
  assign n7593 = n7575 ^ n7566 ^ n134 ;
  assign n7594 = n7575 ^ n7553 ^ n716 ;
  assign n7595 = n7575 ^ n7557 ^ n458 ;
  assign n7596 = n7575 & n7593 ;
  assign n7597 = n7575 & n7581 ;
  assign n7598 = n7575 & n7594 ;
  assign n7599 = n7575 & n7595 ;
  assign n7600 = n7597 ^ n7435 ^ n7121 ;
  assign n7601 = n7592 ^ n7438 ^ n7130 ;
  assign n7602 = n7598 ^ n7432 ^ n7217 ;
  assign n7603 = n7589 ^ n7444 ^ n7139 ;
  assign n7604 = n7599 ^ n7359 ^ n7100 ;
  assign n7605 = n7596 ^ n7446 ^ n7103 ;
  assign n7606 = n7590 ^ n7441 ^ n7136 ;
  assign n7607 = n7588 ^ n7364 ^ n7133 ;
  assign n7608 = n7578 ^ n7367 ^ n7142 ;
  assign n7609 = n7575 ^ n7510 ^ n5964 ;
  assign n7610 = n7503 ^ n6171 ^ 1'b0 ;
  assign n7611 = n7575 ^ n7497 ^ n6630 ;
  assign n7612 = n7512 ^ n5743 ^ 1'b0 ;
  assign n7613 = n7575 ^ n7500 ^ n6401 ;
  assign n7614 = n7575 & n7612 ;
  assign n7615 = n7614 ^ n7575 ^ n7341 ;
  assign n7616 = n7575 & n7613 ;
  assign n7617 = n7542 ^ n1766 ^ 1'b0 ;
  assign n7618 = n7526 ^ n4167 ^ 1'b0 ;
  assign n7619 = n7575 & n7610 ;
  assign n7620 = n7524 ^ n4534 ^ 1'b0 ;
  assign n7621 = n7575 ^ n7521 ^ n5124 ;
  assign n7622 = n7575 & n7609 ;
  assign n7623 = n7575 ^ n7530 ^ n3464 ;
  assign n7624 = n7575 & n7611 ;
  assign n7625 = n7575 & n7617 ;
  assign n7626 = n7619 ^ n7575 ^ n7489 ;
  assign n7627 = n7575 ^ n7520 ^ n5319 ;
  assign n7628 = n7548 ^ n1118 ^ 1'b0 ;
  assign n7629 = n7575 & n7628 ;
  assign n7630 = n7540 ^ n2009 ^ 1'b0 ;
  assign n7631 = n7532 ^ n3141 ^ 1'b0 ;
  assign n7632 = n7575 & n7630 ;
  assign n7633 = n7575 & n7631 ;
  assign n7634 = n7575 & n7627 ;
  assign n7635 = n7575 & n7620 ;
  assign n7636 = n7558 ^ n399 ^ 1'b0 ;
  assign n7637 = n7575 ^ n7528 ^ n3804 ;
  assign n7638 = n7575 & n7618 ;
  assign n7639 = n7575 ^ n7549 ^ n1034 ;
  assign n7640 = n7550 ^ n941 ^ 1'b0 ;
  assign n7641 = n7575 ^ n7552 ^ n785 ;
  assign n7642 = n7575 ^ n7547 ^ n1220 ;
  assign n7643 = n7534 ^ n2839 ^ 1'b0 ;
  assign n7644 = n7575 ^ n7529 ^ n3631 ;
  assign n7645 = n7575 ^ n7535 ^ n2690 ;
  assign n7646 = n7575 & n7640 ;
  assign n7647 = n7575 & n7636 ;
  assign n7648 = n7575 & n7643 ;
  assign n7649 = n7572 & ~n7574 ;
  assign n7650 = n7622 ^ n7460 ^ n7260 ;
  assign n7651 = n7634 ^ n7502 ^ n7175 ;
  assign n7652 = n7616 ^ n7491 ^ n7252 ;
  assign n7653 = n7624 ^ n7339 ^ n7223 ;
  assign n7654 = n7629 ^ n7575 ^ n7353 ;
  assign n7655 = n7575 & n7637 ;
  assign n7656 = n7655 ^ n7499 ^ n7195 ;
  assign n7657 = n7575 & n7645 ;
  assign n7658 = n7657 ^ n7398 ^ n7181 ;
  assign n7659 = n7575 & n7642 ;
  assign n7660 = n7659 ^ n7423 ^ n7188 ;
  assign n7661 = n7575 & n7621 ;
  assign n7662 = n7661 ^ n7343 ^ n7211 ;
  assign n7663 = n7575 & n7639 ;
  assign n7664 = n7663 ^ n7426 ^ n7115 ;
  assign n7665 = n7635 ^ n7575 ^ n7518 ;
  assign n7666 = n7638 ^ n7575 ^ n7448 ;
  assign n7667 = n7575 & n7644 ;
  assign n7668 = n7633 ^ n7575 ^ n7487 ;
  assign n7669 = n7575 & n7623 ;
  assign n7670 = n7669 ^ n7506 ^ n7196 ;
  assign n7671 = n7648 ^ n7575 ^ n7463 ;
  assign n7672 = n7632 ^ n7575 ^ n7349 ;
  assign n7673 = n7625 ^ n7575 ^ n7351 ;
  assign n7674 = n7575 & n7641 ;
  assign n7675 = n7337 & ~n7574 ;
  assign n7676 = n7646 ^ n7575 ^ n7355 ;
  assign n7677 = n7674 ^ n7470 ^ n7205 ;
  assign n7678 = n7667 ^ n7392 ^ n7184 ;
  assign n7679 = n7647 ^ n7575 ^ n7362 ;
  assign n7680 = ~n7492 & n7575 ;
  assign n7681 = n7675 | n7680 ;
  assign n7682 = n7580 ^ n7464 ^ x36 ;
  assign n7683 = n7575 ^ n7496 ^ n6858 ;
  assign n7684 = n7575 & n7683 ;
  assign n7685 = n7684 ^ n7377 ^ x37 ;
  assign n7686 = n7575 ^ n7517 ^ n5527 ;
  assign n7687 = n7575 & n7686 ;
  assign n7688 = n7687 ^ n7513 ^ n7182 ;
  assign n7689 = n7575 ^ n7522 ^ n4915 ;
  assign n7690 = n7575 & n7689 ;
  assign n7691 = n7690 ^ n7382 ^ n7161 ;
  assign n7692 = n7575 ^ n7523 ^ n4728 ;
  assign n7693 = n7575 & n7692 ;
  assign n7694 = n7693 ^ n7346 ^ n7207 ;
  assign n7695 = n7575 ^ n7525 ^ n4346 ;
  assign n7696 = n7575 & n7695 ;
  assign n7697 = n7696 ^ n7385 ^ n7201 ;
  assign n7698 = n7575 ^ n7527 ^ n3986 ;
  assign n7699 = n7575 & n7698 ;
  assign n7700 = n7699 ^ n7390 ^ n7192 ;
  assign n7701 = n7575 ^ n7531 ^ n3302 ;
  assign n7702 = n7575 & n7701 ;
  assign n7703 = n7702 ^ n7474 ^ n7209 ;
  assign n7704 = n7575 ^ n7533 ^ n2995 ;
  assign n7705 = n7575 & n7704 ;
  assign n7706 = n7705 ^ n7395 ^ n7199 ;
  assign n7707 = n7575 ^ n7536 ^ n2544 ;
  assign n7708 = n7575 & n7707 ;
  assign n7709 = n7708 ^ n7402 ^ n7190 ;
  assign n7710 = n7575 ^ n7537 ^ n2404 ;
  assign n7711 = n7575 & n7710 ;
  assign n7712 = n7711 ^ n7478 ^ n7106 ;
  assign n7713 = n7575 ^ n7538 ^ n2269 ;
  assign n7714 = n7575 & n7713 ;
  assign n7715 = n7714 ^ n7405 ^ n7218 ;
  assign n7716 = n7575 ^ n7539 ^ n2139 ;
  assign n7717 = n7575 & n7716 ;
  assign n7718 = n7717 ^ n7408 ^ n7179 ;
  assign n7719 = n7575 ^ n7541 ^ n1885 ;
  assign n7720 = n7575 & n7719 ;
  assign n7721 = n7720 ^ n7411 ^ n7204 ;
  assign n7722 = n7575 ^ n7543 ^ n1652 ;
  assign n7723 = n7575 & n7722 ;
  assign n7724 = n7723 ^ n7458 ^ n7234 ;
  assign n7725 = n7575 ^ n7544 ^ n1534 ;
  assign n7726 = n7575 & n7725 ;
  assign n7727 = n7726 ^ n7414 ^ n7109 ;
  assign n7728 = n7575 ^ n7545 ^ n1416 ;
  assign n7729 = n7575 & n7728 ;
  assign n7730 = n7729 ^ n7417 ^ n7186 ;
  assign n7731 = n7575 ^ n7546 ^ n1318 ;
  assign n7732 = n7575 & n7731 ;
  assign n7733 = n7732 ^ n7420 ^ n7097 ;
  assign n7734 = n7575 ^ n7551 ^ n859 ;
  assign n7735 = n7575 & n7734 ;
  assign n7736 = n7735 ^ n7429 ^ n7219 ;
  assign n7737 = n7575 ^ n7554 ^ n640 ;
  assign n7738 = n7575 & n7737 ;
  assign n7739 = n7738 ^ n7468 ^ n7118 ;
  assign n7740 = n7681 ^ x35 ^ 1'b0 ;
  assign n7741 = x31 | x32 ;
  assign n7742 = x33 & n7575 ;
  assign n7743 = ( x33 & ~n7335 ) | ( x33 & n7741 ) | ( ~n7335 & n7741 ) ;
  assign n7744 = x33 | n7741 ;
  assign n7745 = n7742 ^ n7575 ^ x34 ;
  assign n7746 = ( n7337 & n7742 ) | ( n7337 & ~n7744 ) | ( n7742 & ~n7744 ) ;
  assign n7747 = ( ~n7337 & n7742 ) | ( ~n7337 & n7743 ) | ( n7742 & n7743 ) ;
  assign n7748 = ~n7742 & n7747 ;
  assign n7749 = n7745 | n7748 ;
  assign n7750 = ~n7746 & n7749 ;
  assign n7751 = ( ~n7089 & n7740 ) | ( ~n7089 & n7750 ) | ( n7740 & n7750 ) ;
  assign n7752 = ( ~n6858 & n7682 ) | ( ~n6858 & n7751 ) | ( n7682 & n7751 ) ;
  assign n7753 = ( ~n6630 & n7685 ) | ( ~n6630 & n7752 ) | ( n7685 & n7752 ) ;
  assign n7754 = ( ~n6401 & n7653 ) | ( ~n6401 & n7753 ) | ( n7653 & n7753 ) ;
  assign n7755 = ( ~n6171 & n7652 ) | ( ~n6171 & n7754 ) | ( n7652 & n7754 ) ;
  assign n7756 = ( ~n5964 & n7626 ) | ( ~n5964 & n7755 ) | ( n7626 & n7755 ) ;
  assign n7757 = ( ~n7498 & n7575 ) | ( ~n7498 & n7649 ) | ( n7575 & n7649 ) ;
  assign n7758 = ( ~n5743 & n7650 ) | ( ~n5743 & n7756 ) | ( n7650 & n7756 ) ;
  assign n7759 = ( ~n5527 & n7615 ) | ( ~n5527 & n7758 ) | ( n7615 & n7758 ) ;
  assign n7760 = ( ~n5319 & n7688 ) | ( ~n5319 & n7759 ) | ( n7688 & n7759 ) ;
  assign n7761 = ( ~n5124 & n7651 ) | ( ~n5124 & n7760 ) | ( n7651 & n7760 ) ;
  assign n7762 = ( ~n4915 & n7662 ) | ( ~n4915 & n7761 ) | ( n7662 & n7761 ) ;
  assign n7763 = ( ~n4728 & n7691 ) | ( ~n4728 & n7762 ) | ( n7691 & n7762 ) ;
  assign n7764 = ( ~n4534 & n7694 ) | ( ~n4534 & n7763 ) | ( n7694 & n7763 ) ;
  assign n7765 = ( ~n4346 & n7665 ) | ( ~n4346 & n7764 ) | ( n7665 & n7764 ) ;
  assign n7766 = ( ~n4167 & n7697 ) | ( ~n4167 & n7765 ) | ( n7697 & n7765 ) ;
  assign n7767 = ( ~n3986 & n7666 ) | ( ~n3986 & n7766 ) | ( n7666 & n7766 ) ;
  assign n7768 = ( ~n3804 & n7700 ) | ( ~n3804 & n7767 ) | ( n7700 & n7767 ) ;
  assign n7769 = ( n136 & n7498 ) | ( n136 & n7567 ) | ( n7498 & n7567 ) ;
  assign n7770 = n7567 & ~n7757 ;
  assign n7771 = ( ~n3631 & n7656 ) | ( ~n3631 & n7768 ) | ( n7656 & n7768 ) ;
  assign n7772 = ( ~n3464 & n7678 ) | ( ~n3464 & n7771 ) | ( n7678 & n7771 ) ;
  assign n7773 = ( n7649 & n7769 ) | ( n7649 & ~n7770 ) | ( n7769 & ~n7770 ) ;
  assign n7774 = ( ~n3302 & n7670 ) | ( ~n3302 & n7772 ) | ( n7670 & n7772 ) ;
  assign n7775 = ( ~n3141 & n7703 ) | ( ~n3141 & n7774 ) | ( n7703 & n7774 ) ;
  assign n7776 = ( ~n2995 & n7668 ) | ( ~n2995 & n7775 ) | ( n7668 & n7775 ) ;
  assign n7777 = ( ~n2839 & n7706 ) | ( ~n2839 & n7776 ) | ( n7706 & n7776 ) ;
  assign n7778 = ( ~n2690 & n7671 ) | ( ~n2690 & n7777 ) | ( n7671 & n7777 ) ;
  assign n7779 = ( ~n2544 & n7658 ) | ( ~n2544 & n7778 ) | ( n7658 & n7778 ) ;
  assign n7780 = ( ~n2404 & n7709 ) | ( ~n2404 & n7779 ) | ( n7709 & n7779 ) ;
  assign n7781 = ( ~n2269 & n7712 ) | ( ~n2269 & n7780 ) | ( n7712 & n7780 ) ;
  assign n7782 = ( ~n2139 & n7715 ) | ( ~n2139 & n7781 ) | ( n7715 & n7781 ) ;
  assign n7783 = ( ~n2009 & n7718 ) | ( ~n2009 & n7782 ) | ( n7718 & n7782 ) ;
  assign n7784 = ( ~n1885 & n7672 ) | ( ~n1885 & n7783 ) | ( n7672 & n7783 ) ;
  assign n7785 = ( ~n1766 & n7721 ) | ( ~n1766 & n7784 ) | ( n7721 & n7784 ) ;
  assign n7786 = ( ~n1652 & n7673 ) | ( ~n1652 & n7785 ) | ( n7673 & n7785 ) ;
  assign n7787 = ( ~n1534 & n7724 ) | ( ~n1534 & n7786 ) | ( n7724 & n7786 ) ;
  assign n7788 = ( ~n1416 & n7727 ) | ( ~n1416 & n7787 ) | ( n7727 & n7787 ) ;
  assign n7789 = ( ~n1318 & n7730 ) | ( ~n1318 & n7788 ) | ( n7730 & n7788 ) ;
  assign n7790 = ( ~n1220 & n7733 ) | ( ~n1220 & n7789 ) | ( n7733 & n7789 ) ;
  assign n7791 = ( ~n1118 & n7660 ) | ( ~n1118 & n7790 ) | ( n7660 & n7790 ) ;
  assign n7792 = n7567 ^ n7498 ^ 1'b0 ;
  assign n7793 = ( n7498 & ~n7567 ) | ( n7498 & n7575 ) | ( ~n7567 & n7575 ) ;
  assign n7794 = n7746 | n7748 ;
  assign n7795 = n7791 ^ n1034 ^ 1'b0 ;
  assign n7796 = ( n7567 & ~n7792 ) | ( n7567 & n7793 ) | ( ~n7792 & n7793 ) ;
  assign n7797 = ( n7569 & ~n7773 ) | ( n7569 & n7796 ) | ( ~n7773 & n7796 ) ;
  assign n7798 = ( x11 & x116 ) | ( x11 & ~n7649 ) | ( x116 & ~n7649 ) ;
  assign n7799 = ( ~n1034 & n7654 ) | ( ~n1034 & n7791 ) | ( n7654 & n7791 ) ;
  assign n7800 = ( x127 & ~n7649 ) | ( x127 & n7798 ) | ( ~n7649 & n7798 ) ;
  assign n7801 = ( ~n941 & n7664 ) | ( ~n941 & n7799 ) | ( n7664 & n7799 ) ;
  assign n7802 = ( ~n859 & n7676 ) | ( ~n859 & n7801 ) | ( n7676 & n7801 ) ;
  assign n7803 = ( ~n785 & n7736 ) | ( ~n785 & n7802 ) | ( n7736 & n7802 ) ;
  assign n7804 = ( ~n716 & n7677 ) | ( ~n716 & n7803 ) | ( n7677 & n7803 ) ;
  assign n7805 = ( ~n640 & n7602 ) | ( ~n640 & n7804 ) | ( n7602 & n7804 ) ;
  assign n7806 = ( ~n572 & n7739 ) | ( ~n572 & n7805 ) | ( n7739 & n7805 ) ;
  assign n7807 = ( ~n514 & n7600 ) | ( ~n514 & n7806 ) | ( n7600 & n7806 ) ;
  assign n7808 = ( ~n458 & n7583 ) | ( ~n458 & n7807 ) | ( n7583 & n7807 ) ;
  assign n7809 = ( ~n399 & n7604 ) | ( ~n399 & n7808 ) | ( n7604 & n7808 ) ;
  assign n7810 = ( ~n345 & n7679 ) | ( ~n345 & n7809 ) | ( n7679 & n7809 ) ;
  assign n7811 = ( ~n302 & n7601 ) | ( ~n302 & n7810 ) | ( n7601 & n7810 ) ;
  assign n7812 = ( ~n261 & n7607 ) | ( ~n261 & n7811 ) | ( n7607 & n7811 ) ;
  assign n7813 = ( ~n217 & n7606 ) | ( ~n217 & n7812 ) | ( n7606 & n7812 ) ;
  assign n7814 = ( ~n179 & n7603 ) | ( ~n179 & n7813 ) | ( n7603 & n7813 ) ;
  assign n7815 = ( ~n144 & n7608 ) | ( ~n144 & n7814 ) | ( n7608 & n7814 ) ;
  assign n7816 = ( ~n134 & n7584 ) | ( ~n134 & n7815 ) | ( n7584 & n7815 ) ;
  assign n7817 = ( ~n136 & n7605 ) | ( ~n136 & n7816 ) | ( n7605 & n7816 ) ;
  assign n7818 = n7796 | n7817 ;
  assign n7819 = ~n136 & n7818 ;
  assign n7820 = n7605 & n7816 ;
  assign n7821 = ( n7773 & n7800 ) | ( n7773 & ~n7820 ) | ( n7800 & ~n7820 ) ;
  assign n7822 = ~n7773 & n7821 ;
  assign n7823 = n7819 | n7820 ;
  assign n7824 = n7773 | n7823 ;
  assign n7825 = n7794 & n7824 ;
  assign n7826 = n7824 ^ n7802 ^ n785 ;
  assign n7827 = n7824 ^ n7786 ^ n1534 ;
  assign n7828 = n7795 & n7824 ;
  assign n7829 = n7824 ^ n7813 ^ n179 ;
  assign n7830 = n7824 ^ n7810 ^ n302 ;
  assign n7831 = n7824 & n7830 ;
  assign n7832 = n7824 ^ n7784 ^ n1766 ;
  assign n7833 = n7824 & n7832 ;
  assign n7834 = n7825 ^ n7824 ^ n7745 ;
  assign n7835 = n7824 ^ n7803 ^ n716 ;
  assign n7836 = n7824 ^ n7811 ^ n261 ;
  assign n7837 = ~n7741 & n7824 ;
  assign n7838 = n7824 & n7835 ;
  assign n7839 = n7824 & n7836 ;
  assign n7840 = n7838 ^ n7674 ^ n7515 ;
  assign n7841 = n7824 ^ n7782 ^ n2009 ;
  assign n7842 = n7824 ^ n7806 ^ n514 ;
  assign n7843 = n7824 ^ n7808 ^ n399 ;
  assign n7844 = n7824 ^ n7780 ^ n2269 ;
  assign n7845 = n7824 & n7841 ;
  assign n7846 = n7824 & n7844 ;
  assign n7847 = n7845 ^ n7717 ^ n7409 ;
  assign n7848 = n7824 & n7843 ;
  assign n7849 = n7824 ^ n7774 ^ n3141 ;
  assign n7850 = n7824 & n7842 ;
  assign n7851 = n7846 ^ n7711 ^ n7483 ;
  assign n7852 = n7824 & n7827 ;
  assign n7853 = n7824 ^ n7771 ^ n3464 ;
  assign n7854 = n7852 ^ n7723 ^ n7465 ;
  assign n7855 = n7824 & n7853 ;
  assign n7856 = n7824 ^ n7812 ^ n217 ;
  assign n7857 = n7823 & ~n7837 ;
  assign n7858 = n7824 & n7856 ;
  assign n7859 = ( n7797 & n7837 ) | ( n7797 & ~n7857 ) | ( n7837 & ~n7857 ) ;
  assign n7860 = n7850 ^ n7597 ^ n7436 ;
  assign n7861 = n7824 & n7826 ;
  assign n7862 = n7824 & n7849 ;
  assign n7863 = n7824 ^ n7772 ^ n3302 ;
  assign n7864 = n7862 ^ n7702 ^ n7475 ;
  assign n7865 = n7861 ^ n7735 ^ n7430 ;
  assign n7866 = n7828 ^ n7824 ^ n7654 ;
  assign n7867 = n7824 ^ n7763 ^ n4534 ;
  assign n7868 = n7824 & n7829 ;
  assign n7869 = n7824 & n7867 ;
  assign n7870 = n7855 ^ n7667 ^ n7393 ;
  assign n7871 = n7869 ^ n7693 ^ n7347 ;
  assign n7872 = n7824 & n7863 ;
  assign n7873 = n7872 ^ n7669 ^ n7511 ;
  assign n7874 = n7833 ^ n7720 ^ n7412 ;
  assign n7875 = n7858 ^ n7590 ^ n7442 ;
  assign n7876 = n7848 ^ n7599 ^ n7360 ;
  assign n7877 = n7868 ^ n7589 ^ n7445 ;
  assign n7878 = n7831 ^ n7592 ^ n7439 ;
  assign n7879 = n7839 ^ n7588 ^ n7365 ;
  assign n7880 = n7824 ^ n7751 ^ n6858 ;
  assign n7881 = n7824 & n7880 ;
  assign n7882 = n7881 ^ n7580 ^ n7466 ;
  assign n7883 = n7824 ^ n7754 ^ n6171 ;
  assign n7884 = n7824 ^ n7756 ^ n5743 ;
  assign n7885 = n7824 & n7884 ;
  assign n7886 = n7885 ^ n7622 ^ n7462 ;
  assign n7887 = n7824 ^ n7759 ^ n5319 ;
  assign n7888 = n7824 & n7887 ;
  assign n7889 = n7888 ^ n7687 ^ n7514 ;
  assign n7890 = n7824 ^ n7760 ^ n5124 ;
  assign n7891 = n7824 & n7890 ;
  assign n7892 = n7891 ^ n7634 ^ n7504 ;
  assign n7893 = n7824 ^ n7761 ^ n4915 ;
  assign n7894 = n7824 & n7893 ;
  assign n7895 = n7894 ^ n7661 ^ n7344 ;
  assign n7896 = n7824 ^ n7762 ^ n4728 ;
  assign n7897 = n7824 & n7883 ;
  assign n7898 = n7897 ^ n7616 ^ n7495 ;
  assign n7899 = n7824 & n7896 ;
  assign n7900 = n7899 ^ n7690 ^ n7383 ;
  assign n7901 = n7824 ^ n7767 ^ n3804 ;
  assign n7902 = n7824 & n7901 ;
  assign n7903 = n7902 ^ n7699 ^ n7399 ;
  assign n7904 = n7824 ^ n7768 ^ n3631 ;
  assign n7905 = n7824 & n7904 ;
  assign n7906 = n7905 ^ n7655 ^ n7501 ;
  assign n7907 = n7824 ^ n7778 ^ n2544 ;
  assign n7908 = n7824 & n7907 ;
  assign n7909 = n7908 ^ n7657 ^ n7400 ;
  assign n7910 = n7824 ^ n7781 ^ n2139 ;
  assign n7911 = n7824 & n7910 ;
  assign n7912 = n7911 ^ n7714 ^ n7406 ;
  assign n7913 = n7824 ^ n7787 ^ n1416 ;
  assign n7914 = n7824 & n7913 ;
  assign n7915 = n7914 ^ n7726 ^ n7415 ;
  assign n7916 = n7824 ^ n7788 ^ n1318 ;
  assign n7917 = n7824 & n7916 ;
  assign n7918 = n7917 ^ n7729 ^ n7418 ;
  assign n7919 = n7824 ^ n7789 ^ n1220 ;
  assign n7920 = n7824 & n7919 ;
  assign n7921 = n7920 ^ n7732 ^ n7421 ;
  assign n7922 = n7824 ^ n7790 ^ n1118 ;
  assign n7923 = n7824 & n7922 ;
  assign n7924 = n7923 ^ n7659 ^ n7424 ;
  assign n7925 = n7824 ^ n7799 ^ n941 ;
  assign n7926 = n7824 & n7925 ;
  assign n7927 = n7926 ^ n7663 ^ n7427 ;
  assign n7928 = n7801 ^ n859 ^ 1'b0 ;
  assign n7929 = n7824 & n7928 ;
  assign n7930 = n7929 ^ n7824 ^ n7676 ;
  assign n7931 = n7824 ^ n7804 ^ n640 ;
  assign n7932 = n7824 & n7931 ;
  assign n7933 = n7932 ^ n7598 ^ n7433 ;
  assign n7934 = n7824 ^ n7805 ^ n572 ;
  assign n7935 = n7824 & n7934 ;
  assign n7936 = n7935 ^ n7738 ^ n7481 ;
  assign n7937 = n7807 ^ n458 ^ 1'b0 ;
  assign n7938 = n7824 & n7937 ;
  assign n7939 = n7938 ^ n7824 ^ n7583 ;
  assign n7940 = n7824 ^ n7814 ^ n144 ;
  assign n7941 = n7824 & n7940 ;
  assign n7942 = n7941 ^ n7578 ^ n7368 ;
  assign n7943 = n7824 ^ n7750 ^ n7089 ;
  assign n7944 = n7824 & n7943 ;
  assign n7945 = n7944 ^ n7681 ^ x35 ;
  assign n7946 = n7824 ^ n7752 ^ n6630 ;
  assign n7947 = n7824 & n7946 ;
  assign n7948 = n7947 ^ n7684 ^ n7477 ;
  assign n7949 = n7824 ^ n7753 ^ n6401 ;
  assign n7950 = n7824 & n7949 ;
  assign n7951 = n7950 ^ n7624 ^ n7455 ;
  assign n7952 = n7755 ^ n5964 ^ 1'b0 ;
  assign n7953 = n7824 & n7952 ;
  assign n7954 = n7953 ^ n7824 ^ n7626 ;
  assign n7955 = n7758 ^ n5527 ^ 1'b0 ;
  assign n7956 = n7824 & n7955 ;
  assign n7957 = n7956 ^ n7824 ^ n7615 ;
  assign n7958 = n7764 ^ n4346 ^ 1'b0 ;
  assign n7959 = n7824 & n7958 ;
  assign n7960 = n7824 ^ n7765 ^ n4167 ;
  assign n7961 = n7824 & n7960 ;
  assign n7962 = n7961 ^ n7696 ^ n7386 ;
  assign n7963 = n7766 ^ n3986 ^ 1'b0 ;
  assign n7964 = n7824 & n7963 ;
  assign n7965 = n7964 ^ n7824 ^ n7666 ;
  assign n7966 = n7775 ^ n2995 ^ 1'b0 ;
  assign n7967 = n7824 & n7966 ;
  assign n7968 = n7967 ^ n7824 ^ n7668 ;
  assign n7969 = n7824 ^ n7776 ^ n2839 ;
  assign n7970 = n7824 & n7969 ;
  assign n7971 = n7970 ^ n7705 ^ n7396 ;
  assign n7972 = n7777 ^ n2690 ^ 1'b0 ;
  assign n7973 = n7824 & n7972 ;
  assign n7974 = n7973 ^ n7824 ^ n7671 ;
  assign n7975 = n7824 ^ n7779 ^ n2404 ;
  assign n7976 = n7824 & n7975 ;
  assign n7977 = n7976 ^ n7708 ^ n7403 ;
  assign n7978 = n7783 ^ n1885 ^ 1'b0 ;
  assign n7979 = n7824 & n7978 ;
  assign n7980 = n7979 ^ n7824 ^ n7672 ;
  assign n7981 = n7785 ^ n1652 ^ 1'b0 ;
  assign n7982 = n7824 & n7981 ;
  assign n7983 = n7982 ^ n7824 ^ n7673 ;
  assign n7984 = n7809 ^ n345 ^ 1'b0 ;
  assign n7985 = n7824 & n7984 ;
  assign n7986 = n7985 ^ n7824 ^ n7679 ;
  assign n7987 = n7815 ^ n134 ^ 1'b0 ;
  assign n7988 = n7824 & n7987 ;
  assign n7989 = n7988 ^ n7824 ^ n7584 ;
  assign n7990 = ( n7605 & ~n7816 ) | ( n7605 & n7824 ) | ( ~n7816 & n7824 ) ;
  assign n7991 = n7605 & ~n7816 ;
  assign n7992 = ( n7989 & n7990 ) | ( n7989 & ~n7991 ) | ( n7990 & ~n7991 ) ;
  assign n7993 = ( n7816 & n7817 ) | ( n7816 & n7824 ) | ( n7817 & n7824 ) ;
  assign n7994 = n7605 & ~n7993 ;
  assign n7995 = n7994 ^ n7993 ^ n7817 ;
  assign n7996 = n7959 ^ n7824 ^ n7665 ;
  assign n7997 = n7859 ^ x33 ^ 1'b0 ;
  assign n7998 = x11 | x22 ;
  assign n7999 = ( x31 & n7575 ) | ( x31 & ~n7998 ) | ( n7575 & ~n7998 ) ;
  assign n8000 = ( ~x31 & n7575 ) | ( ~x31 & n7824 ) | ( n7575 & n7824 ) ;
  assign n8001 = n7999 & n8000 ;
  assign n8002 = x31 & n7824 ;
  assign n8003 = n8002 ^ n7824 ^ x32 ;
  assign n8004 = ( x31 & ~n7571 ) | ( x31 & n7998 ) | ( ~n7571 & n7998 ) ;
  assign n8005 = ( ~n7575 & n8002 ) | ( ~n7575 & n8004 ) | ( n8002 & n8004 ) ;
  assign n8006 = ~n8002 & n8005 ;
  assign n8007 = n8003 | n8006 ;
  assign n8008 = ~n8001 & n8007 ;
  assign n8009 = ( ~n7337 & n7997 ) | ( ~n7337 & n8008 ) | ( n7997 & n8008 ) ;
  assign n8010 = ( ~n7089 & n7834 ) | ( ~n7089 & n8009 ) | ( n7834 & n8009 ) ;
  assign n8011 = ( ~n6858 & n7945 ) | ( ~n6858 & n8010 ) | ( n7945 & n8010 ) ;
  assign n8012 = ( ~n6630 & n7882 ) | ( ~n6630 & n8011 ) | ( n7882 & n8011 ) ;
  assign n8013 = ( ~n6401 & n7948 ) | ( ~n6401 & n8012 ) | ( n7948 & n8012 ) ;
  assign n8014 = ( ~n6171 & n7951 ) | ( ~n6171 & n8013 ) | ( n7951 & n8013 ) ;
  assign n8015 = ( ~n5964 & n7898 ) | ( ~n5964 & n8014 ) | ( n7898 & n8014 ) ;
  assign n8016 = ( ~n5743 & n7954 ) | ( ~n5743 & n8015 ) | ( n7954 & n8015 ) ;
  assign n8017 = ( ~n5527 & n7886 ) | ( ~n5527 & n8016 ) | ( n7886 & n8016 ) ;
  assign n8018 = ( ~n5319 & n7957 ) | ( ~n5319 & n8017 ) | ( n7957 & n8017 ) ;
  assign n8019 = ( ~n5124 & n7889 ) | ( ~n5124 & n8018 ) | ( n7889 & n8018 ) ;
  assign n8020 = ( ~n4915 & n7892 ) | ( ~n4915 & n8019 ) | ( n7892 & n8019 ) ;
  assign n8021 = ( ~n4728 & n7895 ) | ( ~n4728 & n8020 ) | ( n7895 & n8020 ) ;
  assign n8022 = ( ~n4534 & n7900 ) | ( ~n4534 & n8021 ) | ( n7900 & n8021 ) ;
  assign n8023 = ( ~n4346 & n7871 ) | ( ~n4346 & n8022 ) | ( n7871 & n8022 ) ;
  assign n8024 = ( ~n4167 & n7996 ) | ( ~n4167 & n8023 ) | ( n7996 & n8023 ) ;
  assign n8025 = ( ~n3986 & n7962 ) | ( ~n3986 & n8024 ) | ( n7962 & n8024 ) ;
  assign n8026 = ( ~n3804 & n7965 ) | ( ~n3804 & n8025 ) | ( n7965 & n8025 ) ;
  assign n8027 = ( ~n3631 & n7903 ) | ( ~n3631 & n8026 ) | ( n7903 & n8026 ) ;
  assign n8028 = ( ~n3464 & n7906 ) | ( ~n3464 & n8027 ) | ( n7906 & n8027 ) ;
  assign n8029 = ( ~n3302 & n7870 ) | ( ~n3302 & n8028 ) | ( n7870 & n8028 ) ;
  assign n8030 = ( ~n3141 & n7873 ) | ( ~n3141 & n8029 ) | ( n7873 & n8029 ) ;
  assign n8031 = ( ~n2995 & n7864 ) | ( ~n2995 & n8030 ) | ( n7864 & n8030 ) ;
  assign n8032 = ( ~n2839 & n7968 ) | ( ~n2839 & n8031 ) | ( n7968 & n8031 ) ;
  assign n8033 = ( ~n2690 & n7971 ) | ( ~n2690 & n8032 ) | ( n7971 & n8032 ) ;
  assign n8034 = ( ~n2544 & n7974 ) | ( ~n2544 & n8033 ) | ( n7974 & n8033 ) ;
  assign n8035 = ( ~n2404 & n7909 ) | ( ~n2404 & n8034 ) | ( n7909 & n8034 ) ;
  assign n8036 = ( ~n2269 & n7977 ) | ( ~n2269 & n8035 ) | ( n7977 & n8035 ) ;
  assign n8037 = ( ~n2139 & n7851 ) | ( ~n2139 & n8036 ) | ( n7851 & n8036 ) ;
  assign n8038 = ( ~n2009 & n7912 ) | ( ~n2009 & n8037 ) | ( n7912 & n8037 ) ;
  assign n8039 = ( ~n1885 & n7847 ) | ( ~n1885 & n8038 ) | ( n7847 & n8038 ) ;
  assign n8040 = ( ~n1766 & n7980 ) | ( ~n1766 & n8039 ) | ( n7980 & n8039 ) ;
  assign n8041 = ( ~n1652 & n7874 ) | ( ~n1652 & n8040 ) | ( n7874 & n8040 ) ;
  assign n8042 = ( ~n1534 & n7983 ) | ( ~n1534 & n8041 ) | ( n7983 & n8041 ) ;
  assign n8043 = ( ~n1416 & n7854 ) | ( ~n1416 & n8042 ) | ( n7854 & n8042 ) ;
  assign n8044 = ( ~n1318 & n7915 ) | ( ~n1318 & n8043 ) | ( n7915 & n8043 ) ;
  assign n8045 = ( ~n1220 & n7918 ) | ( ~n1220 & n8044 ) | ( n7918 & n8044 ) ;
  assign n8046 = ( ~n1118 & n7921 ) | ( ~n1118 & n8045 ) | ( n7921 & n8045 ) ;
  assign n8047 = ( ~n1034 & n7924 ) | ( ~n1034 & n8046 ) | ( n7924 & n8046 ) ;
  assign n8048 = ( ~n941 & n7866 ) | ( ~n941 & n8047 ) | ( n7866 & n8047 ) ;
  assign n8049 = ( ~n859 & n7927 ) | ( ~n859 & n8048 ) | ( n7927 & n8048 ) ;
  assign n8050 = n8001 | n8006 ;
  assign n8051 = ( ~n785 & n7930 ) | ( ~n785 & n8049 ) | ( n7930 & n8049 ) ;
  assign n8052 = ( ~n716 & n7865 ) | ( ~n716 & n8051 ) | ( n7865 & n8051 ) ;
  assign n8053 = ( ~n640 & n7840 ) | ( ~n640 & n8052 ) | ( n7840 & n8052 ) ;
  assign n8054 = ( ~n572 & n7933 ) | ( ~n572 & n8053 ) | ( n7933 & n8053 ) ;
  assign n8055 = ( ~n514 & n7936 ) | ( ~n514 & n8054 ) | ( n7936 & n8054 ) ;
  assign n8056 = ( ~n458 & n7860 ) | ( ~n458 & n8055 ) | ( n7860 & n8055 ) ;
  assign n8057 = ( ~n399 & n7939 ) | ( ~n399 & n8056 ) | ( n7939 & n8056 ) ;
  assign n8058 = ( ~n345 & n7876 ) | ( ~n345 & n8057 ) | ( n7876 & n8057 ) ;
  assign n8059 = ( ~n302 & n7986 ) | ( ~n302 & n8058 ) | ( n7986 & n8058 ) ;
  assign n8060 = ( ~n261 & n7878 ) | ( ~n261 & n8059 ) | ( n7878 & n8059 ) ;
  assign n8061 = ( ~n217 & n7879 ) | ( ~n217 & n8060 ) | ( n7879 & n8060 ) ;
  assign n8062 = ( ~n179 & n7875 ) | ( ~n179 & n8061 ) | ( n7875 & n8061 ) ;
  assign n8063 = ( ~n144 & n7877 ) | ( ~n144 & n8062 ) | ( n7877 & n8062 ) ;
  assign n8064 = ( ~n134 & n7942 ) | ( ~n134 & n8063 ) | ( n7942 & n8063 ) ;
  assign n8065 = ( ~x30 & n7992 ) | ( ~x30 & n8064 ) | ( n7992 & n8064 ) ;
  assign n8066 = ~n136 & n8065 ;
  assign n8067 = n7989 & n8064 ;
  assign n8068 = n7995 | n8067 ;
  assign n8069 = n8066 | n8068 ;
  assign n8070 = n8063 ^ n134 ^ 1'b0 ;
  assign n8071 = n8069 & ~n8070 ;
  assign n8072 = n8071 ^ n7941 ^ n7608 ;
  assign n8073 = n8069 ^ n8010 ^ n6858 ;
  assign n8074 = n8069 & n8073 ;
  assign n8075 = n8074 ^ n7944 ^ n7740 ;
  assign n8076 = n8050 & n8069 ;
  assign n8077 = n8076 ^ n8069 ^ n8003 ;
  assign n8078 = n8069 ^ n8011 ^ n6630 ;
  assign n8079 = n8069 & n8078 ;
  assign n8080 = n8079 ^ n7881 ^ n7682 ;
  assign n8081 = n8069 ^ n8012 ^ n6401 ;
  assign n8082 = n8069 & n8081 ;
  assign n8083 = n8082 ^ n7947 ^ n7685 ;
  assign n8084 = n8069 ^ n8016 ^ n5527 ;
  assign n8085 = n8069 & n8084 ;
  assign n8086 = n8085 ^ n7885 ^ n7650 ;
  assign n8087 = n8069 ^ n8020 ^ n4728 ;
  assign n8088 = n8069 & n8087 ;
  assign n8089 = n8088 ^ n7894 ^ n7662 ;
  assign n8090 = n8069 ^ n8021 ^ n4534 ;
  assign n8091 = n8069 & n8090 ;
  assign n8092 = n8091 ^ n7899 ^ n7691 ;
  assign n8093 = n8069 ^ n8026 ^ n3631 ;
  assign n8094 = n8069 & n8093 ;
  assign n8095 = n8094 ^ n7902 ^ n7700 ;
  assign n8096 = n8069 ^ n8027 ^ n3464 ;
  assign n8097 = n8069 & n8096 ;
  assign n8098 = n8097 ^ n7905 ^ n7656 ;
  assign n8099 = n8069 ^ n8028 ^ n3302 ;
  assign n8100 = n8069 & n8099 ;
  assign n8101 = n8100 ^ n7855 ^ n7678 ;
  assign n8102 = n8069 ^ n8029 ^ n3141 ;
  assign n8103 = n8069 & n8102 ;
  assign n8104 = n8103 ^ n7872 ^ n7670 ;
  assign n8105 = n8069 ^ n8030 ^ n2995 ;
  assign n8106 = n8069 & n8105 ;
  assign n8107 = n8106 ^ n7862 ^ n7703 ;
  assign n8108 = n8069 ^ n8038 ^ n1885 ;
  assign n8109 = n8069 & n8108 ;
  assign n8110 = n8109 ^ n7845 ^ n7718 ;
  assign n8111 = n8069 ^ n8040 ^ n1652 ;
  assign n8112 = n8069 & n8111 ;
  assign n8113 = n8112 ^ n7833 ^ n7721 ;
  assign n8114 = n8069 ^ n8057 ^ n345 ;
  assign n8115 = n8069 & n8114 ;
  assign n8116 = n8115 ^ n7848 ^ n7604 ;
  assign n8117 = n8069 ^ n8062 ^ n144 ;
  assign n8118 = n8069 & n8117 ;
  assign n8119 = n8118 ^ n7868 ^ n7603 ;
  assign n8120 = n8009 ^ n7089 ^ 1'b0 ;
  assign n8121 = n8069 & n8120 ;
  assign n8122 = n8121 ^ n8069 ^ n7834 ;
  assign n8123 = n8017 ^ n5319 ^ 1'b0 ;
  assign n8124 = n8069 & n8123 ;
  assign n8125 = n8124 ^ n8069 ^ n7957 ;
  assign n8126 = n8069 ^ n8022 ^ n4346 ;
  assign n8127 = n8069 & n8126 ;
  assign n8128 = n8127 ^ n7869 ^ n7694 ;
  assign n8129 = n8023 ^ n4167 ^ 1'b0 ;
  assign n8130 = n8069 & n8129 ;
  assign n8131 = n8130 ^ n8069 ^ n7996 ;
  assign n8132 = n8025 ^ n3804 ^ 1'b0 ;
  assign n8133 = n8069 & n8132 ;
  assign n8134 = n8133 ^ n8069 ^ n7965 ;
  assign n8135 = n8031 ^ n2839 ^ 1'b0 ;
  assign n8136 = n8069 & n8135 ;
  assign n8137 = n8136 ^ n8069 ^ n7968 ;
  assign n8138 = n8033 ^ n2544 ^ 1'b0 ;
  assign n8139 = n8069 & n8138 ;
  assign n8140 = n8139 ^ n8069 ^ n7974 ;
  assign n8141 = n8039 ^ n1766 ^ 1'b0 ;
  assign n8142 = n8069 & n8141 ;
  assign n8143 = n8142 ^ n8069 ^ n7980 ;
  assign n8144 = n8041 ^ n1534 ^ 1'b0 ;
  assign n8145 = n8069 & n8144 ;
  assign n8146 = n8145 ^ n8069 ^ n7983 ;
  assign n8147 = n8069 ^ n8044 ^ n1220 ;
  assign n8148 = n8069 & n8147 ;
  assign n8149 = n8148 ^ n7917 ^ n7730 ;
  assign n8150 = n8069 ^ n8045 ^ n1118 ;
  assign n8151 = n8069 & n8150 ;
  assign n8152 = n8151 ^ n7920 ^ n7733 ;
  assign n8153 = n8047 ^ n941 ^ 1'b0 ;
  assign n8154 = n8069 & n8153 ;
  assign n8155 = n8154 ^ n8069 ^ n7866 ;
  assign n8156 = n8069 ^ n8048 ^ n859 ;
  assign n8157 = n8069 & n8156 ;
  assign n8158 = n8157 ^ n7926 ^ n7664 ;
  assign n8159 = n8049 ^ n785 ^ 1'b0 ;
  assign n8160 = n8069 & n8159 ;
  assign n8161 = n8160 ^ n8069 ^ n7930 ;
  assign n8162 = n8069 ^ n8053 ^ n572 ;
  assign n8163 = n8069 & n8162 ;
  assign n8164 = n8163 ^ n7932 ^ n7602 ;
  assign n8165 = n8069 ^ n8054 ^ n514 ;
  assign n8166 = n8069 & n8165 ;
  assign n8167 = n8166 ^ n7935 ^ n7739 ;
  assign n8168 = n8056 ^ n399 ^ 1'b0 ;
  assign n8169 = n8069 & n8168 ;
  assign n8170 = n8169 ^ n8069 ^ n7939 ;
  assign n8171 = n8069 ^ n8059 ^ n261 ;
  assign n8172 = n8069 & n8171 ;
  assign n8173 = n8172 ^ n7831 ^ n7601 ;
  assign n8174 = n8069 ^ n8061 ^ n179 ;
  assign n8175 = n8069 & n8174 ;
  assign n8176 = n8175 ^ n7858 ^ n7606 ;
  assign n8177 = n8069 ^ n8060 ^ n217 ;
  assign n8178 = n8069 ^ n8032 ^ n2690 ;
  assign n8179 = n8069 ^ n8035 ^ n2269 ;
  assign n8180 = n8069 ^ n8019 ^ n4915 ;
  assign n8181 = n8069 ^ n8037 ^ n2009 ;
  assign n8182 = n8069 ^ n8024 ^ n3986 ;
  assign n8183 = n8069 ^ n8036 ^ n2139 ;
  assign n8184 = n8069 ^ n8042 ^ n1416 ;
  assign n8185 = n8069 ^ n8046 ^ n1034 ;
  assign n8186 = n8069 ^ n8043 ^ n1318 ;
  assign n8187 = n8069 ^ n8052 ^ n640 ;
  assign n8188 = n8069 ^ n8055 ^ n458 ;
  assign n8189 = n8069 ^ n8051 ^ n716 ;
  assign n8190 = n8069 ^ n8018 ^ n5124 ;
  assign n8191 = n8069 ^ n8034 ^ n2404 ;
  assign n8192 = n8069 & n8180 ;
  assign n8193 = n8192 ^ n7891 ^ n7651 ;
  assign n8194 = n8069 & n8185 ;
  assign n8195 = n8194 ^ n7923 ^ n7660 ;
  assign n8196 = n8069 & n8191 ;
  assign n8197 = n8196 ^ n7908 ^ n7658 ;
  assign n8198 = n8069 & n8189 ;
  assign n8199 = n8198 ^ n7861 ^ n7736 ;
  assign n8200 = n8069 & n8187 ;
  assign n8201 = n8200 ^ n7838 ^ n7677 ;
  assign n8202 = n8069 & n8190 ;
  assign n8203 = n8202 ^ n7888 ^ n7688 ;
  assign n8204 = n8069 & n8182 ;
  assign n8205 = n8069 & n8188 ;
  assign n8206 = n8069 & n8179 ;
  assign n8207 = n8204 ^ n7961 ^ n7697 ;
  assign n8208 = n8069 & n8178 ;
  assign n8209 = n8069 & n8177 ;
  assign n8210 = n8209 ^ n7839 ^ n7607 ;
  assign n8211 = n8069 & n8181 ;
  assign n8212 = n8211 ^ n7911 ^ n7715 ;
  assign n8213 = n8069 & n8183 ;
  assign n8214 = n8213 ^ n7846 ^ n7712 ;
  assign n8215 = ( x11 & n7819 ) | ( x11 & n8069 ) | ( n7819 & n8069 ) ;
  assign n8216 = ( ~n7819 & n7822 ) | ( ~n7819 & n8215 ) | ( n7822 & n8215 ) ;
  assign n8217 = ~n8215 & n8216 ;
  assign n8218 = n8069 & n8184 ;
  assign n8219 = n8069 & n8186 ;
  assign n8220 = n8208 ^ n7970 ^ n7706 ;
  assign n8221 = n8218 ^ n7852 ^ n7724 ;
  assign n8222 = n8219 ^ n7914 ^ n7727 ;
  assign n8223 = n8206 ^ n7976 ^ n7709 ;
  assign n8224 = n8205 ^ n7850 ^ n7600 ;
  assign n8225 = n8058 ^ n302 ^ 1'b0 ;
  assign n8226 = n8069 & n8225 ;
  assign n8227 = n8069 ^ n8008 ^ n7337 ;
  assign n8228 = x116 | x127 ;
  assign n8229 = n8226 ^ n8069 ^ n7986 ;
  assign n8230 = ( x11 & n7824 ) | ( x11 & ~n8228 ) | ( n7824 & ~n8228 ) ;
  assign n8231 = n8015 ^ n5743 ^ 1'b0 ;
  assign n8232 = n8069 & n8231 ;
  assign n8233 = n8232 ^ n8069 ^ n7954 ;
  assign n8234 = ( ~x11 & n7824 ) | ( ~x11 & n8069 ) | ( n7824 & n8069 ) ;
  assign n8235 = n8230 & n8234 ;
  assign n8236 = n8069 & n8227 ;
  assign n8237 = n8236 ^ n7859 ^ x33 ;
  assign n8238 = ~n7998 & n8069 ;
  assign n8239 = ( n8064 & n8067 ) | ( n8064 & ~n8069 ) | ( n8067 & ~n8069 ) ;
  assign n8240 = ( n7824 & ~n8066 ) | ( n7824 & n8067 ) | ( ~n8066 & n8067 ) ;
  assign n8241 = n8068 & ~n8238 ;
  assign n8242 = ( n8238 & n8240 ) | ( n8238 & ~n8241 ) | ( n8240 & ~n8241 ) ;
  assign n8243 = ( n136 & ~n7989 ) | ( n136 & n8064 ) | ( ~n7989 & n8064 ) ;
  assign n8244 = ( n136 & n7989 ) | ( n136 & n8064 ) | ( n7989 & n8064 ) ;
  assign n8245 = ~n8239 & n8244 ;
  assign n8246 = n6171 & n8013 ;
  assign n8247 = ( ~n7989 & n8064 ) | ( ~n7989 & n8069 ) | ( n8064 & n8069 ) ;
  assign n8248 = ( ~n6171 & n8069 ) | ( ~n6171 & n8246 ) | ( n8069 & n8246 ) ;
  assign n8249 = ( n8072 & ~n8243 ) | ( n8072 & n8247 ) | ( ~n8243 & n8247 ) ;
  assign n8250 = n5964 & n8014 ;
  assign n8251 = ( ~n8013 & n8246 ) | ( ~n8013 & n8248 ) | ( n8246 & n8248 ) ;
  assign n8252 = ~x11 & n8069 ;
  assign n8253 = n8251 ^ n7950 ^ n7653 ;
  assign n8254 = n8242 ^ x31 ^ 1'b0 ;
  assign n8255 = ( ~n5964 & n8069 ) | ( ~n5964 & n8250 ) | ( n8069 & n8250 ) ;
  assign n8256 = ( ~n8014 & n8250 ) | ( ~n8014 & n8255 ) | ( n8250 & n8255 ) ;
  assign n8257 = n8252 ^ x22 ^ 1'b0 ;
  assign n8258 = n8256 ^ n7897 ^ n7652 ;
  assign n8259 = n8217 | n8257 ;
  assign n8260 = ~n8235 & n8259 ;
  assign n8261 = ( ~n7575 & n8254 ) | ( ~n7575 & n8260 ) | ( n8254 & n8260 ) ;
  assign n8262 = ( ~n7337 & n8077 ) | ( ~n7337 & n8261 ) | ( n8077 & n8261 ) ;
  assign n8263 = ( ~n7089 & n8237 ) | ( ~n7089 & n8262 ) | ( n8237 & n8262 ) ;
  assign n8264 = ( ~n6858 & n8122 ) | ( ~n6858 & n8263 ) | ( n8122 & n8263 ) ;
  assign n8265 = ( ~n6630 & n8075 ) | ( ~n6630 & n8264 ) | ( n8075 & n8264 ) ;
  assign n8266 = ( ~n6401 & n8080 ) | ( ~n6401 & n8265 ) | ( n8080 & n8265 ) ;
  assign n8267 = ( ~n6171 & n8083 ) | ( ~n6171 & n8266 ) | ( n8083 & n8266 ) ;
  assign n8268 = ( ~n5964 & n8253 ) | ( ~n5964 & n8267 ) | ( n8253 & n8267 ) ;
  assign n8269 = ( ~n5743 & n8258 ) | ( ~n5743 & n8268 ) | ( n8258 & n8268 ) ;
  assign n8270 = ( ~n5527 & n8233 ) | ( ~n5527 & n8269 ) | ( n8233 & n8269 ) ;
  assign n8271 = ( ~n5319 & n8086 ) | ( ~n5319 & n8270 ) | ( n8086 & n8270 ) ;
  assign n8272 = ( ~n5124 & n8125 ) | ( ~n5124 & n8271 ) | ( n8125 & n8271 ) ;
  assign n8273 = ( ~n4915 & n8203 ) | ( ~n4915 & n8272 ) | ( n8203 & n8272 ) ;
  assign n8274 = ( ~n4728 & n8193 ) | ( ~n4728 & n8273 ) | ( n8193 & n8273 ) ;
  assign n8275 = ( ~n4534 & n8089 ) | ( ~n4534 & n8274 ) | ( n8089 & n8274 ) ;
  assign n8276 = ( ~n4346 & n8092 ) | ( ~n4346 & n8275 ) | ( n8092 & n8275 ) ;
  assign n8277 = ( ~n4167 & n8128 ) | ( ~n4167 & n8276 ) | ( n8128 & n8276 ) ;
  assign n8278 = ( ~n3986 & n8131 ) | ( ~n3986 & n8277 ) | ( n8131 & n8277 ) ;
  assign n8279 = ( ~n3804 & n8207 ) | ( ~n3804 & n8278 ) | ( n8207 & n8278 ) ;
  assign n8280 = ( ~n3631 & n8134 ) | ( ~n3631 & n8279 ) | ( n8134 & n8279 ) ;
  assign n8281 = ( ~n3464 & n8095 ) | ( ~n3464 & n8280 ) | ( n8095 & n8280 ) ;
  assign n8282 = ( ~n3302 & n8098 ) | ( ~n3302 & n8281 ) | ( n8098 & n8281 ) ;
  assign n8283 = ( ~n3141 & n8101 ) | ( ~n3141 & n8282 ) | ( n8101 & n8282 ) ;
  assign n8284 = ( ~n2995 & n8104 ) | ( ~n2995 & n8283 ) | ( n8104 & n8283 ) ;
  assign n8285 = ( ~n2839 & n8107 ) | ( ~n2839 & n8284 ) | ( n8107 & n8284 ) ;
  assign n8286 = ( ~n2690 & n8137 ) | ( ~n2690 & n8285 ) | ( n8137 & n8285 ) ;
  assign n8287 = ( ~n2544 & n8220 ) | ( ~n2544 & n8286 ) | ( n8220 & n8286 ) ;
  assign n8288 = ( ~n2404 & n8140 ) | ( ~n2404 & n8287 ) | ( n8140 & n8287 ) ;
  assign n8289 = ( ~n2269 & n8197 ) | ( ~n2269 & n8288 ) | ( n8197 & n8288 ) ;
  assign n8290 = ( ~n2139 & n8223 ) | ( ~n2139 & n8289 ) | ( n8223 & n8289 ) ;
  assign n8291 = ( ~n2009 & n8214 ) | ( ~n2009 & n8290 ) | ( n8214 & n8290 ) ;
  assign n8292 = ( ~n1885 & n8212 ) | ( ~n1885 & n8291 ) | ( n8212 & n8291 ) ;
  assign n8293 = ( ~n1766 & n8110 ) | ( ~n1766 & n8292 ) | ( n8110 & n8292 ) ;
  assign n8294 = ( ~n1652 & n8143 ) | ( ~n1652 & n8293 ) | ( n8143 & n8293 ) ;
  assign n8295 = ( ~n1534 & n8113 ) | ( ~n1534 & n8294 ) | ( n8113 & n8294 ) ;
  assign n8296 = ( ~n1416 & n8146 ) | ( ~n1416 & n8295 ) | ( n8146 & n8295 ) ;
  assign n8297 = ( ~n1318 & n8221 ) | ( ~n1318 & n8296 ) | ( n8221 & n8296 ) ;
  assign n8298 = ( ~n1220 & n8222 ) | ( ~n1220 & n8297 ) | ( n8222 & n8297 ) ;
  assign n8299 = ( ~n1118 & n8149 ) | ( ~n1118 & n8298 ) | ( n8149 & n8298 ) ;
  assign n8300 = ( ~n1034 & n8152 ) | ( ~n1034 & n8299 ) | ( n8152 & n8299 ) ;
  assign n8301 = ( ~n941 & n8195 ) | ( ~n941 & n8300 ) | ( n8195 & n8300 ) ;
  assign n8302 = ( ~n859 & n8155 ) | ( ~n859 & n8301 ) | ( n8155 & n8301 ) ;
  assign n8303 = ( ~n785 & n8158 ) | ( ~n785 & n8302 ) | ( n8158 & n8302 ) ;
  assign n8304 = ( ~n716 & n8161 ) | ( ~n716 & n8303 ) | ( n8161 & n8303 ) ;
  assign n8305 = n8263 ^ n6858 ^ 1'b0 ;
  assign n8306 = n8287 ^ n2404 ^ 1'b0 ;
  assign n8307 = n8303 ^ n716 ^ 1'b0 ;
  assign n8308 = ( ~n640 & n8199 ) | ( ~n640 & n8304 ) | ( n8199 & n8304 ) ;
  assign n8309 = ( ~n572 & n8201 ) | ( ~n572 & n8308 ) | ( n8201 & n8308 ) ;
  assign n8310 = ( ~n514 & n8164 ) | ( ~n514 & n8309 ) | ( n8164 & n8309 ) ;
  assign n8311 = ( ~n458 & n8167 ) | ( ~n458 & n8310 ) | ( n8167 & n8310 ) ;
  assign n8312 = ( ~n399 & n8224 ) | ( ~n399 & n8311 ) | ( n8224 & n8311 ) ;
  assign n8313 = ( ~n345 & n8170 ) | ( ~n345 & n8312 ) | ( n8170 & n8312 ) ;
  assign n8314 = ( ~n302 & n8116 ) | ( ~n302 & n8313 ) | ( n8116 & n8313 ) ;
  assign n8315 = ( ~n261 & n8229 ) | ( ~n261 & n8314 ) | ( n8229 & n8314 ) ;
  assign n8316 = ( ~n217 & n8173 ) | ( ~n217 & n8315 ) | ( n8173 & n8315 ) ;
  assign n8317 = ( ~n179 & n8210 ) | ( ~n179 & n8316 ) | ( n8210 & n8316 ) ;
  assign n8318 = ( ~n144 & n8176 ) | ( ~n144 & n8317 ) | ( n8176 & n8317 ) ;
  assign n8319 = ( ~n134 & n8119 ) | ( ~n134 & n8318 ) | ( n8119 & n8318 ) ;
  assign n8320 = n8072 & n8319 ;
  assign n8321 = n8245 | n8320 ;
  assign n8322 = ~n136 & n8319 ;
  assign n8323 = ( ~n136 & n8249 ) | ( ~n136 & n8322 ) | ( n8249 & n8322 ) ;
  assign n8324 = n8321 | n8323 ;
  assign n8325 = ( n8069 & n8320 ) | ( n8069 & ~n8323 ) | ( n8320 & ~n8323 ) ;
  assign n8326 = ~n8228 & n8324 ;
  assign n8327 = n8321 & ~n8326 ;
  assign n8328 = ( n8325 & n8326 ) | ( n8325 & ~n8327 ) | ( n8326 & ~n8327 ) ;
  assign n8329 = ( n8217 & ~n8235 ) | ( n8217 & n8324 ) | ( ~n8235 & n8324 ) ;
  assign n8330 = ~n8217 & n8329 ;
  assign n8331 = n8305 & n8324 ;
  assign n8332 = n8331 ^ n8324 ^ n8122 ;
  assign n8333 = n8324 ^ n8267 ^ n5964 ;
  assign n8334 = n8324 & n8333 ;
  assign n8335 = n8334 ^ n8251 ^ n7951 ;
  assign n8336 = n8324 ^ n8272 ^ n4915 ;
  assign n8337 = n8324 & n8336 ;
  assign n8338 = n8337 ^ n8202 ^ n7889 ;
  assign n8339 = n8324 ^ n8281 ^ n3302 ;
  assign n8340 = n8324 & n8339 ;
  assign n8341 = n8340 ^ n8097 ^ n7906 ;
  assign n8342 = n8306 & n8324 ;
  assign n8343 = n8342 ^ n8324 ^ n8140 ;
  assign n8344 = n8324 ^ n8288 ^ n2269 ;
  assign n8345 = n8324 & n8344 ;
  assign n8346 = n8345 ^ n8196 ^ n7909 ;
  assign n8347 = n8324 ^ n8289 ^ n2139 ;
  assign n8348 = n8324 & n8347 ;
  assign n8349 = n8348 ^ n8206 ^ n7977 ;
  assign n8350 = n8324 ^ n8297 ^ n1220 ;
  assign n8351 = n8324 & n8350 ;
  assign n8352 = n8351 ^ n8219 ^ n7915 ;
  assign n8353 = n8307 & n8324 ;
  assign n8354 = n8353 ^ n8324 ^ n8161 ;
  assign n8355 = n8324 ^ n8304 ^ n640 ;
  assign n8356 = n8324 & n8355 ;
  assign n8357 = n8356 ^ n8198 ^ n7865 ;
  assign n8358 = n8324 ^ n8309 ^ n514 ;
  assign n8359 = n8324 & n8358 ;
  assign n8360 = n8359 ^ n8163 ^ n7933 ;
  assign n8361 = n8324 ^ n8318 ^ n134 ;
  assign n8362 = n8324 & n8361 ;
  assign n8363 = n8362 ^ n8118 ^ n7877 ;
  assign n8364 = n8324 ^ n8268 ^ n5743 ;
  assign n8365 = n8324 ^ n8270 ^ n5319 ;
  assign n8366 = n8324 & n8365 ;
  assign n8367 = n8366 ^ n8085 ^ n7886 ;
  assign n8368 = n8324 ^ n8291 ^ n1885 ;
  assign n8369 = n8324 & n8368 ;
  assign n8370 = n8369 ^ n8211 ^ n7912 ;
  assign n8371 = n8324 ^ n8292 ^ n1766 ;
  assign n8372 = n8324 & n8371 ;
  assign n8373 = n8372 ^ n8109 ^ n7847 ;
  assign n8374 = n8324 ^ n8300 ^ n941 ;
  assign n8375 = n8324 & n8374 ;
  assign n8376 = n8375 ^ n8194 ^ n7924 ;
  assign n8377 = n8301 ^ n859 ^ 1'b0 ;
  assign n8378 = n8324 & n8377 ;
  assign n8379 = n8378 ^ n8324 ^ n8155 ;
  assign n8380 = n8324 ^ n8302 ^ n785 ;
  assign n8381 = n8324 & n8364 ;
  assign n8382 = n8381 ^ n8256 ^ n7898 ;
  assign n8383 = n8324 & n8380 ;
  assign n8384 = n8383 ^ n8157 ^ n7927 ;
  assign n8385 = n8324 ^ n8308 ^ n572 ;
  assign n8386 = n8324 ^ n8310 ^ n458 ;
  assign n8387 = n8324 & n8386 ;
  assign n8388 = n8387 ^ n8166 ^ n7936 ;
  assign n8389 = n8324 ^ n8311 ^ n399 ;
  assign n8390 = n8312 ^ n345 ^ 1'b0 ;
  assign n8391 = n8324 & n8390 ;
  assign n8392 = n8391 ^ n8324 ^ n8170 ;
  assign n8393 = n8324 ^ n8313 ^ n302 ;
  assign n8394 = n8324 & n8393 ;
  assign n8395 = n8394 ^ n8115 ^ n7876 ;
  assign n8396 = n8324 & n8389 ;
  assign n8397 = n8396 ^ n8205 ^ n7860 ;
  assign n8398 = n8314 ^ n261 ^ 1'b0 ;
  assign n8399 = n8324 & n8398 ;
  assign n8400 = n8399 ^ n8324 ^ n8229 ;
  assign n8401 = n8324 ^ n8315 ^ n217 ;
  assign n8402 = n8324 & n8401 ;
  assign n8403 = n8402 ^ n8172 ^ n7878 ;
  assign n8404 = n8324 ^ n8316 ^ n179 ;
  assign n8405 = n8324 & n8404 ;
  assign n8406 = n8405 ^ n8209 ^ n7879 ;
  assign n8407 = n8324 ^ n8317 ^ n144 ;
  assign n8408 = n8324 & n8407 ;
  assign n8409 = n8408 ^ n8175 ^ n7875 ;
  assign n8410 = n8324 ^ n8266 ^ n6171 ;
  assign n8411 = n8324 & n8410 ;
  assign n8412 = n8411 ^ n8082 ^ n7948 ;
  assign n8413 = n8261 ^ n7337 ^ 1'b0 ;
  assign n8414 = n8324 & n8413 ;
  assign n8415 = n8414 ^ n8324 ^ n8077 ;
  assign n8416 = n8324 ^ n8264 ^ n6630 ;
  assign n8417 = n8324 & n8416 ;
  assign n8418 = n8417 ^ n8074 ^ n7945 ;
  assign n8419 = n8324 ^ n8265 ^ n6401 ;
  assign n8420 = n8324 & n8419 ;
  assign n8421 = n8420 ^ n8079 ^ n7882 ;
  assign n8422 = n8269 ^ n5527 ^ 1'b0 ;
  assign n8423 = n8324 & n8422 ;
  assign n8424 = n8423 ^ n8324 ^ n8233 ;
  assign n8425 = n8271 ^ n5124 ^ 1'b0 ;
  assign n8426 = n8324 & n8425 ;
  assign n8427 = n8426 ^ n8324 ^ n8125 ;
  assign n8428 = n8324 ^ n8275 ^ n4346 ;
  assign n8429 = n8324 & n8428 ;
  assign n8430 = n8429 ^ n8091 ^ n7900 ;
  assign n8431 = n8277 ^ n3986 ^ 1'b0 ;
  assign n8432 = n8324 & n8431 ;
  assign n8433 = n8432 ^ n8324 ^ n8131 ;
  assign n8434 = n8279 ^ n3631 ^ 1'b0 ;
  assign n8435 = n8324 ^ n8283 ^ n2995 ;
  assign n8436 = n8324 & n8435 ;
  assign n8437 = n8436 ^ n8103 ^ n7873 ;
  assign n8438 = n8285 ^ n2690 ^ 1'b0 ;
  assign n8439 = n8324 & n8438 ;
  assign n8440 = n8439 ^ n8324 ^ n8137 ;
  assign n8441 = n8324 ^ n8290 ^ n2009 ;
  assign n8442 = n8324 & n8441 ;
  assign n8443 = n8324 & n8434 ;
  assign n8444 = n8443 ^ n8324 ^ n8134 ;
  assign n8445 = n8442 ^ n8213 ^ n7851 ;
  assign n8446 = n8293 ^ n1652 ^ 1'b0 ;
  assign n8447 = n8324 & n8446 ;
  assign n8448 = n8447 ^ n8324 ^ n8143 ;
  assign n8449 = n8295 ^ n1416 ^ 1'b0 ;
  assign n8450 = n8324 & n8449 ;
  assign n8451 = n8450 ^ n8324 ^ n8146 ;
  assign n8452 = n8324 ^ n8298 ^ n1118 ;
  assign n8453 = n8324 ^ n8299 ^ n1034 ;
  assign n8454 = n8324 & n8385 ;
  assign n8455 = n8454 ^ n8200 ^ n7840 ;
  assign n8456 = ( x116 & n8066 ) | ( x116 & n8324 ) | ( n8066 & n8324 ) ;
  assign n8457 = n8324 ^ n8262 ^ n7089 ;
  assign n8458 = n8324 & n8457 ;
  assign n8459 = n8458 ^ n8236 ^ n7997 ;
  assign n8460 = n8324 ^ n8273 ^ n4728 ;
  assign n8461 = n8324 & n8460 ;
  assign n8462 = n8461 ^ n8192 ^ n7892 ;
  assign n8463 = n8324 ^ n8274 ^ n4534 ;
  assign n8464 = n8324 & n8463 ;
  assign n8465 = n8464 ^ n8088 ^ n7895 ;
  assign n8466 = n8324 ^ n8276 ^ n4167 ;
  assign n8467 = n8324 & n8466 ;
  assign n8468 = n8467 ^ n8127 ^ n7871 ;
  assign n8469 = n8324 ^ n8278 ^ n3804 ;
  assign n8470 = n8324 & n8469 ;
  assign n8471 = n8470 ^ n8204 ^ n7962 ;
  assign n8472 = n8324 ^ n8280 ^ n3464 ;
  assign n8473 = n8324 & n8472 ;
  assign n8474 = n8473 ^ n8094 ^ n7903 ;
  assign n8475 = n8324 ^ n8282 ^ n3141 ;
  assign n8476 = n8324 & n8475 ;
  assign n8477 = n8476 ^ n8100 ^ n7870 ;
  assign n8478 = n8324 ^ n8284 ^ n2839 ;
  assign n8479 = n8324 & n8478 ;
  assign n8480 = n8479 ^ n8106 ^ n7864 ;
  assign n8481 = n8324 ^ n8286 ^ n2544 ;
  assign n8482 = n8324 & n8481 ;
  assign n8483 = n8482 ^ n8208 ^ n7971 ;
  assign n8484 = n8324 ^ n8294 ^ n1534 ;
  assign n8485 = n8324 & n8484 ;
  assign n8486 = n8485 ^ n8112 ^ n7874 ;
  assign n8487 = n8324 ^ n8296 ^ n1318 ;
  assign n8488 = n8324 & n8487 ;
  assign n8489 = n8488 ^ n8218 ^ n7854 ;
  assign n8490 = n8324 & n8452 ;
  assign n8491 = n8490 ^ n8148 ^ n7918 ;
  assign n8492 = n8324 & n8453 ;
  assign n8493 = n8492 ^ n8151 ^ n7921 ;
  assign n8494 = x94 | x105 ;
  assign n8495 = ~x116 & n8324 ;
  assign n8496 = n8324 ^ n8260 ^ n7575 ;
  assign n8497 = ( x116 & ~n7995 ) | ( x116 & n8494 ) | ( ~n7995 & n8494 ) ;
  assign n8498 = n8495 ^ x127 ^ 1'b0 ;
  assign n8499 = ( ~x116 & n8069 ) | ( ~x116 & n8324 ) | ( n8069 & n8324 ) ;
  assign n8500 = n8324 & n8496 ;
  assign n8501 = ( x116 & n8069 ) | ( x116 & ~n8494 ) | ( n8069 & ~n8494 ) ;
  assign n8502 = n8500 ^ n8242 ^ x31 ;
  assign n8503 = n8330 ^ n8252 ^ x22 ;
  assign n8504 = n8499 & n8501 ;
  assign n8505 = ( ~n8069 & n8456 ) | ( ~n8069 & n8497 ) | ( n8456 & n8497 ) ;
  assign n8506 = ~n8456 & n8505 ;
  assign n8507 = n8072 & ~n8319 ;
  assign n8508 = n8498 | n8506 ;
  assign n8509 = ~n8504 & n8508 ;
  assign n8510 = n8328 ^ x11 ^ 1'b0 ;
  assign n8511 = ( ~n7824 & n8509 ) | ( ~n7824 & n8510 ) | ( n8509 & n8510 ) ;
  assign n8512 = ( ~n7575 & n8503 ) | ( ~n7575 & n8511 ) | ( n8503 & n8511 ) ;
  assign n8513 = ( ~n7337 & n8502 ) | ( ~n7337 & n8512 ) | ( n8502 & n8512 ) ;
  assign n8514 = ( ~n7089 & n8415 ) | ( ~n7089 & n8513 ) | ( n8415 & n8513 ) ;
  assign n8515 = ( ~n6858 & n8459 ) | ( ~n6858 & n8514 ) | ( n8459 & n8514 ) ;
  assign n8516 = ( ~n6630 & n8332 ) | ( ~n6630 & n8515 ) | ( n8332 & n8515 ) ;
  assign n8517 = ( ~n6401 & n8418 ) | ( ~n6401 & n8516 ) | ( n8418 & n8516 ) ;
  assign n8518 = ( ~n6171 & n8421 ) | ( ~n6171 & n8517 ) | ( n8421 & n8517 ) ;
  assign n8519 = ( ~n5964 & n8412 ) | ( ~n5964 & n8518 ) | ( n8412 & n8518 ) ;
  assign n8520 = ( ~n5743 & n8335 ) | ( ~n5743 & n8519 ) | ( n8335 & n8519 ) ;
  assign n8521 = ( ~n5527 & n8382 ) | ( ~n5527 & n8520 ) | ( n8382 & n8520 ) ;
  assign n8522 = ( ~n5319 & n8424 ) | ( ~n5319 & n8521 ) | ( n8424 & n8521 ) ;
  assign n8523 = ( ~n5124 & n8367 ) | ( ~n5124 & n8522 ) | ( n8367 & n8522 ) ;
  assign n8524 = ( ~n4915 & n8427 ) | ( ~n4915 & n8523 ) | ( n8427 & n8523 ) ;
  assign n8525 = ( ~n4728 & n8338 ) | ( ~n4728 & n8524 ) | ( n8338 & n8524 ) ;
  assign n8526 = ( ~n4534 & n8462 ) | ( ~n4534 & n8525 ) | ( n8462 & n8525 ) ;
  assign n8527 = ( ~n4346 & n8465 ) | ( ~n4346 & n8526 ) | ( n8465 & n8526 ) ;
  assign n8528 = ( ~n4167 & n8430 ) | ( ~n4167 & n8527 ) | ( n8430 & n8527 ) ;
  assign n8529 = ( ~n3986 & n8468 ) | ( ~n3986 & n8528 ) | ( n8468 & n8528 ) ;
  assign n8530 = ( ~n3804 & n8433 ) | ( ~n3804 & n8529 ) | ( n8433 & n8529 ) ;
  assign n8531 = ( ~n3631 & n8471 ) | ( ~n3631 & n8530 ) | ( n8471 & n8530 ) ;
  assign n8532 = ( ~n3464 & n8444 ) | ( ~n3464 & n8531 ) | ( n8444 & n8531 ) ;
  assign n8533 = ( ~n3302 & n8474 ) | ( ~n3302 & n8532 ) | ( n8474 & n8532 ) ;
  assign n8534 = ( ~n3141 & n8341 ) | ( ~n3141 & n8533 ) | ( n8341 & n8533 ) ;
  assign n8535 = ( ~n2995 & n8477 ) | ( ~n2995 & n8534 ) | ( n8477 & n8534 ) ;
  assign n8536 = ( ~n2839 & n8437 ) | ( ~n2839 & n8535 ) | ( n8437 & n8535 ) ;
  assign n8537 = ( ~n2690 & n8480 ) | ( ~n2690 & n8536 ) | ( n8480 & n8536 ) ;
  assign n8538 = ( ~n2544 & n8440 ) | ( ~n2544 & n8537 ) | ( n8440 & n8537 ) ;
  assign n8539 = ( ~n2404 & n8483 ) | ( ~n2404 & n8538 ) | ( n8483 & n8538 ) ;
  assign n8540 = ( n8072 & ~n8319 ) | ( n8072 & n8324 ) | ( ~n8319 & n8324 ) ;
  assign n8541 = ( ~n2269 & n8343 ) | ( ~n2269 & n8539 ) | ( n8343 & n8539 ) ;
  assign n8542 = ( ~n2139 & n8346 ) | ( ~n2139 & n8541 ) | ( n8346 & n8541 ) ;
  assign n8543 = ( ~n2009 & n8349 ) | ( ~n2009 & n8542 ) | ( n8349 & n8542 ) ;
  assign n8544 = ( ~n1885 & n8445 ) | ( ~n1885 & n8543 ) | ( n8445 & n8543 ) ;
  assign n8545 = ( ~n1766 & n8370 ) | ( ~n1766 & n8544 ) | ( n8370 & n8544 ) ;
  assign n8546 = ( ~n1652 & n8373 ) | ( ~n1652 & n8545 ) | ( n8373 & n8545 ) ;
  assign n8547 = ( ~n1534 & n8448 ) | ( ~n1534 & n8546 ) | ( n8448 & n8546 ) ;
  assign n8548 = ( ~n1416 & n8486 ) | ( ~n1416 & n8547 ) | ( n8486 & n8547 ) ;
  assign n8549 = n8523 ^ n4915 ^ 1'b0 ;
  assign n8550 = n8537 ^ n2544 ^ 1'b0 ;
  assign n8551 = n8521 ^ n5319 ^ 1'b0 ;
  assign n8552 = n8539 ^ n2269 ^ 1'b0 ;
  assign n8553 = n8529 ^ n3804 ^ 1'b0 ;
  assign n8554 = ( ~n1318 & n8451 ) | ( ~n1318 & n8548 ) | ( n8451 & n8548 ) ;
  assign n8555 = ( ~n1220 & n8489 ) | ( ~n1220 & n8554 ) | ( n8489 & n8554 ) ;
  assign n8556 = ( ~n1118 & n8352 ) | ( ~n1118 & n8555 ) | ( n8352 & n8555 ) ;
  assign n8557 = n8513 ^ n7089 ^ 1'b0 ;
  assign n8558 = n8546 ^ n1534 ^ 1'b0 ;
  assign n8559 = n8515 ^ n6630 ^ 1'b0 ;
  assign n8560 = n8548 ^ n1318 ^ 1'b0 ;
  assign n8561 = ( n8363 & ~n8507 ) | ( n8363 & n8540 ) | ( ~n8507 & n8540 ) ;
  assign n8562 = ( n136 & n8072 ) | ( n136 & n8319 ) | ( n8072 & n8319 ) ;
  assign n8563 = n8531 ^ n3464 ^ 1'b0 ;
  assign n8564 = ( ~n1034 & n8491 ) | ( ~n1034 & n8556 ) | ( n8491 & n8556 ) ;
  assign n8565 = ( ~n941 & n8493 ) | ( ~n941 & n8564 ) | ( n8493 & n8564 ) ;
  assign n8566 = ( ~n859 & n8376 ) | ( ~n859 & n8565 ) | ( n8376 & n8565 ) ;
  assign n8567 = ( ~n785 & n8379 ) | ( ~n785 & n8566 ) | ( n8379 & n8566 ) ;
  assign n8568 = ( ~n716 & n8384 ) | ( ~n716 & n8567 ) | ( n8384 & n8567 ) ;
  assign n8569 = ( ~n640 & n8354 ) | ( ~n640 & n8568 ) | ( n8354 & n8568 ) ;
  assign n8570 = ( ~n572 & n8357 ) | ( ~n572 & n8569 ) | ( n8357 & n8569 ) ;
  assign n8571 = ( ~n514 & n8455 ) | ( ~n514 & n8570 ) | ( n8455 & n8570 ) ;
  assign n8572 = ( ~n458 & n8360 ) | ( ~n458 & n8571 ) | ( n8360 & n8571 ) ;
  assign n8573 = ( ~n399 & n8388 ) | ( ~n399 & n8572 ) | ( n8388 & n8572 ) ;
  assign n8574 = ( ~n345 & n8397 ) | ( ~n345 & n8573 ) | ( n8397 & n8573 ) ;
  assign n8575 = ( ~n302 & n8392 ) | ( ~n302 & n8574 ) | ( n8392 & n8574 ) ;
  assign n8576 = ( ~n261 & n8395 ) | ( ~n261 & n8575 ) | ( n8395 & n8575 ) ;
  assign n8577 = ( ~n217 & n8400 ) | ( ~n217 & n8576 ) | ( n8400 & n8576 ) ;
  assign n8578 = ( ~n179 & n8403 ) | ( ~n179 & n8577 ) | ( n8403 & n8577 ) ;
  assign n8579 = ( ~n144 & n8406 ) | ( ~n144 & n8578 ) | ( n8406 & n8578 ) ;
  assign n8580 = ( ~n134 & n8409 ) | ( ~n134 & n8579 ) | ( n8409 & n8579 ) ;
  assign n8581 = n8363 & n8580 ;
  assign n8582 = ( ~n8072 & n8324 ) | ( ~n8072 & n8581 ) | ( n8324 & n8581 ) ;
  assign n8583 = n8319 & ~n8582 ;
  assign n8584 = ( ~x30 & n8561 ) | ( ~x30 & n8580 ) | ( n8561 & n8580 ) ;
  assign n8585 = ~n136 & n8584 ;
  assign n8586 = ( n8562 & n8581 ) | ( n8562 & ~n8583 ) | ( n8581 & ~n8583 ) ;
  assign n8587 = n8585 | n8586 ;
  assign n8588 = n8553 & n8587 ;
  assign n8589 = n8587 ^ n8579 ^ n134 ;
  assign n8590 = ~n8494 & n8587 ;
  assign n8591 = n8560 & n8587 ;
  assign n8592 = n8591 ^ n8587 ^ n8451 ;
  assign n8593 = n8558 & n8587 ;
  assign n8594 = n8550 & n8587 ;
  assign n8595 = n8593 ^ n8587 ^ n8448 ;
  assign n8596 = n8594 ^ n8587 ^ n8440 ;
  assign n8597 = n8552 & n8587 ;
  assign n8598 = n8597 ^ n8587 ^ n8343 ;
  assign n8599 = n8557 & n8587 ;
  assign n8600 = ( ~n8504 & n8506 ) | ( ~n8504 & n8587 ) | ( n8506 & n8587 ) ;
  assign n8601 = ( n8324 & n8581 ) | ( n8324 & ~n8585 ) | ( n8581 & ~n8585 ) ;
  assign n8602 = n8599 ^ n8587 ^ n8415 ;
  assign n8603 = n8587 ^ n8516 ^ n6401 ;
  assign n8604 = n8587 & n8589 ;
  assign n8605 = n8559 & n8587 ;
  assign n8606 = n8586 & ~n8590 ;
  assign n8607 = n8605 ^ n8587 ^ n8332 ;
  assign n8608 = n8563 & n8587 ;
  assign n8609 = n8551 & n8587 ;
  assign n8610 = n8549 & n8587 ;
  assign n8611 = n8609 ^ n8587 ^ n8424 ;
  assign n8612 = n8610 ^ n8587 ^ n8427 ;
  assign n8613 = n8608 ^ n8587 ^ n8444 ;
  assign n8614 = n8604 ^ n8408 ^ n8176 ;
  assign n8615 = n8587 & n8603 ;
  assign n8616 = n8615 ^ n8417 ^ n8075 ;
  assign n8617 = ( n8590 & n8601 ) | ( n8590 & ~n8606 ) | ( n8601 & ~n8606 ) ;
  assign n8618 = ~n8506 & n8600 ;
  assign n8619 = n8588 ^ n8587 ^ n8433 ;
  assign n8620 = n8587 ^ n8534 ^ n2995 ;
  assign n8621 = n8587 ^ n8524 ^ n4728 ;
  assign n8622 = n8587 ^ n8545 ^ n1652 ;
  assign n8623 = n8587 ^ n8517 ^ n6171 ;
  assign n8624 = n8587 ^ n8535 ^ n2839 ;
  assign n8625 = n8587 ^ n8527 ^ n4167 ;
  assign n8626 = n8587 ^ n8536 ^ n2690 ;
  assign n8627 = n8587 ^ n8556 ^ n1034 ;
  assign n8628 = n8587 ^ n8541 ^ n2139 ;
  assign n8629 = n8587 ^ n8533 ^ n3141 ;
  assign n8630 = n8587 ^ n8573 ^ n345 ;
  assign n8631 = n8587 ^ n8538 ^ n2404 ;
  assign n8632 = n8587 ^ n8555 ^ n1118 ;
  assign n8633 = n8587 ^ n8565 ^ n859 ;
  assign n8634 = n8587 ^ n8532 ^ n3302 ;
  assign n8635 = n8587 & n8625 ;
  assign n8636 = n8635 ^ n8429 ^ n8092 ;
  assign n8637 = n8587 & n8622 ;
  assign n8638 = n8637 ^ n8372 ^ n8110 ;
  assign n8639 = n8587 & n8632 ;
  assign n8640 = n8639 ^ n8351 ^ n8222 ;
  assign n8641 = n8587 & n8624 ;
  assign n8642 = n8641 ^ n8436 ^ n8104 ;
  assign n8643 = n8587 & n8630 ;
  assign n8644 = n8587 & n8627 ;
  assign n8645 = n8644 ^ n8490 ^ n8149 ;
  assign n8646 = n8587 & n8621 ;
  assign n8647 = n8646 ^ n8337 ^ n8203 ;
  assign n8648 = n8587 & n8629 ;
  assign n8649 = n8587 & n8623 ;
  assign n8650 = n8643 ^ n8396 ^ n8224 ;
  assign n8651 = n8649 ^ n8420 ^ n8080 ;
  assign n8652 = n8587 & n8620 ;
  assign n8653 = n8652 ^ n8476 ^ n8101 ;
  assign n8654 = n8587 & n8633 ;
  assign n8655 = n8654 ^ n8375 ^ n8195 ;
  assign n8656 = n8587 & n8634 ;
  assign n8657 = n8656 ^ n8473 ^ n8095 ;
  assign n8658 = n8587 & n8626 ;
  assign n8659 = n8587 & n8628 ;
  assign n8660 = n8659 ^ n8345 ^ n8197 ;
  assign n8661 = n8658 ^ n8479 ^ n8107 ;
  assign n8662 = n8587 & n8631 ;
  assign n8663 = n8662 ^ n8482 ^ n8220 ;
  assign n8664 = n8648 ^ n8340 ^ n8098 ;
  assign n8665 = n8587 ^ n8511 ^ n7575 ;
  assign n8666 = n8587 & n8665 ;
  assign n8667 = n8666 ^ n8330 ^ n8257 ;
  assign n8668 = n8587 ^ n8522 ^ n5124 ;
  assign n8669 = n8587 & n8668 ;
  assign n8670 = n8669 ^ n8366 ^ n8086 ;
  assign n8671 = n8587 ^ n8525 ^ n4534 ;
  assign n8672 = n8587 & n8671 ;
  assign n8673 = n8672 ^ n8461 ^ n8193 ;
  assign n8674 = n8587 ^ n8530 ^ n3631 ;
  assign n8675 = n8587 & n8674 ;
  assign n8676 = n8675 ^ n8470 ^ n8207 ;
  assign n8677 = n8587 ^ n8543 ^ n1885 ;
  assign n8678 = n8587 & n8677 ;
  assign n8679 = n8587 ^ n8544 ^ n1766 ;
  assign n8680 = n8587 & n8679 ;
  assign n8681 = n8680 ^ n8369 ^ n8212 ;
  assign n8682 = n8587 ^ n8547 ^ n1416 ;
  assign n8683 = n8587 & n8682 ;
  assign n8684 = n8683 ^ n8485 ^ n8113 ;
  assign n8685 = n8587 ^ n8564 ^ n941 ;
  assign n8686 = n8587 & n8685 ;
  assign n8687 = n8686 ^ n8492 ^ n8152 ;
  assign n8688 = n8566 ^ n785 ^ 1'b0 ;
  assign n8689 = n8587 & n8688 ;
  assign n8690 = n8689 ^ n8587 ^ n8379 ;
  assign n8691 = n8568 ^ n640 ^ 1'b0 ;
  assign n8692 = n8587 & n8691 ;
  assign n8693 = n8692 ^ n8587 ^ n8354 ;
  assign n8694 = n8587 ^ n8518 ^ n5964 ;
  assign n8695 = n8587 & n8694 ;
  assign n8696 = n8695 ^ n8411 ^ n8083 ;
  assign n8697 = n8587 ^ n8570 ^ n514 ;
  assign n8698 = n8587 & n8697 ;
  assign n8699 = n8678 ^ n8442 ^ n8214 ;
  assign n8700 = n8698 ^ n8454 ^ n8201 ;
  assign n8701 = n8587 ^ n8571 ^ n458 ;
  assign n8702 = n8587 & n8701 ;
  assign n8703 = n8702 ^ n8359 ^ n8164 ;
  assign n8704 = n8574 ^ n302 ^ 1'b0 ;
  assign n8705 = n8587 & n8704 ;
  assign n8706 = n8705 ^ n8587 ^ n8392 ;
  assign n8707 = n8576 ^ n217 ^ 1'b0 ;
  assign n8708 = n8587 & n8707 ;
  assign n8709 = n8708 ^ n8587 ^ n8400 ;
  assign n8710 = n8587 ^ n8578 ^ n144 ;
  assign n8711 = n8587 & n8710 ;
  assign n8712 = n8711 ^ n8405 ^ n8210 ;
  assign n8713 = n8587 ^ n8514 ^ n6858 ;
  assign n8714 = n8587 ^ n8526 ^ n4346 ;
  assign n8715 = n8587 ^ n8542 ^ n2009 ;
  assign n8716 = n8587 ^ n8554 ^ n1220 ;
  assign n8717 = n8587 ^ n8520 ^ n5527 ;
  assign n8718 = n8587 ^ n8519 ^ n5743 ;
  assign n8719 = n8587 ^ n8567 ^ n716 ;
  assign n8720 = n8587 ^ n8528 ^ n3986 ;
  assign n8721 = n8587 ^ n8572 ^ n399 ;
  assign n8722 = n8587 ^ n8577 ^ n179 ;
  assign n8723 = n8587 ^ n8512 ^ n7337 ;
  assign n8724 = n8587 ^ n8569 ^ n572 ;
  assign n8725 = n8587 ^ n8575 ^ n261 ;
  assign n8726 = n8587 & n8716 ;
  assign n8727 = n8587 & n8715 ;
  assign n8728 = n8587 & n8719 ;
  assign n8729 = n8728 ^ n8383 ^ n8158 ;
  assign n8730 = n8587 & n8721 ;
  assign n8731 = n8730 ^ n8387 ^ n8167 ;
  assign n8732 = n8587 & n8724 ;
  assign n8733 = n8732 ^ n8356 ^ n8199 ;
  assign n8734 = n8587 & n8725 ;
  assign n8735 = n8587 & n8720 ;
  assign n8736 = n8727 ^ n8348 ^ n8223 ;
  assign n8737 = n8587 & n8713 ;
  assign n8738 = n8737 ^ n8458 ^ n8237 ;
  assign n8739 = n8735 ^ n8467 ^ n8128 ;
  assign n8740 = n8587 & n8714 ;
  assign n8741 = n8740 ^ n8464 ^ n8089 ;
  assign n8742 = n8587 & n8717 ;
  assign n8743 = n8742 ^ n8381 ^ n8258 ;
  assign n8744 = n8734 ^ n8394 ^ n8116 ;
  assign n8745 = n8587 & n8722 ;
  assign n8746 = n8587 & n8718 ;
  assign n8747 = n8745 ^ n8402 ^ n8173 ;
  assign n8748 = n8587 & n8723 ;
  assign n8749 = n8748 ^ n8500 ^ n8254 ;
  assign n8750 = n8746 ^ n8334 ^ n8253 ;
  assign n8751 = ~x94 & n8587 ;
  assign n8752 = n8751 ^ x105 ^ 1'b0 ;
  assign n8753 = n8617 ^ x116 ^ 1'b0 ;
  assign n8754 = ( ~x94 & n8324 ) | ( ~x94 & n8587 ) | ( n8324 & n8587 ) ;
  assign n8755 = x72 | x83 ;
  assign n8756 = ( x94 & n8324 ) | ( x94 & ~n8755 ) | ( n8324 & ~n8755 ) ;
  assign n8757 = n8754 & n8756 ;
  assign n8758 = ( x94 & ~n8245 ) | ( x94 & n8755 ) | ( ~n8245 & n8755 ) ;
  assign n8759 = ( x94 & n8323 ) | ( x94 & n8587 ) | ( n8323 & n8587 ) ;
  assign n8760 = ( ~n8324 & n8758 ) | ( ~n8324 & n8759 ) | ( n8758 & n8759 ) ;
  assign n8761 = ~n8759 & n8760 ;
  assign n8762 = n8587 ^ n8509 ^ n7824 ;
  assign n8763 = n8587 & n8762 ;
  assign n8764 = n8618 ^ n8495 ^ x127 ;
  assign n8765 = n8752 | n8761 ;
  assign n8766 = ~n8757 & n8765 ;
  assign n8767 = ( ~n8069 & n8753 ) | ( ~n8069 & n8766 ) | ( n8753 & n8766 ) ;
  assign n8768 = ( ~n7824 & n8764 ) | ( ~n7824 & n8767 ) | ( n8764 & n8767 ) ;
  assign n8769 = n8763 ^ n8328 ^ x11 ;
  assign n8770 = ( ~n7575 & n8768 ) | ( ~n7575 & n8769 ) | ( n8768 & n8769 ) ;
  assign n8771 = ( ~n7337 & n8667 ) | ( ~n7337 & n8770 ) | ( n8667 & n8770 ) ;
  assign n8772 = ( ~n7089 & n8749 ) | ( ~n7089 & n8771 ) | ( n8749 & n8771 ) ;
  assign n8773 = ( ~n6858 & n8602 ) | ( ~n6858 & n8772 ) | ( n8602 & n8772 ) ;
  assign n8774 = ( ~n6630 & n8738 ) | ( ~n6630 & n8773 ) | ( n8738 & n8773 ) ;
  assign n8775 = ( ~n6401 & n8607 ) | ( ~n6401 & n8774 ) | ( n8607 & n8774 ) ;
  assign n8776 = ( ~n6171 & n8616 ) | ( ~n6171 & n8775 ) | ( n8616 & n8775 ) ;
  assign n8777 = ( ~n5964 & n8651 ) | ( ~n5964 & n8776 ) | ( n8651 & n8776 ) ;
  assign n8778 = ( ~n5743 & n8696 ) | ( ~n5743 & n8777 ) | ( n8696 & n8777 ) ;
  assign n8779 = ( ~n5527 & n8750 ) | ( ~n5527 & n8778 ) | ( n8750 & n8778 ) ;
  assign n8780 = ( ~n5319 & n8743 ) | ( ~n5319 & n8779 ) | ( n8743 & n8779 ) ;
  assign n8781 = ( ~n5124 & n8611 ) | ( ~n5124 & n8780 ) | ( n8611 & n8780 ) ;
  assign n8782 = ( ~n4915 & n8670 ) | ( ~n4915 & n8781 ) | ( n8670 & n8781 ) ;
  assign n8783 = ( ~n4728 & n8612 ) | ( ~n4728 & n8782 ) | ( n8612 & n8782 ) ;
  assign n8784 = ( ~n4534 & n8647 ) | ( ~n4534 & n8783 ) | ( n8647 & n8783 ) ;
  assign n8785 = ( ~n4346 & n8673 ) | ( ~n4346 & n8784 ) | ( n8673 & n8784 ) ;
  assign n8786 = ( ~n4167 & n8741 ) | ( ~n4167 & n8785 ) | ( n8741 & n8785 ) ;
  assign n8787 = ( ~n3986 & n8636 ) | ( ~n3986 & n8786 ) | ( n8636 & n8786 ) ;
  assign n8788 = ( ~n8363 & n8580 ) | ( ~n8363 & n8587 ) | ( n8580 & n8587 ) ;
  assign n8789 = ( ~n3804 & n8739 ) | ( ~n3804 & n8787 ) | ( n8739 & n8787 ) ;
  assign n8790 = ( ~n3631 & n8619 ) | ( ~n3631 & n8789 ) | ( n8619 & n8789 ) ;
  assign n8791 = n8726 ^ n8488 ^ n8221 ;
  assign n8792 = ( ~n3464 & n8676 ) | ( ~n3464 & n8790 ) | ( n8676 & n8790 ) ;
  assign n8793 = ( ~n3302 & n8613 ) | ( ~n3302 & n8792 ) | ( n8613 & n8792 ) ;
  assign n8794 = ( ~n3141 & n8657 ) | ( ~n3141 & n8793 ) | ( n8657 & n8793 ) ;
  assign n8795 = ( ~n2995 & n8664 ) | ( ~n2995 & n8794 ) | ( n8664 & n8794 ) ;
  assign n8796 = ( ~n2839 & n8653 ) | ( ~n2839 & n8795 ) | ( n8653 & n8795 ) ;
  assign n8797 = ( ~n2690 & n8642 ) | ( ~n2690 & n8796 ) | ( n8642 & n8796 ) ;
  assign n8798 = ( ~n2544 & n8661 ) | ( ~n2544 & n8797 ) | ( n8661 & n8797 ) ;
  assign n8799 = ( ~n2404 & n8596 ) | ( ~n2404 & n8798 ) | ( n8596 & n8798 ) ;
  assign n8800 = ( ~n2269 & n8663 ) | ( ~n2269 & n8799 ) | ( n8663 & n8799 ) ;
  assign n8801 = ~n8363 & n8580 ;
  assign n8802 = ( ~n2139 & n8598 ) | ( ~n2139 & n8800 ) | ( n8598 & n8800 ) ;
  assign n8803 = ( ~n2009 & n8660 ) | ( ~n2009 & n8802 ) | ( n8660 & n8802 ) ;
  assign n8804 = ( ~n1885 & n8736 ) | ( ~n1885 & n8803 ) | ( n8736 & n8803 ) ;
  assign n8805 = ( ~n1766 & n8699 ) | ( ~n1766 & n8804 ) | ( n8699 & n8804 ) ;
  assign n8806 = ( ~n1652 & n8681 ) | ( ~n1652 & n8805 ) | ( n8681 & n8805 ) ;
  assign n8807 = ( ~n1534 & n8638 ) | ( ~n1534 & n8806 ) | ( n8638 & n8806 ) ;
  assign n8808 = ( ~n1416 & n8595 ) | ( ~n1416 & n8807 ) | ( n8595 & n8807 ) ;
  assign n8809 = ( ~n1318 & n8684 ) | ( ~n1318 & n8808 ) | ( n8684 & n8808 ) ;
  assign n8810 = ( ~n1220 & n8592 ) | ( ~n1220 & n8809 ) | ( n8592 & n8809 ) ;
  assign n8811 = ( ~n1118 & n8791 ) | ( ~n1118 & n8810 ) | ( n8791 & n8810 ) ;
  assign n8812 = ( ~n1034 & n8640 ) | ( ~n1034 & n8811 ) | ( n8640 & n8811 ) ;
  assign n8813 = ( ~n941 & n8645 ) | ( ~n941 & n8812 ) | ( n8645 & n8812 ) ;
  assign n8814 = ( ~n859 & n8687 ) | ( ~n859 & n8813 ) | ( n8687 & n8813 ) ;
  assign n8815 = ( ~n785 & n8655 ) | ( ~n785 & n8814 ) | ( n8655 & n8814 ) ;
  assign n8816 = ( ~n716 & n8690 ) | ( ~n716 & n8815 ) | ( n8690 & n8815 ) ;
  assign n8817 = ( n8614 & n8788 ) | ( n8614 & ~n8801 ) | ( n8788 & ~n8801 ) ;
  assign n8818 = ( ~n640 & n8729 ) | ( ~n640 & n8816 ) | ( n8729 & n8816 ) ;
  assign n8819 = ( ~n572 & n8693 ) | ( ~n572 & n8818 ) | ( n8693 & n8818 ) ;
  assign n8820 = ( ~n514 & n8733 ) | ( ~n514 & n8819 ) | ( n8733 & n8819 ) ;
  assign n8821 = ( ~n458 & n8700 ) | ( ~n458 & n8820 ) | ( n8700 & n8820 ) ;
  assign n8822 = ( ~n399 & n8703 ) | ( ~n399 & n8821 ) | ( n8703 & n8821 ) ;
  assign n8823 = ( ~n345 & n8731 ) | ( ~n345 & n8822 ) | ( n8731 & n8822 ) ;
  assign n8824 = ( ~n302 & n8650 ) | ( ~n302 & n8823 ) | ( n8650 & n8823 ) ;
  assign n8825 = ( ~n261 & n8706 ) | ( ~n261 & n8824 ) | ( n8706 & n8824 ) ;
  assign n8826 = ( ~n217 & n8744 ) | ( ~n217 & n8825 ) | ( n8744 & n8825 ) ;
  assign n8827 = ( ~n179 & n8709 ) | ( ~n179 & n8826 ) | ( n8709 & n8826 ) ;
  assign n8828 = ( ~n144 & n8747 ) | ( ~n144 & n8827 ) | ( n8747 & n8827 ) ;
  assign n8829 = ( ~n134 & n8712 ) | ( ~n134 & n8828 ) | ( n8712 & n8828 ) ;
  assign n8830 = ( ~x30 & n8817 ) | ( ~x30 & n8829 ) | ( n8817 & n8829 ) ;
  assign n8831 = ~n136 & n8830 ;
  assign n8832 = n8614 & n8829 ;
  assign n8833 = ( n136 & n8363 ) | ( n136 & n8580 ) | ( n8363 & n8580 ) ;
  assign n8834 = ( ~n8363 & n8587 ) | ( ~n8363 & n8832 ) | ( n8587 & n8832 ) ;
  assign n8835 = n8580 & ~n8834 ;
  assign n8836 = ( n8832 & n8833 ) | ( n8832 & ~n8835 ) | ( n8833 & ~n8835 ) ;
  assign n8837 = n8831 | n8836 ;
  assign n8838 = ( n8587 & ~n8831 ) | ( n8587 & n8832 ) | ( ~n8831 & n8832 ) ;
  assign n8839 = ~n8755 & n8837 ;
  assign n8840 = n8836 & ~n8839 ;
  assign n8841 = ( n8838 & n8839 ) | ( n8838 & ~n8840 ) | ( n8839 & ~n8840 ) ;
  assign n8842 = ( ~n8757 & n8761 ) | ( ~n8757 & n8837 ) | ( n8761 & n8837 ) ;
  assign n8843 = ~n8761 & n8842 ;
  assign n8844 = n8837 ^ n8776 ^ n5964 ;
  assign n8845 = n8837 & n8844 ;
  assign n8846 = n8845 ^ n8649 ^ n8421 ;
  assign n8847 = n8837 ^ n8784 ^ n4346 ;
  assign n8848 = n8837 & n8847 ;
  assign n8849 = n8848 ^ n8672 ^ n8462 ;
  assign n8850 = n8837 ^ n8790 ^ n3464 ;
  assign n8851 = n8837 & n8850 ;
  assign n8852 = n8851 ^ n8675 ^ n8471 ;
  assign n8853 = n8837 ^ n8795 ^ n2839 ;
  assign n8854 = n8837 & n8853 ;
  assign n8855 = n8854 ^ n8652 ^ n8477 ;
  assign n8856 = n8837 ^ n8799 ^ n2269 ;
  assign n8857 = n8837 & n8856 ;
  assign n8858 = n8857 ^ n8662 ^ n8483 ;
  assign n8859 = n8837 ^ n8810 ^ n1118 ;
  assign n8860 = n8837 & n8859 ;
  assign n8861 = n8860 ^ n8726 ^ n8489 ;
  assign n8862 = n8837 ^ n8828 ^ n134 ;
  assign n8863 = n8837 & n8862 ;
  assign n8864 = n8863 ^ n8711 ^ n8406 ;
  assign n8865 = n8837 ^ n8767 ^ n7824 ;
  assign n8866 = n8837 & n8865 ;
  assign n8867 = n8866 ^ n8618 ^ n8498 ;
  assign n8868 = n8837 ^ n8777 ^ n5743 ;
  assign n8869 = n8837 & n8868 ;
  assign n8870 = n8869 ^ n8695 ^ n8412 ;
  assign n8871 = n8837 ^ n8779 ^ n5319 ;
  assign n8872 = n8837 & n8871 ;
  assign n8873 = n8872 ^ n8742 ^ n8382 ;
  assign n8874 = n8837 ^ n8785 ^ n4167 ;
  assign n8875 = n8837 & n8874 ;
  assign n8876 = n8875 ^ n8740 ^ n8465 ;
  assign n8877 = n8837 ^ n8794 ^ n2995 ;
  assign n8878 = n8837 & n8877 ;
  assign n8879 = n8878 ^ n8648 ^ n8341 ;
  assign n8880 = n8837 ^ n8796 ^ n2690 ;
  assign n8881 = n8837 & n8880 ;
  assign n8882 = n8881 ^ n8641 ^ n8437 ;
  assign n8883 = n8837 ^ n8797 ^ n2544 ;
  assign n8884 = n8837 & n8883 ;
  assign n8885 = n8884 ^ n8658 ^ n8480 ;
  assign n8886 = n8837 ^ n8802 ^ n2009 ;
  assign n8887 = n8837 & n8886 ;
  assign n8888 = n8887 ^ n8659 ^ n8346 ;
  assign n8889 = n8837 ^ n8803 ^ n1885 ;
  assign n8890 = n8837 & n8889 ;
  assign n8891 = n8890 ^ n8727 ^ n8349 ;
  assign n8892 = n8837 ^ n8813 ^ n859 ;
  assign n8893 = n8837 & n8892 ;
  assign n8894 = n8893 ^ n8686 ^ n8493 ;
  assign n8895 = n8837 ^ n8822 ^ n345 ;
  assign n8896 = n8837 & n8895 ;
  assign n8897 = n8896 ^ n8730 ^ n8388 ;
  assign n8898 = n8837 ^ n8825 ^ n217 ;
  assign n8899 = n8837 & n8898 ;
  assign n8900 = n8899 ^ n8734 ^ n8395 ;
  assign n8901 = n8837 ^ n8827 ^ n144 ;
  assign n8902 = n8837 & n8901 ;
  assign n8903 = n8902 ^ n8745 ^ n8403 ;
  assign n8904 = n8768 ^ n7575 ^ 1'b0 ;
  assign n8905 = n8837 & ~n8904 ;
  assign n8906 = n8905 ^ n8763 ^ n8510 ;
  assign n8907 = n8837 ^ n8770 ^ n7337 ;
  assign n8908 = n8837 & n8907 ;
  assign n8909 = n8908 ^ n8666 ^ n8503 ;
  assign n8910 = n8837 ^ n8773 ^ n6630 ;
  assign n8911 = n8837 & n8910 ;
  assign n8912 = n8911 ^ n8737 ^ n8459 ;
  assign n8913 = n8774 ^ n6401 ^ 1'b0 ;
  assign n8914 = n8837 & n8913 ;
  assign n8915 = n8914 ^ n8837 ^ n8607 ;
  assign n8916 = n8837 ^ n8778 ^ n5527 ;
  assign n8917 = n8837 & n8916 ;
  assign n8918 = n8917 ^ n8746 ^ n8335 ;
  assign n8919 = n8780 ^ n5124 ^ 1'b0 ;
  assign n8920 = n8837 & n8919 ;
  assign n8921 = n8920 ^ n8837 ^ n8611 ;
  assign n8922 = n8837 ^ n8781 ^ n4915 ;
  assign n8923 = n8837 & n8922 ;
  assign n8924 = n8923 ^ n8669 ^ n8367 ;
  assign n8925 = n8782 ^ n4728 ^ 1'b0 ;
  assign n8926 = n8837 & n8925 ;
  assign n8927 = n8926 ^ n8837 ^ n8612 ;
  assign n8928 = n8837 ^ n8783 ^ n4534 ;
  assign n8929 = n8837 & n8928 ;
  assign n8930 = n8929 ^ n8646 ^ n8338 ;
  assign n8931 = n8837 ^ n8786 ^ n3986 ;
  assign n8932 = n8837 & n8931 ;
  assign n8933 = n8932 ^ n8635 ^ n8430 ;
  assign n8934 = n8837 ^ n8793 ^ n3141 ;
  assign n8935 = n8837 & n8934 ;
  assign n8936 = n8935 ^ n8656 ^ n8474 ;
  assign n8937 = n8800 ^ n2139 ^ 1'b0 ;
  assign n8938 = n8837 & n8937 ;
  assign n8939 = n8938 ^ n8837 ^ n8598 ;
  assign n8940 = n8837 ^ n8804 ^ n1766 ;
  assign n8941 = n8837 & n8940 ;
  assign n8942 = n8941 ^ n8678 ^ n8445 ;
  assign n8943 = n8837 ^ n8805 ^ n1652 ;
  assign n8944 = n8837 & n8943 ;
  assign n8945 = n8944 ^ n8680 ^ n8370 ;
  assign n8946 = n8837 ^ n8806 ^ n1534 ;
  assign n8947 = n8837 & n8946 ;
  assign n8948 = n8947 ^ n8637 ^ n8373 ;
  assign n8949 = n8809 ^ n1220 ^ 1'b0 ;
  assign n8950 = n8837 & n8949 ;
  assign n8951 = n8950 ^ n8837 ^ n8592 ;
  assign n8952 = n8837 ^ n8811 ^ n1034 ;
  assign n8953 = n8837 & n8952 ;
  assign n8954 = n8953 ^ n8639 ^ n8352 ;
  assign n8955 = n8837 ^ n8812 ^ n941 ;
  assign n8956 = n8837 & n8955 ;
  assign n8957 = n8956 ^ n8644 ^ n8491 ;
  assign n8958 = n8837 ^ n8814 ^ n785 ;
  assign n8959 = n8837 & n8958 ;
  assign n8960 = n8959 ^ n8654 ^ n8376 ;
  assign n8961 = n8837 ^ n8816 ^ n640 ;
  assign n8962 = n8837 & n8961 ;
  assign n8963 = n8962 ^ n8728 ^ n8384 ;
  assign n8964 = n8818 ^ n572 ^ 1'b0 ;
  assign n8965 = n8837 & n8964 ;
  assign n8966 = n8965 ^ n8837 ^ n8693 ;
  assign n8967 = n8837 ^ n8821 ^ n399 ;
  assign n8968 = n8837 & n8967 ;
  assign n8969 = n8968 ^ n8702 ^ n8360 ;
  assign n8970 = n8837 ^ n8823 ^ n302 ;
  assign n8971 = n8837 & n8970 ;
  assign n8972 = n8971 ^ n8643 ^ n8397 ;
  assign n8973 = ( n8829 & n8832 ) | ( n8829 & ~n8837 ) | ( n8832 & ~n8837 ) ;
  assign n8974 = n8792 ^ n3302 ^ 1'b0 ;
  assign n8975 = n8837 & n8974 ;
  assign n8976 = n8807 ^ n1416 ^ 1'b0 ;
  assign n8977 = n8975 ^ n8837 ^ n8613 ;
  assign n8978 = ~n8614 & n8829 ;
  assign n8979 = n8815 ^ n716 ^ 1'b0 ;
  assign n8980 = n8772 ^ n6858 ^ 1'b0 ;
  assign n8981 = n8837 ^ n8771 ^ n7089 ;
  assign n8982 = n8798 ^ n2404 ^ 1'b0 ;
  assign n8983 = n8837 & n8982 ;
  assign n8984 = n8837 & n8980 ;
  assign n8985 = n8837 ^ n8819 ^ n514 ;
  assign n8986 = n8983 ^ n8837 ^ n8596 ;
  assign n8987 = n8837 & n8976 ;
  assign n8988 = n8984 ^ n8837 ^ n8602 ;
  assign n8989 = n8837 ^ n8787 ^ n3804 ;
  assign n8990 = n8837 & n8989 ;
  assign n8991 = ( ~x50 & x61 ) | ( ~x50 & x72 ) | ( x61 & x72 ) ;
  assign n8992 = x50 | n8991 ;
  assign n8993 = x72 & n8837 ;
  assign n8994 = n8837 ^ n8808 ^ n1318 ;
  assign n8995 = n8837 & n8994 ;
  assign n8996 = n8837 ^ n8820 ^ n458 ;
  assign n8997 = n8995 ^ n8683 ^ n8486 ;
  assign n8998 = ( n8587 & ~n8992 ) | ( n8587 & n8993 ) | ( ~n8992 & n8993 ) ;
  assign n8999 = n8990 ^ n8735 ^ n8468 ;
  assign n9000 = ( ~n8587 & n8992 ) | ( ~n8587 & n8993 ) | ( n8992 & n8993 ) ;
  assign n9001 = n8824 ^ n261 ^ 1'b0 ;
  assign n9002 = n8837 & n9001 ;
  assign n9003 = ( ~n8614 & n8829 ) | ( ~n8614 & n8837 ) | ( n8829 & n8837 ) ;
  assign n9004 = ( n8864 & ~n8978 ) | ( n8864 & n9003 ) | ( ~n8978 & n9003 ) ;
  assign n9005 = ( n136 & n8614 ) | ( n136 & n8829 ) | ( n8614 & n8829 ) ;
  assign n9006 = n8826 ^ n179 ^ 1'b0 ;
  assign n9007 = n8789 ^ n3631 ^ 1'b0 ;
  assign n9008 = ~n8993 & n9000 ;
  assign n9009 = ~n8973 & n9005 ;
  assign n9010 = n8843 ^ n8751 ^ x105 ;
  assign n9011 = n8837 & n9006 ;
  assign n9012 = n8837 ^ n8775 ^ n6171 ;
  assign n9013 = n8837 & n9012 ;
  assign n9014 = n8837 ^ n8766 ^ n8069 ;
  assign n9015 = n8837 & n9007 ;
  assign n9016 = n9015 ^ n8837 ^ n8619 ;
  assign n9017 = n8993 ^ n8837 ^ x83 ;
  assign n9018 = n8837 & n8996 ;
  assign n9019 = n8837 & n8981 ;
  assign n9020 = n9018 ^ n8698 ^ n8455 ;
  assign n9021 = n8837 & n8979 ;
  assign n9022 = n9019 ^ n8748 ^ n8502 ;
  assign n9023 = n9002 ^ n8837 ^ n8706 ;
  assign n9024 = n9013 ^ n8615 ^ n8418 ;
  assign n9025 = n9011 ^ n8837 ^ n8709 ;
  assign n9026 = n8837 & n8985 ;
  assign n9027 = n8837 & n9014 ;
  assign n9028 = n8987 ^ n8837 ^ n8595 ;
  assign n9029 = n9021 ^ n8837 ^ n8690 ;
  assign n9030 = n9026 ^ n8732 ^ n8357 ;
  assign n9031 = n9027 ^ n8617 ^ x116 ;
  assign n9032 = n8841 ^ x94 ^ 1'b0 ;
  assign n9033 = n9008 | n9017 ;
  assign n9034 = ~n8998 & n9033 ;
  assign n9035 = ( ~n8324 & n9032 ) | ( ~n8324 & n9034 ) | ( n9032 & n9034 ) ;
  assign n9036 = ( ~n8069 & n9010 ) | ( ~n8069 & n9035 ) | ( n9010 & n9035 ) ;
  assign n9037 = ( ~n7824 & n9031 ) | ( ~n7824 & n9036 ) | ( n9031 & n9036 ) ;
  assign n9038 = ( ~n7575 & n8867 ) | ( ~n7575 & n9037 ) | ( n8867 & n9037 ) ;
  assign n9039 = ( ~n7337 & n8906 ) | ( ~n7337 & n9038 ) | ( n8906 & n9038 ) ;
  assign n9040 = ( ~n7089 & n8909 ) | ( ~n7089 & n9039 ) | ( n8909 & n9039 ) ;
  assign n9041 = ( ~n6858 & n9022 ) | ( ~n6858 & n9040 ) | ( n9022 & n9040 ) ;
  assign n9042 = ( ~n6630 & n8988 ) | ( ~n6630 & n9041 ) | ( n8988 & n9041 ) ;
  assign n9043 = ( ~n6401 & n8912 ) | ( ~n6401 & n9042 ) | ( n8912 & n9042 ) ;
  assign n9044 = ( ~n6171 & n8915 ) | ( ~n6171 & n9043 ) | ( n8915 & n9043 ) ;
  assign n9045 = ( ~n5964 & n9024 ) | ( ~n5964 & n9044 ) | ( n9024 & n9044 ) ;
  assign n9046 = ( ~n5743 & n8846 ) | ( ~n5743 & n9045 ) | ( n8846 & n9045 ) ;
  assign n9047 = ( ~n5527 & n8870 ) | ( ~n5527 & n9046 ) | ( n8870 & n9046 ) ;
  assign n9048 = ( ~n5319 & n8918 ) | ( ~n5319 & n9047 ) | ( n8918 & n9047 ) ;
  assign n9049 = ( ~n5124 & n8873 ) | ( ~n5124 & n9048 ) | ( n8873 & n9048 ) ;
  assign n9050 = ( ~n4915 & n8921 ) | ( ~n4915 & n9049 ) | ( n8921 & n9049 ) ;
  assign n9051 = ( ~n4728 & n8924 ) | ( ~n4728 & n9050 ) | ( n8924 & n9050 ) ;
  assign n9052 = ( ~n4534 & n8927 ) | ( ~n4534 & n9051 ) | ( n8927 & n9051 ) ;
  assign n9053 = ( ~n4346 & n8930 ) | ( ~n4346 & n9052 ) | ( n8930 & n9052 ) ;
  assign n9054 = ( ~n4167 & n8849 ) | ( ~n4167 & n9053 ) | ( n8849 & n9053 ) ;
  assign n9055 = ( ~n3986 & n8876 ) | ( ~n3986 & n9054 ) | ( n8876 & n9054 ) ;
  assign n9056 = ( ~n3804 & n8933 ) | ( ~n3804 & n9055 ) | ( n8933 & n9055 ) ;
  assign n9057 = ( ~n3631 & n8999 ) | ( ~n3631 & n9056 ) | ( n8999 & n9056 ) ;
  assign n9058 = ( ~n3464 & n9016 ) | ( ~n3464 & n9057 ) | ( n9016 & n9057 ) ;
  assign n9059 = ( ~n3302 & n8852 ) | ( ~n3302 & n9058 ) | ( n8852 & n9058 ) ;
  assign n9060 = ( ~n3141 & n8977 ) | ( ~n3141 & n9059 ) | ( n8977 & n9059 ) ;
  assign n9061 = ( ~n2995 & n8936 ) | ( ~n2995 & n9060 ) | ( n8936 & n9060 ) ;
  assign n9062 = ( ~n2839 & n8879 ) | ( ~n2839 & n9061 ) | ( n8879 & n9061 ) ;
  assign n9063 = ( ~n2690 & n8855 ) | ( ~n2690 & n9062 ) | ( n8855 & n9062 ) ;
  assign n9064 = ( ~n2544 & n8882 ) | ( ~n2544 & n9063 ) | ( n8882 & n9063 ) ;
  assign n9065 = ( ~n2404 & n8885 ) | ( ~n2404 & n9064 ) | ( n8885 & n9064 ) ;
  assign n9066 = ( ~n2269 & n8986 ) | ( ~n2269 & n9065 ) | ( n8986 & n9065 ) ;
  assign n9067 = ( ~n2139 & n8858 ) | ( ~n2139 & n9066 ) | ( n8858 & n9066 ) ;
  assign n9068 = ( ~n2009 & n8939 ) | ( ~n2009 & n9067 ) | ( n8939 & n9067 ) ;
  assign n9069 = ( ~n1885 & n8888 ) | ( ~n1885 & n9068 ) | ( n8888 & n9068 ) ;
  assign n9070 = ( ~n1766 & n8891 ) | ( ~n1766 & n9069 ) | ( n8891 & n9069 ) ;
  assign n9071 = ( ~n1652 & n8942 ) | ( ~n1652 & n9070 ) | ( n8942 & n9070 ) ;
  assign n9072 = ( ~n1534 & n8945 ) | ( ~n1534 & n9071 ) | ( n8945 & n9071 ) ;
  assign n9073 = ( ~n1416 & n8948 ) | ( ~n1416 & n9072 ) | ( n8948 & n9072 ) ;
  assign n9074 = ( ~n1318 & n9028 ) | ( ~n1318 & n9073 ) | ( n9028 & n9073 ) ;
  assign n9075 = ( ~n1220 & n8997 ) | ( ~n1220 & n9074 ) | ( n8997 & n9074 ) ;
  assign n9076 = ( ~n1118 & n8951 ) | ( ~n1118 & n9075 ) | ( n8951 & n9075 ) ;
  assign n9077 = ( ~n1034 & n8861 ) | ( ~n1034 & n9076 ) | ( n8861 & n9076 ) ;
  assign n9078 = ( ~n941 & n8954 ) | ( ~n941 & n9077 ) | ( n8954 & n9077 ) ;
  assign n9079 = ( ~n859 & n8957 ) | ( ~n859 & n9078 ) | ( n8957 & n9078 ) ;
  assign n9080 = ( ~n785 & n8894 ) | ( ~n785 & n9079 ) | ( n8894 & n9079 ) ;
  assign n9081 = ( ~n716 & n8960 ) | ( ~n716 & n9080 ) | ( n8960 & n9080 ) ;
  assign n9082 = ( ~n640 & n9029 ) | ( ~n640 & n9081 ) | ( n9029 & n9081 ) ;
  assign n9083 = ( ~n572 & n8963 ) | ( ~n572 & n9082 ) | ( n8963 & n9082 ) ;
  assign n9084 = ( ~n514 & n8966 ) | ( ~n514 & n9083 ) | ( n8966 & n9083 ) ;
  assign n9085 = ( ~n458 & n9030 ) | ( ~n458 & n9084 ) | ( n9030 & n9084 ) ;
  assign n9086 = ( ~n399 & n9020 ) | ( ~n399 & n9085 ) | ( n9020 & n9085 ) ;
  assign n9087 = ( ~n345 & n8969 ) | ( ~n345 & n9086 ) | ( n8969 & n9086 ) ;
  assign n9088 = ( ~n302 & n8897 ) | ( ~n302 & n9087 ) | ( n8897 & n9087 ) ;
  assign n9089 = ( ~n261 & n8972 ) | ( ~n261 & n9088 ) | ( n8972 & n9088 ) ;
  assign n9090 = ( ~n217 & n9023 ) | ( ~n217 & n9089 ) | ( n9023 & n9089 ) ;
  assign n9091 = ( ~n179 & n8900 ) | ( ~n179 & n9090 ) | ( n8900 & n9090 ) ;
  assign n9092 = ( ~n144 & n9025 ) | ( ~n144 & n9091 ) | ( n9025 & n9091 ) ;
  assign n9093 = ( ~n134 & n8903 ) | ( ~n134 & n9092 ) | ( n8903 & n9092 ) ;
  assign n9094 = ( ~x30 & n9004 ) | ( ~x30 & n9093 ) | ( n9004 & n9093 ) ;
  assign n9095 = ~n136 & n9094 ;
  assign n9096 = n8864 & n9093 ;
  assign n9097 = n9009 | n9096 ;
  assign n9098 = n9095 | n9097 ;
  assign n9099 = n9098 ^ n9085 ^ n399 ;
  assign n9100 = n9098 & n9099 ;
  assign n9101 = n9100 ^ n9018 ^ n8700 ;
  assign n9102 = n9098 ^ n9071 ^ n1534 ;
  assign n9103 = n9098 & n9102 ;
  assign n9104 = n9103 ^ n8944 ^ n8681 ;
  assign n9105 = n9098 ^ n9063 ^ n2544 ;
  assign n9106 = n9098 & n9105 ;
  assign n9107 = n9106 ^ n8881 ^ n8642 ;
  assign n9108 = n9098 ^ n9062 ^ n2690 ;
  assign n9109 = n9098 & n9108 ;
  assign n9110 = n9109 ^ n8854 ^ n8653 ;
  assign n9111 = n9098 ^ n9061 ^ n2839 ;
  assign n9112 = n9098 & n9111 ;
  assign n9113 = n9112 ^ n8878 ^ n8664 ;
  assign n9114 = n9098 ^ n9058 ^ n3302 ;
  assign n9115 = n9098 & n9114 ;
  assign n9116 = n9115 ^ n8851 ^ n8676 ;
  assign n9117 = n9098 ^ n9054 ^ n3986 ;
  assign n9118 = n9098 & n9117 ;
  assign n9119 = n9118 ^ n8875 ^ n8741 ;
  assign n9120 = n9098 ^ n9053 ^ n4167 ;
  assign n9121 = n9098 & n9120 ;
  assign n9122 = n9121 ^ n8848 ^ n8673 ;
  assign n9123 = n9098 ^ n9045 ^ n5743 ;
  assign n9124 = n9098 & n9123 ;
  assign n9125 = n9124 ^ n8845 ^ n8651 ;
  assign n9126 = n9098 ^ n9036 ^ n7824 ;
  assign n9127 = n9098 & n9126 ;
  assign n9128 = n9127 ^ n9027 ^ n8753 ;
  assign n9129 = n9008 & n9098 ;
  assign n9130 = ( n8998 & n9098 ) | ( n8998 & ~n9129 ) | ( n9098 & ~n9129 ) ;
  assign n9131 = n9130 ^ n9017 ^ n8998 ;
  assign n9132 = n9098 ^ n9090 ^ n179 ;
  assign n9133 = n9098 & n9132 ;
  assign n9134 = n9133 ^ n8899 ^ n8744 ;
  assign n9135 = n9098 ^ n9088 ^ n261 ;
  assign n9136 = n9098 & n9135 ;
  assign n9137 = n9136 ^ n8971 ^ n8650 ;
  assign n9138 = n9098 ^ n9086 ^ n345 ;
  assign n9139 = n9098 & n9138 ;
  assign n9140 = n9139 ^ n8968 ^ n8703 ;
  assign n9141 = n9098 ^ n9080 ^ n716 ;
  assign n9142 = n9098 & n9141 ;
  assign n9143 = n9142 ^ n8959 ^ n8655 ;
  assign n9144 = n9098 ^ n9079 ^ n785 ;
  assign n9145 = n9098 & n9144 ;
  assign n9146 = n9145 ^ n8893 ^ n8687 ;
  assign n9147 = n9098 ^ n9076 ^ n1034 ;
  assign n9148 = n9098 & n9147 ;
  assign n9149 = n9148 ^ n8860 ^ n8791 ;
  assign n9150 = n9098 ^ n9069 ^ n1766 ;
  assign n9151 = n9098 & n9150 ;
  assign n9152 = n9151 ^ n8890 ^ n8736 ;
  assign n9153 = n9098 ^ n9068 ^ n1885 ;
  assign n9154 = n9098 & n9153 ;
  assign n9155 = n9154 ^ n8887 ^ n8660 ;
  assign n9156 = n9098 ^ n9066 ^ n2139 ;
  assign n9157 = n9098 & n9156 ;
  assign n9158 = n9157 ^ n8857 ^ n8663 ;
  assign n9159 = n9098 ^ n9052 ^ n4346 ;
  assign n9160 = n9098 & n9159 ;
  assign n9161 = n9160 ^ n8929 ^ n8647 ;
  assign n9162 = n9098 ^ n9042 ^ n6401 ;
  assign n9163 = n9098 & n9162 ;
  assign n9164 = n9163 ^ n8911 ^ n8738 ;
  assign n9165 = n9098 ^ n9039 ^ n7089 ;
  assign n9166 = n9098 & n9165 ;
  assign n9167 = n9166 ^ n8908 ^ n8667 ;
  assign n9168 = n9098 ^ n9038 ^ n7337 ;
  assign n9169 = n9098 & n9168 ;
  assign n9170 = n9169 ^ n8905 ^ n8769 ;
  assign n9171 = n9098 ^ n9037 ^ n7575 ;
  assign n9172 = n9098 & n9171 ;
  assign n9173 = n9172 ^ n8866 ^ n8764 ;
  assign n9174 = n9098 ^ n9035 ^ n8069 ;
  assign n9175 = n9098 & n9174 ;
  assign n9176 = n9175 ^ n8843 ^ n8752 ;
  assign n9177 = n9092 ^ n134 ^ 1'b0 ;
  assign n9178 = n9098 & ~n9177 ;
  assign n9179 = n9178 ^ n8902 ^ n8747 ;
  assign n9180 = n9098 ^ n9087 ^ n302 ;
  assign n9181 = n9098 & n9180 ;
  assign n9182 = n9181 ^ n8896 ^ n8731 ;
  assign n9183 = n9098 ^ n9084 ^ n458 ;
  assign n9184 = n9098 & n9183 ;
  assign n9185 = n9184 ^ n9026 ^ n8733 ;
  assign n9186 = n9098 ^ n9082 ^ n572 ;
  assign n9187 = n9098 & n9186 ;
  assign n9188 = n9187 ^ n8962 ^ n8729 ;
  assign n9189 = n9098 ^ n9078 ^ n859 ;
  assign n9190 = n9098 & n9189 ;
  assign n9191 = n9190 ^ n8956 ^ n8645 ;
  assign n9192 = n9098 ^ n9077 ^ n941 ;
  assign n9193 = n9098 & n9192 ;
  assign n9194 = n9193 ^ n8953 ^ n8640 ;
  assign n9195 = n9098 ^ n9074 ^ n1220 ;
  assign n9196 = n9098 & n9195 ;
  assign n9197 = n9196 ^ n8995 ^ n8684 ;
  assign n9198 = n9098 ^ n9072 ^ n1416 ;
  assign n9199 = n9098 & n9198 ;
  assign n9200 = n9199 ^ n8947 ^ n8638 ;
  assign n9201 = n9098 ^ n9070 ^ n1652 ;
  assign n9202 = n9098 & n9201 ;
  assign n9203 = n9202 ^ n8941 ^ n8699 ;
  assign n9204 = n9098 ^ n9064 ^ n2404 ;
  assign n9205 = n9098 & n9204 ;
  assign n9206 = n9205 ^ n8884 ^ n8661 ;
  assign n9207 = n9098 ^ n9055 ^ n3804 ;
  assign n9208 = n9098 & n9207 ;
  assign n9209 = n9208 ^ n8932 ^ n8636 ;
  assign n9210 = n9098 ^ n9048 ^ n5124 ;
  assign n9211 = n9098 & n9210 ;
  assign n9212 = n9211 ^ n8872 ^ n8743 ;
  assign n9213 = n9098 ^ n9047 ^ n5319 ;
  assign n9214 = n9098 & n9213 ;
  assign n9215 = n9214 ^ n8917 ^ n8750 ;
  assign n9216 = n9098 ^ n9060 ^ n2995 ;
  assign n9217 = n9098 & n9216 ;
  assign n9218 = n9217 ^ n8935 ^ n8657 ;
  assign n9219 = n9098 ^ n9056 ^ n3631 ;
  assign n9220 = n9098 & n9219 ;
  assign n9221 = n9220 ^ n8990 ^ n8739 ;
  assign n9222 = n9098 ^ n9050 ^ n4728 ;
  assign n9223 = n9098 ^ n9046 ^ n5527 ;
  assign n9224 = n9098 & n9223 ;
  assign n9225 = n9224 ^ n8869 ^ n8696 ;
  assign n9226 = n9098 ^ n9044 ^ n5964 ;
  assign n9227 = n9098 & n9226 ;
  assign n9228 = n9227 ^ n9013 ^ n8616 ;
  assign n9229 = n9098 ^ n9040 ^ n6858 ;
  assign n9230 = n9098 ^ n9034 ^ n8324 ;
  assign n9231 = n9098 & n9230 ;
  assign n9232 = n9231 ^ n8841 ^ x94 ;
  assign n9233 = x50 | n9098 ;
  assign n9234 = n9233 ^ x61 ^ x50 ;
  assign n9235 = ( x50 & n9095 ) | ( x50 & n9096 ) | ( n9095 & n9096 ) ;
  assign n9236 = ( x50 & n9009 ) | ( x50 & n9235 ) | ( n9009 & n9235 ) ;
  assign n9237 = ( ~x0 & x39 ) | ( ~x0 & x50 ) | ( x39 & x50 ) ;
  assign n9238 = x0 | n9237 ;
  assign n9239 = ~x50 & n9238 ;
  assign n9240 = ( ~n9236 & n9238 ) | ( ~n9236 & n9239 ) | ( n9238 & n9239 ) ;
  assign n9241 = ( ~n8837 & n9234 ) | ( ~n8837 & n9240 ) | ( n9234 & n9240 ) ;
  assign n9242 = ( n8837 & ~n9095 ) | ( n8837 & n9096 ) | ( ~n9095 & n9096 ) ;
  assign n9243 = ~n9097 & n9242 ;
  assign n9244 = x50 & ~x61 ;
  assign n9245 = ( ~x61 & n9098 ) | ( ~x61 & n9244 ) | ( n9098 & n9244 ) ;
  assign n9246 = ( n9243 & ~n9244 ) | ( n9243 & n9245 ) | ( ~n9244 & n9245 ) ;
  assign n9247 = n9246 ^ x72 ^ 1'b0 ;
  assign n9248 = ( ~n8587 & n9241 ) | ( ~n8587 & n9247 ) | ( n9241 & n9247 ) ;
  assign n9249 = ( ~n8324 & n9131 ) | ( ~n8324 & n9248 ) | ( n9131 & n9248 ) ;
  assign n9250 = n9098 & n9229 ;
  assign n9251 = n9250 ^ n9019 ^ n8749 ;
  assign n9252 = ( ~n8069 & n9232 ) | ( ~n8069 & n9249 ) | ( n9232 & n9249 ) ;
  assign n9253 = ( ~n7824 & n9176 ) | ( ~n7824 & n9252 ) | ( n9176 & n9252 ) ;
  assign n9254 = ( ~n7575 & n9128 ) | ( ~n7575 & n9253 ) | ( n9128 & n9253 ) ;
  assign n9255 = n9098 & n9222 ;
  assign n9256 = n9255 ^ n8923 ^ n8670 ;
  assign n9257 = ( ~n7337 & n9173 ) | ( ~n7337 & n9254 ) | ( n9173 & n9254 ) ;
  assign n9258 = ( ~n7089 & n9170 ) | ( ~n7089 & n9257 ) | ( n9170 & n9257 ) ;
  assign n9259 = ( ~n6858 & n9167 ) | ( ~n6858 & n9258 ) | ( n9167 & n9258 ) ;
  assign n9260 = ( ~n6630 & n9251 ) | ( ~n6630 & n9259 ) | ( n9251 & n9259 ) ;
  assign n9261 = n9059 ^ n3141 ^ 1'b0 ;
  assign n9262 = n9098 & n9261 ;
  assign n9263 = n9262 ^ n9098 ^ n8977 ;
  assign n9264 = n9057 ^ n3464 ^ 1'b0 ;
  assign n9265 = n9098 & n9264 ;
  assign n9266 = n9265 ^ n9098 ^ n9016 ;
  assign n9267 = n9051 ^ n4534 ^ 1'b0 ;
  assign n9268 = n9098 & n9267 ;
  assign n9269 = n9268 ^ n9098 ^ n8927 ;
  assign n9270 = n9049 ^ n4915 ^ 1'b0 ;
  assign n9271 = n9098 & n9270 ;
  assign n9272 = n9271 ^ n9098 ^ n8921 ;
  assign n9273 = n9043 ^ n6171 ^ 1'b0 ;
  assign n9274 = n9098 & n9273 ;
  assign n9275 = n9274 ^ n9098 ^ n8915 ;
  assign n9276 = n9041 ^ n6630 ^ 1'b0 ;
  assign n9277 = n9098 & n9276 ;
  assign n9278 = n9277 ^ n9098 ^ n8988 ;
  assign n9279 = ( ~n6401 & n9260 ) | ( ~n6401 & n9278 ) | ( n9260 & n9278 ) ;
  assign n9280 = ( ~n6171 & n9164 ) | ( ~n6171 & n9279 ) | ( n9164 & n9279 ) ;
  assign n9281 = ( ~n5964 & n9275 ) | ( ~n5964 & n9280 ) | ( n9275 & n9280 ) ;
  assign n9282 = ( ~n5743 & n9228 ) | ( ~n5743 & n9281 ) | ( n9228 & n9281 ) ;
  assign n9283 = ( ~n5527 & n9125 ) | ( ~n5527 & n9282 ) | ( n9125 & n9282 ) ;
  assign n9284 = ( ~n5319 & n9225 ) | ( ~n5319 & n9283 ) | ( n9225 & n9283 ) ;
  assign n9285 = ( ~n5124 & n9215 ) | ( ~n5124 & n9284 ) | ( n9215 & n9284 ) ;
  assign n9286 = ( ~n4915 & n9212 ) | ( ~n4915 & n9285 ) | ( n9212 & n9285 ) ;
  assign n9287 = ( ~n4728 & n9272 ) | ( ~n4728 & n9286 ) | ( n9272 & n9286 ) ;
  assign n9288 = ( ~n4534 & n9256 ) | ( ~n4534 & n9287 ) | ( n9256 & n9287 ) ;
  assign n9289 = ( ~n4346 & n9269 ) | ( ~n4346 & n9288 ) | ( n9269 & n9288 ) ;
  assign n9290 = ( ~n4167 & n9161 ) | ( ~n4167 & n9289 ) | ( n9161 & n9289 ) ;
  assign n9291 = ( ~n3986 & n9122 ) | ( ~n3986 & n9290 ) | ( n9122 & n9290 ) ;
  assign n9292 = ( ~n3804 & n9119 ) | ( ~n3804 & n9291 ) | ( n9119 & n9291 ) ;
  assign n9293 = ( ~n3631 & n9209 ) | ( ~n3631 & n9292 ) | ( n9209 & n9292 ) ;
  assign n9294 = ( ~n3464 & n9221 ) | ( ~n3464 & n9293 ) | ( n9221 & n9293 ) ;
  assign n9295 = ( ~n3302 & n9266 ) | ( ~n3302 & n9294 ) | ( n9266 & n9294 ) ;
  assign n9296 = ( ~n3141 & n9116 ) | ( ~n3141 & n9295 ) | ( n9116 & n9295 ) ;
  assign n9297 = ( ~n2995 & n9263 ) | ( ~n2995 & n9296 ) | ( n9263 & n9296 ) ;
  assign n9298 = ( ~n2839 & n9218 ) | ( ~n2839 & n9297 ) | ( n9218 & n9297 ) ;
  assign n9299 = ( ~n2690 & n9113 ) | ( ~n2690 & n9298 ) | ( n9113 & n9298 ) ;
  assign n9300 = ( ~n2544 & n9110 ) | ( ~n2544 & n9299 ) | ( n9110 & n9299 ) ;
  assign n9301 = n9089 ^ n217 ^ 1'b0 ;
  assign n9302 = n9098 & n9301 ;
  assign n9303 = n9302 ^ n9098 ^ n9023 ;
  assign n9304 = n9091 ^ n144 ^ 1'b0 ;
  assign n9305 = n9098 & n9304 ;
  assign n9306 = n9305 ^ n9098 ^ n9025 ;
  assign n9307 = n9065 ^ n2269 ^ 1'b0 ;
  assign n9308 = n9098 & n9307 ;
  assign n9309 = n9308 ^ n9098 ^ n8986 ;
  assign n9310 = ( ~n2404 & n9107 ) | ( ~n2404 & n9300 ) | ( n9107 & n9300 ) ;
  assign n9311 = n9083 ^ n514 ^ 1'b0 ;
  assign n9312 = n9098 & n9311 ;
  assign n9313 = n9312 ^ n9098 ^ n8966 ;
  assign n9314 = n9081 ^ n640 ^ 1'b0 ;
  assign n9315 = n9098 & n9314 ;
  assign n9316 = n9315 ^ n9098 ^ n9029 ;
  assign n9317 = n9075 ^ n1118 ^ 1'b0 ;
  assign n9318 = n9098 & n9317 ;
  assign n9319 = n9318 ^ n9098 ^ n8951 ;
  assign n9320 = n9073 ^ n1318 ^ 1'b0 ;
  assign n9321 = n9098 & n9320 ;
  assign n9322 = n9321 ^ n9098 ^ n9028 ;
  assign n9323 = n9067 ^ n2009 ^ 1'b0 ;
  assign n9324 = n9098 & n9323 ;
  assign n9325 = n9324 ^ n9098 ^ n8939 ;
  assign n9326 = ( ~n2269 & n9206 ) | ( ~n2269 & n9310 ) | ( n9206 & n9310 ) ;
  assign n9327 = ( ~n2139 & n9309 ) | ( ~n2139 & n9326 ) | ( n9309 & n9326 ) ;
  assign n9328 = ( ~n2009 & n9158 ) | ( ~n2009 & n9327 ) | ( n9158 & n9327 ) ;
  assign n9329 = ( ~n1885 & n9325 ) | ( ~n1885 & n9328 ) | ( n9325 & n9328 ) ;
  assign n9330 = ( n136 & n8864 ) | ( n136 & n9093 ) | ( n8864 & n9093 ) ;
  assign n9331 = ( n136 & n9093 ) | ( n136 & n9096 ) | ( n9093 & n9096 ) ;
  assign n9332 = ( ~n1766 & n9155 ) | ( ~n1766 & n9329 ) | ( n9155 & n9329 ) ;
  assign n9333 = ( ~n1652 & n9152 ) | ( ~n1652 & n9332 ) | ( n9152 & n9332 ) ;
  assign n9334 = ( ~n1534 & n9203 ) | ( ~n1534 & n9333 ) | ( n9203 & n9333 ) ;
  assign n9335 = ( ~n1416 & n9104 ) | ( ~n1416 & n9334 ) | ( n9104 & n9334 ) ;
  assign n9336 = ( ~n1318 & n9200 ) | ( ~n1318 & n9335 ) | ( n9200 & n9335 ) ;
  assign n9337 = ( ~n1220 & n9322 ) | ( ~n1220 & n9336 ) | ( n9322 & n9336 ) ;
  assign n9338 = ( ~n1118 & n9197 ) | ( ~n1118 & n9337 ) | ( n9197 & n9337 ) ;
  assign n9339 = ( ~n1034 & n9319 ) | ( ~n1034 & n9338 ) | ( n9319 & n9338 ) ;
  assign n9340 = ( ~n941 & n9149 ) | ( ~n941 & n9339 ) | ( n9149 & n9339 ) ;
  assign n9341 = ( ~n859 & n9194 ) | ( ~n859 & n9340 ) | ( n9194 & n9340 ) ;
  assign n9342 = ( ~n785 & n9191 ) | ( ~n785 & n9341 ) | ( n9191 & n9341 ) ;
  assign n9343 = ( ~n716 & n9146 ) | ( ~n716 & n9342 ) | ( n9146 & n9342 ) ;
  assign n9344 = ( ~n640 & n9143 ) | ( ~n640 & n9343 ) | ( n9143 & n9343 ) ;
  assign n9345 = ( ~n572 & n9316 ) | ( ~n572 & n9344 ) | ( n9316 & n9344 ) ;
  assign n9346 = ( ~n514 & n9188 ) | ( ~n514 & n9345 ) | ( n9188 & n9345 ) ;
  assign n9347 = ( ~n458 & n9313 ) | ( ~n458 & n9346 ) | ( n9313 & n9346 ) ;
  assign n9348 = ( n9096 & ~n9098 ) | ( n9096 & n9331 ) | ( ~n9098 & n9331 ) ;
  assign n9349 = ( ~n399 & n9185 ) | ( ~n399 & n9347 ) | ( n9185 & n9347 ) ;
  assign n9350 = ( ~n345 & n9101 ) | ( ~n345 & n9349 ) | ( n9101 & n9349 ) ;
  assign n9351 = ( ~n302 & n9140 ) | ( ~n302 & n9350 ) | ( n9140 & n9350 ) ;
  assign n9352 = ( ~n261 & n9182 ) | ( ~n261 & n9351 ) | ( n9182 & n9351 ) ;
  assign n9353 = ( ~n217 & n9137 ) | ( ~n217 & n9352 ) | ( n9137 & n9352 ) ;
  assign n9354 = ( ~n179 & n9303 ) | ( ~n179 & n9353 ) | ( n9303 & n9353 ) ;
  assign n9355 = ( ~n144 & n9134 ) | ( ~n144 & n9354 ) | ( n9134 & n9354 ) ;
  assign n9356 = ( ~n134 & n9306 ) | ( ~n134 & n9355 ) | ( n9306 & n9355 ) ;
  assign n9357 = n9306 & n9355 ;
  assign n9358 = ~n134 & n9356 ;
  assign n9359 = ( ~n9093 & n9096 ) | ( ~n9093 & n9098 ) | ( n9096 & n9098 ) ;
  assign n9360 = n9179 & ~n9356 ;
  assign n9361 = ( ~n8864 & n9096 ) | ( ~n8864 & n9359 ) | ( n9096 & n9359 ) ;
  assign n9362 = ( ~n9179 & n9358 ) | ( ~n9179 & n9361 ) | ( n9358 & n9361 ) ;
  assign n9363 = n9179 & ~n9362 ;
  assign n9364 = ( ~n9357 & n9362 ) | ( ~n9357 & n9363 ) | ( n9362 & n9363 ) ;
  assign n9365 = ( ~n136 & n9357 ) | ( ~n136 & n9364 ) | ( n9357 & n9364 ) ;
  assign n9366 = ( n9179 & ~n9360 ) | ( n9179 & n9365 ) | ( ~n9360 & n9365 ) ;
  assign n9367 = n9366 ^ n9348 ^ n9330 ;
  assign n9368 = n9366 | n9367 ;
  assign y0 = n9368 ;
  assign y1 = n6858 ;
  assign y2 = n6630 ;
  assign y3 = n6401 ;
  assign y4 = n6171 ;
  assign y5 = n5964 ;
  assign y6 = n5743 ;
  assign y7 = n5527 ;
  assign y8 = n5319 ;
  assign y9 = n5124 ;
  assign y10 = n4915 ;
  assign y11 = n9098 ;
  assign y12 = n4728 ;
  assign y13 = n4534 ;
  assign y14 = n4346 ;
  assign y15 = n4167 ;
  assign y16 = n3986 ;
  assign y17 = n3804 ;
  assign y18 = n3631 ;
  assign y19 = n3464 ;
  assign y20 = n3302 ;
  assign y21 = n3141 ;
  assign y22 = n8837 ;
  assign y23 = n2995 ;
  assign y24 = n2839 ;
  assign y25 = n2690 ;
  assign y26 = n2544 ;
  assign y27 = n2404 ;
  assign y28 = n2269 ;
  assign y29 = n2139 ;
  assign y30 = n2009 ;
  assign y31 = n1885 ;
  assign y32 = n1766 ;
  assign y33 = n8587 ;
  assign y34 = n1652 ;
  assign y35 = n1534 ;
  assign y36 = n1416 ;
  assign y37 = n1318 ;
  assign y38 = n1220 ;
  assign y39 = n1118 ;
  assign y40 = n1034 ;
  assign y41 = n941 ;
  assign y42 = n859 ;
  assign y43 = n785 ;
  assign y44 = n8324 ;
  assign y45 = n716 ;
  assign y46 = n640 ;
  assign y47 = n572 ;
  assign y48 = n514 ;
  assign y49 = n458 ;
  assign y50 = n399 ;
  assign y51 = n345 ;
  assign y52 = n302 ;
  assign y53 = n261 ;
  assign y54 = n217 ;
  assign y55 = n8069 ;
  assign y56 = n179 ;
  assign y57 = n144 ;
  assign y58 = n134 ;
  assign y59 = n136 ;
  assign y60 = n7824 ;
  assign y61 = n7575 ;
  assign y62 = n7337 ;
  assign y63 = n7089 ;
endmodule
