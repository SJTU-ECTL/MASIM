module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 ;
  assign n257 = x0 & x128 ;
  assign n258 = n257 ^ x129 ^ x1 ;
  assign n259 = ( x1 & x129 ) | ( x1 & n257 ) | ( x129 & n257 ) ;
  assign n260 = n259 ^ x130 ^ x2 ;
  assign n261 = ( x2 & x130 ) | ( x2 & n259 ) | ( x130 & n259 ) ;
  assign n262 = n261 ^ x131 ^ x3 ;
  assign n263 = ( x3 & x131 ) | ( x3 & n261 ) | ( x131 & n261 ) ;
  assign n264 = n263 ^ x132 ^ x4 ;
  assign n265 = ( x4 & x132 ) | ( x4 & n263 ) | ( x132 & n263 ) ;
  assign n266 = n265 ^ x133 ^ x5 ;
  assign n267 = ( x5 & x133 ) | ( x5 & n265 ) | ( x133 & n265 ) ;
  assign n268 = ( x6 & x134 ) | ( x6 & n267 ) | ( x134 & n267 ) ;
  assign n269 = ( x7 & x135 ) | ( x7 & n268 ) | ( x135 & n268 ) ;
  assign n270 = n269 ^ x136 ^ x8 ;
  assign n271 = ( x8 & x136 ) | ( x8 & n269 ) | ( x136 & n269 ) ;
  assign n272 = n271 ^ x137 ^ x9 ;
  assign n273 = ( x9 & x137 ) | ( x9 & n271 ) | ( x137 & n271 ) ;
  assign n274 = n273 ^ x138 ^ x10 ;
  assign n275 = ( x10 & x138 ) | ( x10 & n273 ) | ( x138 & n273 ) ;
  assign n276 = n275 ^ x139 ^ x11 ;
  assign n277 = ( x11 & x139 ) | ( x11 & n275 ) | ( x139 & n275 ) ;
  assign n278 = n277 ^ x140 ^ x12 ;
  assign n279 = ( x12 & x140 ) | ( x12 & n277 ) | ( x140 & n277 ) ;
  assign n280 = n279 ^ x141 ^ x13 ;
  assign n281 = ( x13 & x141 ) | ( x13 & n279 ) | ( x141 & n279 ) ;
  assign n282 = n281 ^ x142 ^ x14 ;
  assign n283 = ( x14 & x142 ) | ( x14 & n281 ) | ( x142 & n281 ) ;
  assign n284 = n283 ^ x143 ^ x15 ;
  assign n285 = ( x15 & x143 ) | ( x15 & n283 ) | ( x143 & n283 ) ;
  assign n286 = n285 ^ x144 ^ x16 ;
  assign n287 = n268 ^ x135 ^ x7 ;
  assign n288 = ( x16 & x144 ) | ( x16 & n285 ) | ( x144 & n285 ) ;
  assign n289 = n288 ^ x145 ^ x17 ;
  assign n290 = n267 ^ x134 ^ x6 ;
  assign n291 = ( x17 & x145 ) | ( x17 & n288 ) | ( x145 & n288 ) ;
  assign n292 = n291 ^ x146 ^ x18 ;
  assign n293 = ( x18 & x146 ) | ( x18 & n291 ) | ( x146 & n291 ) ;
  assign n294 = n293 ^ x147 ^ x19 ;
  assign n295 = ( x19 & x147 ) | ( x19 & n293 ) | ( x147 & n293 ) ;
  assign n296 = n295 ^ x148 ^ x20 ;
  assign n297 = ( x20 & x148 ) | ( x20 & n295 ) | ( x148 & n295 ) ;
  assign n298 = n297 ^ x149 ^ x21 ;
  assign n299 = ( x21 & x149 ) | ( x21 & n297 ) | ( x149 & n297 ) ;
  assign n300 = n299 ^ x150 ^ x22 ;
  assign n301 = ( x22 & x150 ) | ( x22 & n299 ) | ( x150 & n299 ) ;
  assign n302 = n301 ^ x151 ^ x23 ;
  assign n303 = ( x23 & x151 ) | ( x23 & n301 ) | ( x151 & n301 ) ;
  assign n304 = n303 ^ x152 ^ x24 ;
  assign n305 = ( x24 & x152 ) | ( x24 & n303 ) | ( x152 & n303 ) ;
  assign n306 = n305 ^ x153 ^ x25 ;
  assign n307 = ( x25 & x153 ) | ( x25 & n305 ) | ( x153 & n305 ) ;
  assign n308 = n307 ^ x154 ^ x26 ;
  assign n309 = ( x26 & x154 ) | ( x26 & n307 ) | ( x154 & n307 ) ;
  assign n310 = n309 ^ x155 ^ x27 ;
  assign n311 = ( x27 & x155 ) | ( x27 & n309 ) | ( x155 & n309 ) ;
  assign n312 = n311 ^ x156 ^ x28 ;
  assign n313 = ( x28 & x156 ) | ( x28 & n311 ) | ( x156 & n311 ) ;
  assign n314 = n313 ^ x157 ^ x29 ;
  assign n315 = ( x29 & x157 ) | ( x29 & n313 ) | ( x157 & n313 ) ;
  assign n316 = n315 ^ x158 ^ x30 ;
  assign n317 = ( x30 & x158 ) | ( x30 & n315 ) | ( x158 & n315 ) ;
  assign n318 = n317 ^ x159 ^ x31 ;
  assign n319 = ( x31 & x159 ) | ( x31 & n317 ) | ( x159 & n317 ) ;
  assign n320 = n319 ^ x160 ^ x32 ;
  assign n321 = ( x32 & x160 ) | ( x32 & n319 ) | ( x160 & n319 ) ;
  assign n322 = n321 ^ x161 ^ x33 ;
  assign n323 = ( x33 & x161 ) | ( x33 & n321 ) | ( x161 & n321 ) ;
  assign n324 = n323 ^ x162 ^ x34 ;
  assign n325 = ( x34 & x162 ) | ( x34 & n323 ) | ( x162 & n323 ) ;
  assign n326 = n325 ^ x163 ^ x35 ;
  assign n327 = ( x35 & x163 ) | ( x35 & n325 ) | ( x163 & n325 ) ;
  assign n328 = n327 ^ x164 ^ x36 ;
  assign n329 = ( x36 & x164 ) | ( x36 & n327 ) | ( x164 & n327 ) ;
  assign n330 = n329 ^ x165 ^ x37 ;
  assign n331 = ( x37 & x165 ) | ( x37 & n329 ) | ( x165 & n329 ) ;
  assign n332 = n331 ^ x166 ^ x38 ;
  assign n333 = ( x38 & x166 ) | ( x38 & n331 ) | ( x166 & n331 ) ;
  assign n334 = n333 ^ x167 ^ x39 ;
  assign n335 = ( x39 & x167 ) | ( x39 & n333 ) | ( x167 & n333 ) ;
  assign n336 = n335 ^ x168 ^ x40 ;
  assign n337 = ( x40 & x168 ) | ( x40 & n335 ) | ( x168 & n335 ) ;
  assign n338 = n337 ^ x169 ^ x41 ;
  assign n339 = ( x41 & x169 ) | ( x41 & n337 ) | ( x169 & n337 ) ;
  assign n340 = n339 ^ x170 ^ x42 ;
  assign n341 = ( x42 & x170 ) | ( x42 & n339 ) | ( x170 & n339 ) ;
  assign n342 = n341 ^ x171 ^ x43 ;
  assign n343 = ( x43 & x171 ) | ( x43 & n341 ) | ( x171 & n341 ) ;
  assign n344 = n343 ^ x172 ^ x44 ;
  assign n345 = ( x44 & x172 ) | ( x44 & n343 ) | ( x172 & n343 ) ;
  assign n346 = n345 ^ x173 ^ x45 ;
  assign n347 = ( x45 & x173 ) | ( x45 & n345 ) | ( x173 & n345 ) ;
  assign n348 = n347 ^ x174 ^ x46 ;
  assign n349 = ( x46 & x174 ) | ( x46 & n347 ) | ( x174 & n347 ) ;
  assign n350 = n349 ^ x175 ^ x47 ;
  assign n351 = ( x47 & x175 ) | ( x47 & n349 ) | ( x175 & n349 ) ;
  assign n352 = n351 ^ x176 ^ x48 ;
  assign n353 = ( x48 & x176 ) | ( x48 & n351 ) | ( x176 & n351 ) ;
  assign n354 = n353 ^ x177 ^ x49 ;
  assign n355 = ( x49 & x177 ) | ( x49 & n353 ) | ( x177 & n353 ) ;
  assign n356 = n355 ^ x178 ^ x50 ;
  assign n357 = ( x50 & x178 ) | ( x50 & n355 ) | ( x178 & n355 ) ;
  assign n358 = n357 ^ x179 ^ x51 ;
  assign n359 = ( x51 & x179 ) | ( x51 & n357 ) | ( x179 & n357 ) ;
  assign n360 = n359 ^ x180 ^ x52 ;
  assign n361 = ( x52 & x180 ) | ( x52 & n359 ) | ( x180 & n359 ) ;
  assign n362 = n361 ^ x181 ^ x53 ;
  assign n363 = ( x53 & x181 ) | ( x53 & n361 ) | ( x181 & n361 ) ;
  assign n364 = n363 ^ x182 ^ x54 ;
  assign n365 = ( x54 & x182 ) | ( x54 & n363 ) | ( x182 & n363 ) ;
  assign n366 = n365 ^ x183 ^ x55 ;
  assign n367 = ( x55 & x183 ) | ( x55 & n365 ) | ( x183 & n365 ) ;
  assign n368 = n367 ^ x184 ^ x56 ;
  assign n369 = ( x56 & x184 ) | ( x56 & n367 ) | ( x184 & n367 ) ;
  assign n370 = n369 ^ x185 ^ x57 ;
  assign n371 = ( x57 & x185 ) | ( x57 & n369 ) | ( x185 & n369 ) ;
  assign n372 = n371 ^ x186 ^ x58 ;
  assign n373 = ( x58 & x186 ) | ( x58 & n371 ) | ( x186 & n371 ) ;
  assign n374 = n373 ^ x187 ^ x59 ;
  assign n375 = ( x59 & x187 ) | ( x59 & n373 ) | ( x187 & n373 ) ;
  assign n376 = n375 ^ x188 ^ x60 ;
  assign n377 = ( x60 & x188 ) | ( x60 & n375 ) | ( x188 & n375 ) ;
  assign n378 = n377 ^ x189 ^ x61 ;
  assign n379 = ( x61 & x189 ) | ( x61 & n377 ) | ( x189 & n377 ) ;
  assign n380 = n379 ^ x190 ^ x62 ;
  assign n381 = ( x62 & x190 ) | ( x62 & n379 ) | ( x190 & n379 ) ;
  assign n382 = n381 ^ x191 ^ x63 ;
  assign n383 = ( x63 & x191 ) | ( x63 & n381 ) | ( x191 & n381 ) ;
  assign n384 = n383 ^ x192 ^ x64 ;
  assign n385 = ( x64 & x192 ) | ( x64 & n383 ) | ( x192 & n383 ) ;
  assign n386 = n385 ^ x193 ^ x65 ;
  assign n387 = ( x65 & x193 ) | ( x65 & n385 ) | ( x193 & n385 ) ;
  assign n388 = n387 ^ x194 ^ x66 ;
  assign n389 = ( x66 & x194 ) | ( x66 & n387 ) | ( x194 & n387 ) ;
  assign n390 = n389 ^ x195 ^ x67 ;
  assign n391 = ( x67 & x195 ) | ( x67 & n389 ) | ( x195 & n389 ) ;
  assign n392 = n391 ^ x196 ^ x68 ;
  assign n393 = ( x68 & x196 ) | ( x68 & n391 ) | ( x196 & n391 ) ;
  assign n394 = n393 ^ x197 ^ x69 ;
  assign n395 = ( x69 & x197 ) | ( x69 & n393 ) | ( x197 & n393 ) ;
  assign n396 = n395 ^ x198 ^ x70 ;
  assign n397 = ( x70 & x198 ) | ( x70 & n395 ) | ( x198 & n395 ) ;
  assign n398 = n397 ^ x199 ^ x71 ;
  assign n399 = ( x71 & x199 ) | ( x71 & n397 ) | ( x199 & n397 ) ;
  assign n400 = n399 ^ x200 ^ x72 ;
  assign n401 = ( x72 & x200 ) | ( x72 & n399 ) | ( x200 & n399 ) ;
  assign n402 = n401 ^ x201 ^ x73 ;
  assign n403 = ( x73 & x201 ) | ( x73 & n401 ) | ( x201 & n401 ) ;
  assign n404 = n403 ^ x202 ^ x74 ;
  assign n405 = ( x74 & x202 ) | ( x74 & n403 ) | ( x202 & n403 ) ;
  assign n406 = n405 ^ x203 ^ x75 ;
  assign n407 = ( x75 & x203 ) | ( x75 & n405 ) | ( x203 & n405 ) ;
  assign n408 = n407 ^ x204 ^ x76 ;
  assign n409 = ( x76 & x204 ) | ( x76 & n407 ) | ( x204 & n407 ) ;
  assign n410 = n409 ^ x205 ^ x77 ;
  assign n411 = ( x77 & x205 ) | ( x77 & n409 ) | ( x205 & n409 ) ;
  assign n412 = n411 ^ x206 ^ x78 ;
  assign n413 = ( x78 & x206 ) | ( x78 & n411 ) | ( x206 & n411 ) ;
  assign n414 = n413 ^ x207 ^ x79 ;
  assign n415 = ( x79 & x207 ) | ( x79 & n413 ) | ( x207 & n413 ) ;
  assign n416 = n415 ^ x208 ^ x80 ;
  assign n417 = ( x80 & x208 ) | ( x80 & n415 ) | ( x208 & n415 ) ;
  assign n418 = n417 ^ x209 ^ x81 ;
  assign n419 = ( x81 & x209 ) | ( x81 & n417 ) | ( x209 & n417 ) ;
  assign n420 = n419 ^ x210 ^ x82 ;
  assign n421 = ( x82 & x210 ) | ( x82 & n419 ) | ( x210 & n419 ) ;
  assign n422 = n421 ^ x211 ^ x83 ;
  assign n423 = ( x83 & x211 ) | ( x83 & n421 ) | ( x211 & n421 ) ;
  assign n424 = n423 ^ x212 ^ x84 ;
  assign n425 = ( x84 & x212 ) | ( x84 & n423 ) | ( x212 & n423 ) ;
  assign n426 = n425 ^ x213 ^ x85 ;
  assign n427 = ( x85 & x213 ) | ( x85 & n425 ) | ( x213 & n425 ) ;
  assign n428 = n427 ^ x214 ^ x86 ;
  assign n429 = ( x86 & x214 ) | ( x86 & n427 ) | ( x214 & n427 ) ;
  assign n430 = n429 ^ x215 ^ x87 ;
  assign n431 = ( x87 & x215 ) | ( x87 & n429 ) | ( x215 & n429 ) ;
  assign n432 = n431 ^ x216 ^ x88 ;
  assign n433 = ( x88 & x216 ) | ( x88 & n431 ) | ( x216 & n431 ) ;
  assign n434 = n433 ^ x217 ^ x89 ;
  assign n435 = ( x89 & x217 ) | ( x89 & n433 ) | ( x217 & n433 ) ;
  assign n436 = n435 ^ x218 ^ x90 ;
  assign n437 = ( x90 & x218 ) | ( x90 & n435 ) | ( x218 & n435 ) ;
  assign n438 = n437 ^ x219 ^ x91 ;
  assign n439 = ( x91 & x219 ) | ( x91 & n437 ) | ( x219 & n437 ) ;
  assign n440 = ( x92 & x220 ) | ( x92 & n439 ) | ( x220 & n439 ) ;
  assign n441 = ( x93 & x221 ) | ( x93 & n440 ) | ( x221 & n440 ) ;
  assign n442 = ( x94 & x222 ) | ( x94 & n441 ) | ( x222 & n441 ) ;
  assign n443 = ( x95 & x223 ) | ( x95 & n442 ) | ( x223 & n442 ) ;
  assign n444 = ( x96 & x224 ) | ( x96 & n443 ) | ( x224 & n443 ) ;
  assign n445 = ( x97 & x225 ) | ( x97 & n444 ) | ( x225 & n444 ) ;
  assign n446 = ( x98 & x226 ) | ( x98 & n445 ) | ( x226 & n445 ) ;
  assign n447 = ( x99 & x227 ) | ( x99 & n446 ) | ( x227 & n446 ) ;
  assign n448 = ( x100 & x228 ) | ( x100 & n447 ) | ( x228 & n447 ) ;
  assign n449 = ( x101 & x229 ) | ( x101 & n448 ) | ( x229 & n448 ) ;
  assign n450 = ( x102 & x230 ) | ( x102 & n449 ) | ( x230 & n449 ) ;
  assign n451 = ( x103 & x231 ) | ( x103 & n450 ) | ( x231 & n450 ) ;
  assign n452 = ( x104 & x232 ) | ( x104 & n451 ) | ( x232 & n451 ) ;
  assign n453 = ( x105 & x233 ) | ( x105 & n452 ) | ( x233 & n452 ) ;
  assign n454 = ( x106 & x234 ) | ( x106 & n453 ) | ( x234 & n453 ) ;
  assign n455 = ( x107 & x235 ) | ( x107 & n454 ) | ( x235 & n454 ) ;
  assign n456 = ( x108 & x236 ) | ( x108 & n455 ) | ( x236 & n455 ) ;
  assign n457 = ( x109 & x237 ) | ( x109 & n456 ) | ( x237 & n456 ) ;
  assign n458 = ( x110 & x238 ) | ( x110 & n457 ) | ( x238 & n457 ) ;
  assign n459 = ( x111 & x239 ) | ( x111 & n458 ) | ( x239 & n458 ) ;
  assign n460 = ( x112 & x240 ) | ( x112 & n459 ) | ( x240 & n459 ) ;
  assign n461 = ( x113 & x241 ) | ( x113 & n460 ) | ( x241 & n460 ) ;
  assign n462 = ( x114 & x242 ) | ( x114 & n461 ) | ( x242 & n461 ) ;
  assign n463 = ( x115 & x243 ) | ( x115 & n462 ) | ( x243 & n462 ) ;
  assign n464 = ( x116 & x244 ) | ( x116 & n463 ) | ( x244 & n463 ) ;
  assign n465 = ( x117 & x245 ) | ( x117 & n464 ) | ( x245 & n464 ) ;
  assign n466 = ( x118 & x246 ) | ( x118 & n465 ) | ( x246 & n465 ) ;
  assign n467 = ( x119 & x247 ) | ( x119 & n466 ) | ( x247 & n466 ) ;
  assign n468 = ( x120 & x248 ) | ( x120 & n467 ) | ( x248 & n467 ) ;
  assign n469 = ( x121 & x249 ) | ( x121 & n468 ) | ( x249 & n468 ) ;
  assign n470 = ( x122 & x250 ) | ( x122 & n469 ) | ( x250 & n469 ) ;
  assign n471 = ( x123 & x251 ) | ( x123 & n470 ) | ( x251 & n470 ) ;
  assign n472 = ( x124 & x252 ) | ( x124 & n471 ) | ( x252 & n471 ) ;
  assign n473 = ( x125 & x253 ) | ( x125 & n472 ) | ( x253 & n472 ) ;
  assign n474 = ( x126 & x254 ) | ( x126 & n473 ) | ( x254 & n473 ) ;
  assign n475 = n474 ^ x255 ^ x127 ;
  assign n476 = n439 ^ x220 ^ x92 ;
  assign n477 = n440 ^ x221 ^ x93 ;
  assign n478 = n441 ^ x222 ^ x94 ;
  assign n479 = n442 ^ x223 ^ x95 ;
  assign n480 = n443 ^ x224 ^ x96 ;
  assign n481 = n444 ^ x225 ^ x97 ;
  assign n482 = n445 ^ x226 ^ x98 ;
  assign n483 = n446 ^ x227 ^ x99 ;
  assign n484 = n447 ^ x228 ^ x100 ;
  assign n485 = n448 ^ x229 ^ x101 ;
  assign n486 = n449 ^ x230 ^ x102 ;
  assign n487 = n450 ^ x231 ^ x103 ;
  assign n488 = n451 ^ x232 ^ x104 ;
  assign n489 = n452 ^ x233 ^ x105 ;
  assign n490 = n453 ^ x234 ^ x106 ;
  assign n491 = n454 ^ x235 ^ x107 ;
  assign n492 = n455 ^ x236 ^ x108 ;
  assign n493 = n456 ^ x237 ^ x109 ;
  assign n494 = n457 ^ x238 ^ x110 ;
  assign n495 = n458 ^ x239 ^ x111 ;
  assign n496 = n459 ^ x240 ^ x112 ;
  assign n497 = n460 ^ x241 ^ x113 ;
  assign n498 = ( x127 & x255 ) | ( x127 & n474 ) | ( x255 & n474 ) ;
  assign n499 = n462 ^ x243 ^ x115 ;
  assign n500 = n463 ^ x244 ^ x116 ;
  assign n501 = n464 ^ x245 ^ x117 ;
  assign n502 = n465 ^ x246 ^ x118 ;
  assign n503 = n466 ^ x247 ^ x119 ;
  assign n504 = n467 ^ x248 ^ x120 ;
  assign n505 = n468 ^ x249 ^ x121 ;
  assign n506 = n469 ^ x250 ^ x122 ;
  assign n507 = n470 ^ x251 ^ x123 ;
  assign n508 = n471 ^ x252 ^ x124 ;
  assign n509 = n472 ^ x253 ^ x125 ;
  assign n510 = x128 ^ x0 ^ 1'b0 ;
  assign n511 = n461 ^ x242 ^ x114 ;
  assign n512 = n473 ^ x254 ^ x126 ;
  assign y0 = n510 ;
  assign y1 = n258 ;
  assign y2 = n260 ;
  assign y3 = n262 ;
  assign y4 = n264 ;
  assign y5 = n266 ;
  assign y6 = n290 ;
  assign y7 = n287 ;
  assign y8 = n270 ;
  assign y9 = n272 ;
  assign y10 = n274 ;
  assign y11 = n276 ;
  assign y12 = n278 ;
  assign y13 = n280 ;
  assign y14 = n282 ;
  assign y15 = n284 ;
  assign y16 = n286 ;
  assign y17 = n289 ;
  assign y18 = n292 ;
  assign y19 = n294 ;
  assign y20 = n296 ;
  assign y21 = n298 ;
  assign y22 = n300 ;
  assign y23 = n302 ;
  assign y24 = n304 ;
  assign y25 = n306 ;
  assign y26 = n308 ;
  assign y27 = n310 ;
  assign y28 = n312 ;
  assign y29 = n314 ;
  assign y30 = n316 ;
  assign y31 = n318 ;
  assign y32 = n320 ;
  assign y33 = n322 ;
  assign y34 = n324 ;
  assign y35 = n326 ;
  assign y36 = n328 ;
  assign y37 = n330 ;
  assign y38 = n332 ;
  assign y39 = n334 ;
  assign y40 = n336 ;
  assign y41 = n338 ;
  assign y42 = n340 ;
  assign y43 = n342 ;
  assign y44 = n344 ;
  assign y45 = n346 ;
  assign y46 = n348 ;
  assign y47 = n350 ;
  assign y48 = n352 ;
  assign y49 = n354 ;
  assign y50 = n356 ;
  assign y51 = n358 ;
  assign y52 = n360 ;
  assign y53 = n362 ;
  assign y54 = n364 ;
  assign y55 = n366 ;
  assign y56 = n368 ;
  assign y57 = n370 ;
  assign y58 = n372 ;
  assign y59 = n374 ;
  assign y60 = n376 ;
  assign y61 = n378 ;
  assign y62 = n380 ;
  assign y63 = n382 ;
  assign y64 = n384 ;
  assign y65 = n386 ;
  assign y66 = n388 ;
  assign y67 = n390 ;
  assign y68 = n392 ;
  assign y69 = n394 ;
  assign y70 = n396 ;
  assign y71 = n398 ;
  assign y72 = n400 ;
  assign y73 = n402 ;
  assign y74 = n404 ;
  assign y75 = n406 ;
  assign y76 = n408 ;
  assign y77 = n410 ;
  assign y78 = n412 ;
  assign y79 = n414 ;
  assign y80 = n416 ;
  assign y81 = n418 ;
  assign y82 = n420 ;
  assign y83 = n422 ;
  assign y84 = n424 ;
  assign y85 = n426 ;
  assign y86 = n428 ;
  assign y87 = n430 ;
  assign y88 = n432 ;
  assign y89 = n434 ;
  assign y90 = n436 ;
  assign y91 = n438 ;
  assign y92 = n476 ;
  assign y93 = n477 ;
  assign y94 = n478 ;
  assign y95 = n479 ;
  assign y96 = n480 ;
  assign y97 = n481 ;
  assign y98 = n482 ;
  assign y99 = n483 ;
  assign y100 = n484 ;
  assign y101 = n485 ;
  assign y102 = n486 ;
  assign y103 = n487 ;
  assign y104 = n488 ;
  assign y105 = n489 ;
  assign y106 = n490 ;
  assign y107 = n491 ;
  assign y108 = n492 ;
  assign y109 = n493 ;
  assign y110 = n494 ;
  assign y111 = n495 ;
  assign y112 = n496 ;
  assign y113 = n497 ;
  assign y114 = n511 ;
  assign y115 = n499 ;
  assign y116 = n500 ;
  assign y117 = n501 ;
  assign y118 = n502 ;
  assign y119 = n503 ;
  assign y120 = n504 ;
  assign y121 = n505 ;
  assign y122 = n506 ;
  assign y123 = n507 ;
  assign y124 = n508 ;
  assign y125 = n509 ;
  assign y126 = n512 ;
  assign y127 = n475 ;
  assign y128 = n498 ;
endmodule
