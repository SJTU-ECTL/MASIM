module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 ;
  assign n61 = x3 | x4 ;
  assign n62 = x1 | x2 ;
  assign n63 = n61 | n62 ;
  assign n64 = x5 | x6 ;
  assign n65 = x10 ^ x9 ^ 1'b0 ;
  assign n66 = ( x9 & x10 ) | ( x9 & x11 ) | ( x10 & x11 ) ;
  assign n67 = n63 | n64 ;
  assign n68 = ( x11 & n65 ) | ( x11 & n66 ) | ( n65 & n66 ) ;
  assign n69 = ( ~x12 & x13 ) | ( ~x12 & n68 ) | ( x13 & n68 ) ;
  assign n70 = n69 ^ x12 ^ 1'b0 ;
  assign n71 = ( x12 & n69 ) | ( x12 & n70 ) | ( n69 & n70 ) ;
  assign n72 = x7 | x8 ;
  assign n73 = n67 | n72 ;
  assign n74 = n68 ^ x12 ^ 1'b0 ;
  assign n75 = ( x11 & n65 ) | ( x11 & n73 ) | ( n65 & n73 ) ;
  assign n76 = ~n73 & n75 ;
  assign n77 = n71 ^ x14 ^ 1'b0 ;
  assign n78 = ( x13 & n74 ) | ( x13 & n76 ) | ( n74 & n76 ) ;
  assign n79 = ~x13 & n78 ;
  assign n80 = ~n77 & n79 ;
  assign n81 = x14 & n71 ;
  assign n82 = ( x15 & x16 ) | ( x15 & n81 ) | ( x16 & n81 ) ;
  assign n83 = x16 | n82 ;
  assign n84 = x17 & n83 ;
  assign n85 = n84 ^ x18 ^ 1'b0 ;
  assign n86 = n66 ^ x11 ^ 1'b0 ;
  assign n87 = ( ~x15 & x16 ) | ( ~x15 & n81 ) | ( x16 & n81 ) ;
  assign n88 = n87 ^ n81 ^ 1'b0 ;
  assign n89 = n83 ^ x17 ^ 1'b0 ;
  assign n90 = n80 & n88 ;
  assign n91 = n85 & ~n89 ;
  assign n92 = n90 & n91 ;
  assign n93 = n81 ^ x15 ^ 1'b0 ;
  assign n94 = x18 | n84 ;
  assign n95 = x19 & n94 ;
  assign n96 = n94 ^ x19 ^ 1'b0 ;
  assign n97 = ~n85 & n96 ;
  assign n98 = n92 & ~n96 ;
  assign n99 = ( ~x20 & x21 ) | ( ~x20 & n95 ) | ( x21 & n95 ) ;
  assign n100 = n99 ^ n95 ^ 1'b0 ;
  assign n101 = n98 & n100 ;
  assign n102 = ( x20 & x21 ) | ( x20 & n95 ) | ( x21 & n95 ) ;
  assign n103 = n95 ^ x20 ^ 1'b0 ;
  assign n104 = x21 | n102 ;
  assign n105 = n104 ^ x22 ^ 1'b0 ;
  assign n106 = x22 | n104 ;
  assign n107 = n101 & n105 ;
  assign n108 = x23 & n106 ;
  assign n109 = x24 & n108 ;
  assign n110 = n106 ^ x23 ^ 1'b0 ;
  assign n111 = ( x25 & x26 ) | ( x25 & n109 ) | ( x26 & n109 ) ;
  assign n112 = n107 & ~n110 ;
  assign n113 = x26 | n111 ;
  assign n114 = x27 & n113 ;
  assign n115 = n108 ^ x24 ^ 1'b0 ;
  assign n116 = n110 & n115 ;
  assign n117 = n112 & ~n115 ;
  assign n118 = ( ~x25 & x26 ) | ( ~x25 & n109 ) | ( x26 & n109 ) ;
  assign n119 = n118 ^ n109 ^ 1'b0 ;
  assign n120 = n117 & n119 ;
  assign n121 = x28 & x29 ;
  assign n122 = n114 & n121 ;
  assign n123 = n113 ^ x27 ^ 1'b0 ;
  assign n124 = n120 & ~n123 ;
  assign n125 = n114 ^ x28 ^ 1'b0 ;
  assign n126 = n124 & ~n125 ;
  assign n127 = ~x9 & n125 ;
  assign n128 = x29 & n123 ;
  assign n129 = x9 & n126 ;
  assign n130 = n109 ^ x25 ^ 1'b0 ;
  assign n131 = n127 & n128 ;
  assign n132 = x5 & x6 ;
  assign n133 = ( x26 & n130 ) | ( x26 & n131 ) | ( n130 & n131 ) ;
  assign n134 = ~x26 & n133 ;
  assign n135 = n116 & n134 ;
  assign n136 = ~n105 & n135 ;
  assign n137 = ( x21 & n103 ) | ( x21 & n136 ) | ( n103 & n136 ) ;
  assign n138 = n122 & ~n129 ;
  assign n139 = x7 & x8 ;
  assign n140 = ~x21 & n137 ;
  assign n141 = n97 & n140 ;
  assign n142 = n89 & n141 ;
  assign n143 = ( x16 & n93 ) | ( x16 & n142 ) | ( n93 & n142 ) ;
  assign n144 = ~x16 & n143 ;
  assign n145 = n77 & n144 ;
  assign n146 = ~n70 & n145 ;
  assign n147 = x1 & x2 ;
  assign n148 = n86 & n146 ;
  assign n149 = n139 & n148 ;
  assign n150 = n132 & n149 ;
  assign n151 = x3 & x4 ;
  assign n152 = n150 & n151 ;
  assign n153 = n147 & n152 ;
  assign n154 = x0 & n153 ;
  assign n155 = n122 | n154 ;
  assign n156 = x31 | x32 ;
  assign n157 = ( x39 & x40 ) | ( x39 & x41 ) | ( x40 & x41 ) ;
  assign n158 = x35 | x36 ;
  assign n159 = x37 | x38 ;
  assign n160 = x33 | x34 ;
  assign n161 = x40 ^ x39 ^ 1'b0 ;
  assign n162 = ( x41 & n157 ) | ( x41 & n161 ) | ( n157 & n161 ) ;
  assign n163 = ( ~x42 & x43 ) | ( ~x42 & n162 ) | ( x43 & n162 ) ;
  assign n164 = n163 ^ x42 ^ 1'b0 ;
  assign n165 = ( x42 & n163 ) | ( x42 & n164 ) | ( n163 & n164 ) ;
  assign n166 = x44 & n165 ;
  assign n167 = ( ~x45 & x46 ) | ( ~x45 & n166 ) | ( x46 & n166 ) ;
  assign n168 = n157 ^ x41 ^ 1'b0 ;
  assign n169 = n156 | n160 ;
  assign n170 = n158 | n169 ;
  assign n171 = ( x45 & x46 ) | ( x45 & n166 ) | ( x46 & n166 ) ;
  assign n172 = n166 ^ x45 ^ 1'b0 ;
  assign n173 = n162 ^ x42 ^ 1'b0 ;
  assign n174 = x46 | n171 ;
  assign n175 = n167 ^ n166 ^ 1'b0 ;
  assign n176 = n174 ^ x47 ^ 1'b0 ;
  assign n177 = x47 & n174 ;
  assign n178 = n159 | n170 ;
  assign n179 = ( x41 & n161 ) | ( x41 & n178 ) | ( n161 & n178 ) ;
  assign n180 = ~n178 & n179 ;
  assign n181 = n177 ^ x48 ^ 1'b0 ;
  assign n182 = n165 ^ x44 ^ 1'b0 ;
  assign n183 = ( x43 & n173 ) | ( x43 & n180 ) | ( n173 & n180 ) ;
  assign n184 = x48 | n177 ;
  assign n185 = x49 & n184 ;
  assign n186 = ( x50 & x51 ) | ( x50 & n185 ) | ( x51 & n185 ) ;
  assign n187 = ~x43 & n183 ;
  assign n188 = ~n182 & n187 ;
  assign n189 = n175 & n188 ;
  assign n190 = ~n176 & n181 ;
  assign n191 = n184 ^ x49 ^ 1'b0 ;
  assign n192 = n189 & n190 ;
  assign n193 = x51 | n186 ;
  assign n194 = ( ~x50 & x51 ) | ( ~x50 & n185 ) | ( x51 & n185 ) ;
  assign n195 = n194 ^ n185 ^ 1'b0 ;
  assign n196 = n185 ^ x50 ^ 1'b0 ;
  assign n197 = ~n191 & n192 ;
  assign n198 = n195 & n197 ;
  assign n199 = n193 ^ x52 ^ 1'b0 ;
  assign n200 = n198 & n199 ;
  assign n201 = x52 | n193 ;
  assign n202 = ~n181 & n191 ;
  assign n203 = x53 & n201 ;
  assign n204 = n201 ^ x53 ^ 1'b0 ;
  assign n205 = n200 & ~n204 ;
  assign n206 = n203 ^ x54 ^ 1'b0 ;
  assign n207 = x54 & n203 ;
  assign n208 = n205 & ~n206 ;
  assign n209 = ( x55 & x56 ) | ( x55 & n207 ) | ( x56 & n207 ) ;
  assign n210 = x56 | n209 ;
  assign n211 = ( ~x55 & x56 ) | ( ~x55 & n207 ) | ( x56 & n207 ) ;
  assign n212 = n204 & n206 ;
  assign n213 = x57 & n210 ;
  assign n214 = n211 ^ n207 ^ 1'b0 ;
  assign n215 = n210 ^ x57 ^ 1'b0 ;
  assign n216 = n208 & n214 ;
  assign n217 = ~n215 & n216 ;
  assign n218 = n213 ^ x58 ^ 1'b0 ;
  assign n219 = n217 & ~n218 ;
  assign n220 = n215 & n218 ;
  assign n221 = n207 ^ x55 ^ 1'b0 ;
  assign n222 = x30 & x59 ;
  assign n223 = ~x39 & n222 ;
  assign n224 = n220 & n223 ;
  assign n225 = x35 & x36 ;
  assign n226 = ( x56 & n221 ) | ( x56 & n224 ) | ( n221 & n224 ) ;
  assign n227 = ~x56 & n226 ;
  assign n228 = n212 & n227 ;
  assign n229 = ~n199 & n228 ;
  assign n230 = ( x51 & n196 ) | ( x51 & n229 ) | ( n196 & n229 ) ;
  assign n231 = x58 & x59 ;
  assign n232 = x39 & n219 ;
  assign n233 = ~x0 & n232 ;
  assign n234 = n213 & n231 ;
  assign n235 = ~x30 & n233 ;
  assign n236 = n234 | n235 ;
  assign n237 = x31 & x32 ;
  assign n238 = x0 & ~n234 ;
  assign n239 = ~x51 & n230 ;
  assign n240 = n202 & n239 ;
  assign n241 = ~n138 & n155 ;
  assign n242 = n234 & n241 ;
  assign n243 = n176 & n240 ;
  assign n244 = ( x0 & x30 ) | ( x0 & ~n232 ) | ( x30 & ~n232 ) ;
  assign n245 = ~n232 & n242 ;
  assign n246 = ( n242 & n244 ) | ( n242 & n245 ) | ( n244 & n245 ) ;
  assign n247 = x37 & x38 ;
  assign n248 = ( x46 & n172 ) | ( x46 & n243 ) | ( n172 & n243 ) ;
  assign n249 = ~x46 & n248 ;
  assign n250 = x33 & x34 ;
  assign n251 = n182 & n249 ;
  assign n252 = ~n164 & n251 ;
  assign n253 = n168 & n252 ;
  assign n254 = n247 & n253 ;
  assign n255 = n225 & n254 ;
  assign n256 = n250 & n255 ;
  assign n257 = n237 & n256 ;
  assign n258 = ( ~n235 & n236 ) | ( ~n235 & n257 ) | ( n236 & n257 ) ;
  assign n259 = n155 & n258 ;
  assign n260 = ~n238 & n259 ;
  assign n261 = n138 | n260 ;
  assign y0 = ~n241 ;
  assign y1 = ~n261 ;
  assign y2 = n246 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
