module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 ;
  assign n9 = x4 | x5 ;
  assign n10 = ~x6 & x7 ;
  assign n11 = ~n9 & n10 ;
  assign n12 = x0 & x2 ;
  assign n13 = x0 | x2 ;
  assign n14 = x1 | x3 ;
  assign n15 = x1 & ~x3 ;
  assign n16 = n13 | n14 ;
  assign n17 = ~n13 & n15 ;
  assign n18 = ~x0 & x2 ;
  assign n19 = ~n14 & n18 ;
  assign n20 = x0 & ~x2 ;
  assign n21 = ~n14 & n20 ;
  assign n22 = n15 & n20 ;
  assign n23 = n15 & n18 ;
  assign n24 = n12 & n15 ;
  assign n25 = ~x1 & x3 ;
  assign n26 = ~n13 & n25 ;
  assign n27 = n20 & n25 ;
  assign n28 = x1 & x3 ;
  assign n29 = ~n13 & n28 ;
  assign n30 = n20 & n28 ;
  assign n31 = n18 & n25 ;
  assign n32 = n12 & n25 ;
  assign n33 = n18 & n28 ;
  assign n34 = n12 & n28 ;
  assign n35 = x4 & ~x5 ;
  assign n36 = n10 & n35 ;
  assign n37 = ~x4 & x5 ;
  assign n38 = n10 & n37 ;
  assign n39 = n21 & n38 ;
  assign n40 = x4 & x5 ;
  assign n41 = n10 & n40 ;
  assign n42 = x6 & x7 ;
  assign n43 = ~n9 & n42 ;
  assign n44 = n35 & n42 ;
  assign n45 = n37 & n42 ;
  assign n46 = n40 & n42 ;
  assign n47 = x6 | x7 ;
  assign n48 = n9 | n47 ;
  assign n49 = n21 & ~n48 ;
  assign n50 = n19 & ~n48 ;
  assign n51 = n35 & ~n47 ;
  assign n52 = n21 & n51 ;
  assign n53 = n37 & ~n47 ;
  assign n54 = n40 & ~n47 ;
  assign n55 = x6 & ~x7 ;
  assign n56 = ~n9 & n55 ;
  assign n57 = n35 & n55 ;
  assign n58 = n29 & n57 ;
  assign n59 = n30 & n57 ;
  assign n60 = n31 & n57 ;
  assign n61 = n32 & n57 ;
  assign n62 = n33 & n57 ;
  assign n63 = n34 & n57 ;
  assign n64 = n37 & n55 ;
  assign n65 = ~n16 & n64 ;
  assign n66 = n17 & n64 ;
  assign n67 = n22 & n64 ;
  assign n68 = n40 & n55 ;
  assign n69 = n12 & ~n14 ;
  assign n70 = n64 & n69 ;
  assign n71 = n11 & n21 ;
  assign n72 = n11 & n19 ;
  assign n73 = n21 & n36 ;
  assign n74 = n19 & n36 ;
  assign n75 = n19 & n38 ;
  assign n76 = n21 & n41 ;
  assign n77 = n19 & n41 ;
  assign n78 = n21 & n43 ;
  assign n79 = n19 & n43 ;
  assign n80 = n19 & n44 ;
  assign n81 = n21 & n45 ;
  assign n82 = n19 & n45 ;
  assign n83 = n21 & n46 ;
  assign n84 = n19 & n46 ;
  assign n85 = n19 & n51 ;
  assign n86 = n21 & n53 ;
  assign n87 = n19 & n53 ;
  assign n88 = n30 & n53 ;
  assign n89 = ~n16 & n54 ;
  assign n90 = n21 & n54 ;
  assign n91 = n17 & n54 ;
  assign n92 = n22 & n54 ;
  assign n93 = n19 & n54 ;
  assign n94 = n54 & n69 ;
  assign n95 = n23 & n54 ;
  assign n96 = n24 & n54 ;
  assign n97 = n26 & n54 ;
  assign n98 = n27 & n54 ;
  assign n99 = n29 & n54 ;
  assign n100 = n30 & n54 ;
  assign n101 = n31 & n54 ;
  assign n102 = n32 & n54 ;
  assign n103 = n33 & n54 ;
  assign n104 = n34 & n54 ;
  assign n105 = ~n16 & n56 ;
  assign n106 = n21 & n56 ;
  assign n107 = n17 & n56 ;
  assign n108 = n22 & n56 ;
  assign n109 = n19 & n56 ;
  assign n110 = n56 & n69 ;
  assign n111 = n23 & n56 ;
  assign n112 = n24 & n56 ;
  assign n113 = n26 & n56 ;
  assign n114 = n27 & n56 ;
  assign n115 = n29 & n56 ;
  assign n116 = n30 & n56 ;
  assign n117 = n31 & n56 ;
  assign n118 = n32 & n56 ;
  assign n119 = n33 & n56 ;
  assign n120 = n34 & n56 ;
  assign n121 = ~n16 & n57 ;
  assign n122 = n21 & n57 ;
  assign n123 = n17 & n57 ;
  assign n124 = n22 & n57 ;
  assign n125 = n19 & n57 ;
  assign n126 = n57 & n69 ;
  assign n127 = n23 & n57 ;
  assign n128 = n24 & n57 ;
  assign n129 = n26 & n57 ;
  assign n130 = n27 & n57 ;
  assign n131 = n21 & n64 ;
  assign n132 = n19 & n64 ;
  assign n133 = n23 & n64 ;
  assign n134 = n24 & n64 ;
  assign n135 = n26 & n64 ;
  assign n136 = n27 & n64 ;
  assign n137 = n29 & n64 ;
  assign n138 = n30 & n64 ;
  assign n139 = n31 & n64 ;
  assign n140 = n32 & n64 ;
  assign n141 = n33 & n64 ;
  assign n142 = n34 & n64 ;
  assign n143 = n21 & n44 ;
  assign n144 = n21 & n68 ;
  assign n145 = n19 & n68 ;
  assign n146 = n11 & ~n16 ;
  assign n147 = n11 & n22 ;
  assign n148 = n11 & n69 ;
  assign n149 = n11 & n23 ;
  assign n150 = n11 & n24 ;
  assign n151 = n11 & n26 ;
  assign n152 = n11 & n27 ;
  assign n153 = n11 & n29 ;
  assign n154 = n11 & n30 ;
  assign n155 = n11 & n31 ;
  assign n156 = n11 & n32 ;
  assign n157 = n11 & n33 ;
  assign n158 = n11 & n34 ;
  assign n159 = n30 & n36 ;
  assign n160 = n32 & n36 ;
  assign n161 = n33 & n36 ;
  assign n162 = n34 & n36 ;
  assign n163 = ~n16 & n38 ;
  assign n164 = n17 & n38 ;
  assign n165 = n22 & n38 ;
  assign n166 = n38 & n69 ;
  assign n167 = n23 & n38 ;
  assign n168 = n24 & n38 ;
  assign n169 = n26 & n38 ;
  assign n170 = n27 & n38 ;
  assign n171 = n29 & n38 ;
  assign n172 = n30 & n38 ;
  assign n173 = n31 & n38 ;
  assign n174 = n32 & n38 ;
  assign n175 = n33 & n38 ;
  assign n176 = n34 & n38 ;
  assign n177 = n30 & n41 ;
  assign n178 = n32 & n41 ;
  assign n179 = n33 & n41 ;
  assign n180 = n34 & n41 ;
  assign n181 = n30 & n43 ;
  assign n182 = n32 & n43 ;
  assign n183 = n33 & n43 ;
  assign n184 = n34 & n43 ;
  assign n185 = n30 & n44 ;
  assign n186 = n32 & n44 ;
  assign n187 = n33 & n44 ;
  assign n188 = n34 & n44 ;
  assign n189 = n30 & n45 ;
  assign n190 = n32 & n45 ;
  assign n191 = n33 & n45 ;
  assign n192 = n34 & n45 ;
  assign n193 = n30 & n46 ;
  assign n194 = n32 & n46 ;
  assign n195 = n33 & n46 ;
  assign n196 = n34 & n46 ;
  assign n197 = n30 & ~n48 ;
  assign n198 = n32 & ~n48 ;
  assign n199 = n33 & ~n48 ;
  assign n200 = n34 & ~n48 ;
  assign n201 = n30 & n51 ;
  assign n202 = n32 & n51 ;
  assign n203 = n33 & n51 ;
  assign n204 = n34 & n51 ;
  assign n205 = n32 & n53 ;
  assign n206 = n33 & n53 ;
  assign n207 = n34 & n53 ;
  assign n208 = ~n16 & n68 ;
  assign n209 = n11 & n17 ;
  assign n210 = n17 & n68 ;
  assign n211 = n22 & n68 ;
  assign n212 = n68 & n69 ;
  assign n213 = n23 & n68 ;
  assign n214 = n24 & n68 ;
  assign n215 = n26 & n68 ;
  assign n216 = n27 & n68 ;
  assign n217 = n29 & n68 ;
  assign n218 = n30 & n68 ;
  assign n219 = n32 & n68 ;
  assign n220 = n33 & n68 ;
  assign n221 = n34 & n68 ;
  assign n222 = ~n16 & n46 ;
  assign n223 = n17 & n46 ;
  assign n224 = n22 & n46 ;
  assign n225 = n46 & n69 ;
  assign n226 = n23 & n46 ;
  assign n227 = n24 & n46 ;
  assign n228 = n26 & n46 ;
  assign n229 = n27 & n46 ;
  assign n230 = n29 & n46 ;
  assign n231 = n31 & n46 ;
  assign n232 = n16 | n48 ;
  assign n233 = n17 & ~n48 ;
  assign n234 = n22 & ~n48 ;
  assign n235 = ~n48 & n69 ;
  assign n236 = n23 & ~n48 ;
  assign n237 = n24 & ~n48 ;
  assign n238 = n26 & ~n48 ;
  assign n239 = n27 & ~n48 ;
  assign n240 = n29 & ~n48 ;
  assign n241 = n31 & ~n48 ;
  assign n242 = ~n16 & n51 ;
  assign n243 = n17 & n51 ;
  assign n244 = n22 & n51 ;
  assign n245 = n51 & n69 ;
  assign n246 = n23 & n51 ;
  assign n247 = n24 & n51 ;
  assign n248 = n26 & n51 ;
  assign n249 = n27 & n51 ;
  assign n250 = n29 & n51 ;
  assign n251 = n31 & n51 ;
  assign n252 = ~n16 & n53 ;
  assign n253 = n17 & n53 ;
  assign n254 = n22 & n53 ;
  assign n255 = n53 & n69 ;
  assign n256 = n23 & n53 ;
  assign n257 = n24 & n53 ;
  assign n258 = n26 & n53 ;
  assign n259 = n27 & n53 ;
  assign n260 = n29 & n53 ;
  assign n261 = n31 & n53 ;
  assign n262 = n31 & n68 ;
  assign n263 = ~n16 & n36 ;
  assign n264 = n17 & n36 ;
  assign n265 = n22 & n36 ;
  assign n266 = n36 & n69 ;
  assign n267 = n23 & n36 ;
  assign n268 = n24 & n36 ;
  assign n269 = n26 & n36 ;
  assign n270 = n29 & n36 ;
  assign n271 = n31 & n36 ;
  assign n272 = ~n16 & n41 ;
  assign n273 = n17 & n41 ;
  assign n274 = n22 & n41 ;
  assign n275 = n41 & n69 ;
  assign n276 = n23 & n41 ;
  assign n277 = n24 & n41 ;
  assign n278 = n26 & n41 ;
  assign n279 = n27 & n41 ;
  assign n280 = n29 & n41 ;
  assign n281 = n31 & n41 ;
  assign n282 = n27 & n36 ;
  assign n283 = ~n16 & n43 ;
  assign n284 = n17 & n43 ;
  assign n285 = n22 & n43 ;
  assign n286 = n43 & n69 ;
  assign n287 = n23 & n43 ;
  assign n288 = n24 & n43 ;
  assign n289 = n26 & n43 ;
  assign n290 = n27 & n43 ;
  assign n291 = n29 & n43 ;
  assign n292 = n31 & n43 ;
  assign n293 = ~n16 & n44 ;
  assign n294 = n17 & n44 ;
  assign n295 = n22 & n44 ;
  assign n296 = n44 & n69 ;
  assign n297 = n23 & n44 ;
  assign n298 = n24 & n44 ;
  assign n299 = n26 & n44 ;
  assign n300 = n27 & n44 ;
  assign n301 = n29 & n44 ;
  assign n302 = n31 & n44 ;
  assign n303 = ~n16 & n45 ;
  assign n304 = n17 & n45 ;
  assign n305 = n22 & n45 ;
  assign n306 = n45 & n69 ;
  assign n307 = n23 & n45 ;
  assign n308 = n24 & n45 ;
  assign n309 = n26 & n45 ;
  assign n310 = n27 & n45 ;
  assign n311 = n29 & n45 ;
  assign n312 = n31 & n45 ;
  assign y0 = n146 ;
  assign y1 = n71 ;
  assign y2 = n209 ;
  assign y3 = n147 ;
  assign y4 = n72 ;
  assign y5 = n148 ;
  assign y6 = n149 ;
  assign y7 = n150 ;
  assign y8 = n151 ;
  assign y9 = n152 ;
  assign y10 = n153 ;
  assign y11 = n154 ;
  assign y12 = n155 ;
  assign y13 = n156 ;
  assign y14 = n157 ;
  assign y15 = n158 ;
  assign y16 = n263 ;
  assign y17 = n73 ;
  assign y18 = n264 ;
  assign y19 = n265 ;
  assign y20 = n74 ;
  assign y21 = n266 ;
  assign y22 = n267 ;
  assign y23 = n268 ;
  assign y24 = n269 ;
  assign y25 = n282 ;
  assign y26 = n270 ;
  assign y27 = n159 ;
  assign y28 = n271 ;
  assign y29 = n160 ;
  assign y30 = n161 ;
  assign y31 = n162 ;
  assign y32 = n163 ;
  assign y33 = n39 ;
  assign y34 = n164 ;
  assign y35 = n165 ;
  assign y36 = n75 ;
  assign y37 = n166 ;
  assign y38 = n167 ;
  assign y39 = n168 ;
  assign y40 = n169 ;
  assign y41 = n170 ;
  assign y42 = n171 ;
  assign y43 = n172 ;
  assign y44 = n173 ;
  assign y45 = n174 ;
  assign y46 = n175 ;
  assign y47 = n176 ;
  assign y48 = n272 ;
  assign y49 = n76 ;
  assign y50 = n273 ;
  assign y51 = n274 ;
  assign y52 = n77 ;
  assign y53 = n275 ;
  assign y54 = n276 ;
  assign y55 = n277 ;
  assign y56 = n278 ;
  assign y57 = n279 ;
  assign y58 = n280 ;
  assign y59 = n177 ;
  assign y60 = n281 ;
  assign y61 = n178 ;
  assign y62 = n179 ;
  assign y63 = n180 ;
  assign y64 = n283 ;
  assign y65 = n78 ;
  assign y66 = n284 ;
  assign y67 = n285 ;
  assign y68 = n79 ;
  assign y69 = n286 ;
  assign y70 = n287 ;
  assign y71 = n288 ;
  assign y72 = n289 ;
  assign y73 = n290 ;
  assign y74 = n291 ;
  assign y75 = n181 ;
  assign y76 = n292 ;
  assign y77 = n182 ;
  assign y78 = n183 ;
  assign y79 = n184 ;
  assign y80 = n293 ;
  assign y81 = n143 ;
  assign y82 = n294 ;
  assign y83 = n295 ;
  assign y84 = n80 ;
  assign y85 = n296 ;
  assign y86 = n297 ;
  assign y87 = n298 ;
  assign y88 = n299 ;
  assign y89 = n300 ;
  assign y90 = n301 ;
  assign y91 = n185 ;
  assign y92 = n302 ;
  assign y93 = n186 ;
  assign y94 = n187 ;
  assign y95 = n188 ;
  assign y96 = n303 ;
  assign y97 = n81 ;
  assign y98 = n304 ;
  assign y99 = n305 ;
  assign y100 = n82 ;
  assign y101 = n306 ;
  assign y102 = n307 ;
  assign y103 = n308 ;
  assign y104 = n309 ;
  assign y105 = n310 ;
  assign y106 = n311 ;
  assign y107 = n189 ;
  assign y108 = n312 ;
  assign y109 = n190 ;
  assign y110 = n191 ;
  assign y111 = n192 ;
  assign y112 = n222 ;
  assign y113 = n83 ;
  assign y114 = n223 ;
  assign y115 = n224 ;
  assign y116 = n84 ;
  assign y117 = n225 ;
  assign y118 = n226 ;
  assign y119 = n227 ;
  assign y120 = n228 ;
  assign y121 = n229 ;
  assign y122 = n230 ;
  assign y123 = n193 ;
  assign y124 = n231 ;
  assign y125 = n194 ;
  assign y126 = n195 ;
  assign y127 = n196 ;
  assign y128 = ~n232 ;
  assign y129 = n49 ;
  assign y130 = n233 ;
  assign y131 = n234 ;
  assign y132 = n50 ;
  assign y133 = n235 ;
  assign y134 = n236 ;
  assign y135 = n237 ;
  assign y136 = n238 ;
  assign y137 = n239 ;
  assign y138 = n240 ;
  assign y139 = n197 ;
  assign y140 = n241 ;
  assign y141 = n198 ;
  assign y142 = n199 ;
  assign y143 = n200 ;
  assign y144 = n242 ;
  assign y145 = n52 ;
  assign y146 = n243 ;
  assign y147 = n244 ;
  assign y148 = n85 ;
  assign y149 = n245 ;
  assign y150 = n246 ;
  assign y151 = n247 ;
  assign y152 = n248 ;
  assign y153 = n249 ;
  assign y154 = n250 ;
  assign y155 = n201 ;
  assign y156 = n251 ;
  assign y157 = n202 ;
  assign y158 = n203 ;
  assign y159 = n204 ;
  assign y160 = n252 ;
  assign y161 = n86 ;
  assign y162 = n253 ;
  assign y163 = n254 ;
  assign y164 = n87 ;
  assign y165 = n255 ;
  assign y166 = n256 ;
  assign y167 = n257 ;
  assign y168 = n258 ;
  assign y169 = n259 ;
  assign y170 = n260 ;
  assign y171 = n88 ;
  assign y172 = n261 ;
  assign y173 = n205 ;
  assign y174 = n206 ;
  assign y175 = n207 ;
  assign y176 = n89 ;
  assign y177 = n90 ;
  assign y178 = n91 ;
  assign y179 = n92 ;
  assign y180 = n93 ;
  assign y181 = n94 ;
  assign y182 = n95 ;
  assign y183 = n96 ;
  assign y184 = n97 ;
  assign y185 = n98 ;
  assign y186 = n99 ;
  assign y187 = n100 ;
  assign y188 = n101 ;
  assign y189 = n102 ;
  assign y190 = n103 ;
  assign y191 = n104 ;
  assign y192 = n105 ;
  assign y193 = n106 ;
  assign y194 = n107 ;
  assign y195 = n108 ;
  assign y196 = n109 ;
  assign y197 = n110 ;
  assign y198 = n111 ;
  assign y199 = n112 ;
  assign y200 = n113 ;
  assign y201 = n114 ;
  assign y202 = n115 ;
  assign y203 = n116 ;
  assign y204 = n117 ;
  assign y205 = n118 ;
  assign y206 = n119 ;
  assign y207 = n120 ;
  assign y208 = n121 ;
  assign y209 = n122 ;
  assign y210 = n123 ;
  assign y211 = n124 ;
  assign y212 = n125 ;
  assign y213 = n126 ;
  assign y214 = n127 ;
  assign y215 = n128 ;
  assign y216 = n129 ;
  assign y217 = n130 ;
  assign y218 = n58 ;
  assign y219 = n59 ;
  assign y220 = n60 ;
  assign y221 = n61 ;
  assign y222 = n62 ;
  assign y223 = n63 ;
  assign y224 = n65 ;
  assign y225 = n131 ;
  assign y226 = n66 ;
  assign y227 = n67 ;
  assign y228 = n132 ;
  assign y229 = n70 ;
  assign y230 = n133 ;
  assign y231 = n134 ;
  assign y232 = n135 ;
  assign y233 = n136 ;
  assign y234 = n137 ;
  assign y235 = n138 ;
  assign y236 = n139 ;
  assign y237 = n140 ;
  assign y238 = n141 ;
  assign y239 = n142 ;
  assign y240 = n208 ;
  assign y241 = n144 ;
  assign y242 = n210 ;
  assign y243 = n211 ;
  assign y244 = n145 ;
  assign y245 = n212 ;
  assign y246 = n213 ;
  assign y247 = n214 ;
  assign y248 = n215 ;
  assign y249 = n216 ;
  assign y250 = n217 ;
  assign y251 = n218 ;
  assign y252 = n262 ;
  assign y253 = n219 ;
  assign y254 = n220 ;
  assign y255 = n221 ;
endmodule
