module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 ;
  wire n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 ;
  assign n513 = x0 & ~x128 ;
  assign n514 = ( x1 & ~x129 ) | ( x1 & n513 ) | ( ~x129 & n513 ) ;
  assign n515 = ~x35 & x163 ;
  assign n516 = ~x33 & x161 ;
  assign n517 = ~x34 & x162 ;
  assign n518 = ( n515 & ~n516 ) | ( n515 & n517 ) | ( ~n516 & n517 ) ;
  assign n519 = x38 & x166 ;
  assign n520 = ~x39 & x167 ;
  assign n521 = ( x166 & ~n519 ) | ( x166 & n520 ) | ( ~n519 & n520 ) ;
  assign n522 = ( x2 & ~x130 ) | ( x2 & n514 ) | ( ~x130 & n514 ) ;
  assign n523 = ( x3 & ~x131 ) | ( x3 & n522 ) | ( ~x131 & n522 ) ;
  assign n524 = ( x4 & ~x132 ) | ( x4 & n523 ) | ( ~x132 & n523 ) ;
  assign n525 = ( x5 & ~x133 ) | ( x5 & n524 ) | ( ~x133 & n524 ) ;
  assign n526 = ( x6 & ~x134 ) | ( x6 & n525 ) | ( ~x134 & n525 ) ;
  assign n527 = ( x7 & ~x135 ) | ( x7 & n526 ) | ( ~x135 & n526 ) ;
  assign n528 = ( x8 & ~x136 ) | ( x8 & n527 ) | ( ~x136 & n527 ) ;
  assign n529 = ( x9 & ~x137 ) | ( x9 & n528 ) | ( ~x137 & n528 ) ;
  assign n530 = ( x10 & ~x138 ) | ( x10 & n529 ) | ( ~x138 & n529 ) ;
  assign n531 = ( x11 & ~x139 ) | ( x11 & n530 ) | ( ~x139 & n530 ) ;
  assign n532 = ( x12 & ~x140 ) | ( x12 & n531 ) | ( ~x140 & n531 ) ;
  assign n533 = ( n516 & n518 ) | ( n516 & ~n521 ) | ( n518 & ~n521 ) ;
  assign n534 = ~x36 & x164 ;
  assign n535 = ( x13 & ~x141 ) | ( x13 & n532 ) | ( ~x141 & n532 ) ;
  assign n536 = ( x14 & ~x142 ) | ( x14 & n535 ) | ( ~x142 & n535 ) ;
  assign n537 = ( x15 & ~x143 ) | ( x15 & n536 ) | ( ~x143 & n536 ) ;
  assign n538 = ( x16 & ~x144 ) | ( x16 & n537 ) | ( ~x144 & n537 ) ;
  assign n539 = ( x17 & ~x145 ) | ( x17 & n538 ) | ( ~x145 & n538 ) ;
  assign n540 = ( x18 & ~x146 ) | ( x18 & n539 ) | ( ~x146 & n539 ) ;
  assign n541 = ( x19 & ~x147 ) | ( x19 & n540 ) | ( ~x147 & n540 ) ;
  assign n542 = ( x20 & ~x148 ) | ( x20 & n541 ) | ( ~x148 & n541 ) ;
  assign n543 = ( x21 & ~x149 ) | ( x21 & n542 ) | ( ~x149 & n542 ) ;
  assign n544 = ( x22 & ~x150 ) | ( x22 & n543 ) | ( ~x150 & n543 ) ;
  assign n545 = ( x23 & ~x151 ) | ( x23 & n544 ) | ( ~x151 & n544 ) ;
  assign n546 = ( x24 & ~x152 ) | ( x24 & n545 ) | ( ~x152 & n545 ) ;
  assign n547 = ( x25 & ~x153 ) | ( x25 & n546 ) | ( ~x153 & n546 ) ;
  assign n548 = ( x26 & ~x154 ) | ( x26 & n547 ) | ( ~x154 & n547 ) ;
  assign n549 = ( x27 & ~x155 ) | ( x27 & n548 ) | ( ~x155 & n548 ) ;
  assign n550 = ( x28 & ~x156 ) | ( x28 & n549 ) | ( ~x156 & n549 ) ;
  assign n551 = ( x29 & ~x157 ) | ( x29 & n550 ) | ( ~x157 & n550 ) ;
  assign n552 = ( x30 & ~x158 ) | ( x30 & n551 ) | ( ~x158 & n551 ) ;
  assign n553 = ( x31 & ~x159 ) | ( x31 & n552 ) | ( ~x159 & n552 ) ;
  assign n554 = ~n533 & n553 ;
  assign n555 = ~x37 & x165 ;
  assign n556 = ( ~n521 & n534 ) | ( ~n521 & n555 ) | ( n534 & n555 ) ;
  assign n557 = x32 & x160 ;
  assign n558 = ( ~n521 & n554 ) | ( ~n521 & n556 ) | ( n554 & n556 ) ;
  assign n559 = ~n556 & n558 ;
  assign n560 = ( ~x160 & n557 ) | ( ~x160 & n559 ) | ( n557 & n559 ) ;
  assign n561 = n521 | n556 ;
  assign n562 = x36 & ~x164 ;
  assign n563 = ( x37 & ~x165 ) | ( x37 & n562 ) | ( ~x165 & n562 ) ;
  assign n564 = x32 & ~x160 ;
  assign n565 = ( x33 & ~x161 ) | ( x33 & n564 ) | ( ~x161 & n564 ) ;
  assign n566 = ( x34 & ~x162 ) | ( x34 & n565 ) | ( ~x162 & n565 ) ;
  assign n567 = ( x38 & ~x166 ) | ( x38 & n563 ) | ( ~x166 & n563 ) ;
  assign n568 = ~n520 & n567 ;
  assign n569 = ( x35 & ~x163 ) | ( x35 & n566 ) | ( ~x163 & n566 ) ;
  assign n570 = x39 & ~x167 ;
  assign n571 = n561 & n569 ;
  assign n572 = ( n568 & n569 ) | ( n568 & ~n571 ) | ( n569 & ~n571 ) ;
  assign n573 = x43 & x171 ;
  assign n574 = ~x42 & x170 ;
  assign n575 = ( x171 & ~n573 ) | ( x171 & n574 ) | ( ~n573 & n574 ) ;
  assign n576 = ( ~n560 & n570 ) | ( ~n560 & n572 ) | ( n570 & n572 ) ;
  assign n577 = ~x41 & x169 ;
  assign n578 = ~x40 & x168 ;
  assign n579 = ( ~n575 & n577 ) | ( ~n575 & n578 ) | ( n577 & n578 ) ;
  assign n580 = ~x47 & x175 ;
  assign n581 = n560 | n576 ;
  assign n582 = x46 & x174 ;
  assign n583 = ( x174 & n580 ) | ( x174 & ~n582 ) | ( n580 & ~n582 ) ;
  assign n584 = ( n575 & n579 ) | ( n575 & ~n583 ) | ( n579 & ~n583 ) ;
  assign n585 = n581 & ~n584 ;
  assign n586 = ~x45 & x173 ;
  assign n587 = ~x44 & x172 ;
  assign n588 = ( ~n583 & n586 ) | ( ~n583 & n587 ) | ( n586 & n587 ) ;
  assign n589 = ( ~n583 & n585 ) | ( ~n583 & n588 ) | ( n585 & n588 ) ;
  assign n590 = ~n588 & n589 ;
  assign n591 = x40 & ~x168 ;
  assign n592 = ( x41 & ~x169 ) | ( x41 & n591 ) | ( ~x169 & n591 ) ;
  assign n593 = ( x42 & ~x170 ) | ( x42 & n592 ) | ( ~x170 & n592 ) ;
  assign n594 = ( x43 & ~x171 ) | ( x43 & n593 ) | ( ~x171 & n593 ) ;
  assign n595 = ( ~n583 & n588 ) | ( ~n583 & n594 ) | ( n588 & n594 ) ;
  assign n596 = x44 & ~x172 ;
  assign n597 = ( x45 & ~x173 ) | ( x45 & n596 ) | ( ~x173 & n596 ) ;
  assign n598 = ( x46 & ~x174 ) | ( x46 & n597 ) | ( ~x174 & n597 ) ;
  assign n599 = ~n588 & n595 ;
  assign n600 = x80 & ~x208 ;
  assign n601 = n580 & n598 ;
  assign n602 = ( n590 & n598 ) | ( n590 & ~n601 ) | ( n598 & ~n601 ) ;
  assign n603 = x47 & ~x175 ;
  assign n604 = ( n599 & ~n602 ) | ( n599 & n603 ) | ( ~n602 & n603 ) ;
  assign n605 = n602 | n604 ;
  assign n606 = x55 & x183 ;
  assign n607 = ~x54 & x182 ;
  assign n608 = ~x50 & x178 ;
  assign n609 = ( x183 & ~n606 ) | ( x183 & n607 ) | ( ~n606 & n607 ) ;
  assign n610 = ~x52 & x180 ;
  assign n611 = ~x53 & x181 ;
  assign n612 = ~x51 & x179 ;
  assign n613 = ( ~n609 & n610 ) | ( ~n609 & n611 ) | ( n610 & n611 ) ;
  assign n614 = ~x49 & x177 ;
  assign n615 = ( n608 & n612 ) | ( n608 & ~n614 ) | ( n612 & ~n614 ) ;
  assign n616 = ( ~n609 & n614 ) | ( ~n609 & n615 ) | ( n614 & n615 ) ;
  assign n617 = ~x63 & x191 ;
  assign n618 = ( ~n609 & n613 ) | ( ~n609 & n616 ) | ( n613 & n616 ) ;
  assign n619 = ( x81 & ~x209 ) | ( x81 & n600 ) | ( ~x209 & n600 ) ;
  assign n620 = x48 & x176 ;
  assign n621 = n609 | n618 ;
  assign n622 = ( x176 & ~n620 ) | ( x176 & n621 ) | ( ~n620 & n621 ) ;
  assign n623 = n605 & ~n622 ;
  assign n624 = ~x60 & x188 ;
  assign n625 = x62 & x190 ;
  assign n626 = ( x190 & n617 ) | ( x190 & ~n625 ) | ( n617 & ~n625 ) ;
  assign n627 = ( x82 & ~x210 ) | ( x82 & n619 ) | ( ~x210 & n619 ) ;
  assign n628 = ( x83 & ~x211 ) | ( x83 & n627 ) | ( ~x211 & n627 ) ;
  assign n629 = n609 | n613 ;
  assign n630 = ~x61 & x189 ;
  assign n631 = ( ~n624 & n626 ) | ( ~n624 & n630 ) | ( n626 & n630 ) ;
  assign n632 = n624 | n631 ;
  assign n633 = x48 & ~x176 ;
  assign n634 = ( x49 & ~x177 ) | ( x49 & n633 ) | ( ~x177 & n633 ) ;
  assign n635 = ( x50 & ~x178 ) | ( x50 & n634 ) | ( ~x178 & n634 ) ;
  assign n636 = ( x51 & ~x179 ) | ( x51 & n635 ) | ( ~x179 & n635 ) ;
  assign n637 = x55 & ~x183 ;
  assign n638 = ( ~n629 & n636 ) | ( ~n629 & n637 ) | ( n636 & n637 ) ;
  assign n639 = x56 & ~x184 ;
  assign n640 = x52 & ~x180 ;
  assign n641 = ( x53 & ~x181 ) | ( x53 & n640 ) | ( ~x181 & n640 ) ;
  assign n642 = ( x54 & ~x182 ) | ( x54 & n641 ) | ( ~x182 & n641 ) ;
  assign n643 = ( x55 & ~x183 ) | ( x55 & n642 ) | ( ~x183 & n642 ) ;
  assign n644 = ( x57 & ~x185 ) | ( x57 & n639 ) | ( ~x185 & n639 ) ;
  assign n645 = ( x58 & ~x186 ) | ( x58 & n644 ) | ( ~x186 & n644 ) ;
  assign n646 = ( x59 & ~x187 ) | ( x59 & n645 ) | ( ~x187 & n645 ) ;
  assign n647 = ( ~n623 & n638 ) | ( ~n623 & n643 ) | ( n638 & n643 ) ;
  assign n648 = ( ~x57 & x185 ) | ( ~x57 & n632 ) | ( x185 & n632 ) ;
  assign n649 = n623 | n647 ;
  assign n650 = x56 & x184 ;
  assign n651 = ~n632 & n646 ;
  assign n652 = ( x184 & n632 ) | ( x184 & ~n650 ) | ( n632 & ~n650 ) ;
  assign n653 = ~x59 & x187 ;
  assign n654 = n648 | n652 ;
  assign n655 = ~x58 & x186 ;
  assign n656 = ( ~n653 & n654 ) | ( ~n653 & n655 ) | ( n654 & n655 ) ;
  assign n657 = ( n649 & ~n653 ) | ( n649 & n656 ) | ( ~n653 & n656 ) ;
  assign n658 = x60 & ~x188 ;
  assign n659 = ( x61 & ~x189 ) | ( x61 & n658 ) | ( ~x189 & n658 ) ;
  assign n660 = ( x62 & ~x190 ) | ( x62 & n659 ) | ( ~x190 & n659 ) ;
  assign n661 = ~n656 & n657 ;
  assign n662 = x63 & ~x191 ;
  assign n663 = n617 & n660 ;
  assign n664 = ( n660 & n661 ) | ( n660 & ~n663 ) | ( n661 & ~n663 ) ;
  assign n665 = ( n651 & n662 ) | ( n651 & ~n664 ) | ( n662 & ~n664 ) ;
  assign n666 = n664 | n665 ;
  assign n667 = ( x64 & ~x192 ) | ( x64 & n666 ) | ( ~x192 & n666 ) ;
  assign n668 = x71 & x199 ;
  assign n669 = ~x70 & x198 ;
  assign n670 = ( x65 & ~x193 ) | ( x65 & n667 ) | ( ~x193 & n667 ) ;
  assign n671 = ( x66 & ~x194 ) | ( x66 & n670 ) | ( ~x194 & n670 ) ;
  assign n672 = ( x199 & ~n668 ) | ( x199 & n669 ) | ( ~n668 & n669 ) ;
  assign n673 = ~x69 & x197 ;
  assign n674 = ( x67 & ~x195 ) | ( x67 & n671 ) | ( ~x195 & n671 ) ;
  assign n675 = ~x68 & x196 ;
  assign n676 = ( ~n672 & n673 ) | ( ~n672 & n675 ) | ( n673 & n675 ) ;
  assign n677 = n674 & ~n676 ;
  assign n678 = n672 & n677 ;
  assign n679 = x68 & ~x196 ;
  assign n680 = ( x69 & ~x197 ) | ( x69 & n679 ) | ( ~x197 & n679 ) ;
  assign n681 = ( x70 & ~x198 ) | ( x70 & n680 ) | ( ~x198 & n680 ) ;
  assign n682 = ( x71 & ~x199 ) | ( x71 & n681 ) | ( ~x199 & n681 ) ;
  assign n683 = ( n677 & ~n678 ) | ( n677 & n682 ) | ( ~n678 & n682 ) ;
  assign n684 = ~x74 & x202 ;
  assign n685 = x75 & x203 ;
  assign n686 = ( x203 & n684 ) | ( x203 & ~n685 ) | ( n684 & ~n685 ) ;
  assign n687 = ~x72 & x200 ;
  assign n688 = ~x73 & x201 ;
  assign n689 = ( ~n686 & n687 ) | ( ~n686 & n688 ) | ( n687 & n688 ) ;
  assign n690 = x72 & ~x200 ;
  assign n691 = ( x73 & ~x201 ) | ( x73 & n690 ) | ( ~x201 & n690 ) ;
  assign n692 = ( x74 & ~x202 ) | ( x74 & n691 ) | ( ~x202 & n691 ) ;
  assign n693 = ( n683 & ~n686 ) | ( n683 & n689 ) | ( ~n686 & n689 ) ;
  assign n694 = n689 & n693 ;
  assign n695 = ( x75 & ~x203 ) | ( x75 & n692 ) | ( ~x203 & n692 ) ;
  assign n696 = x79 & x207 ;
  assign n697 = ( n693 & ~n694 ) | ( n693 & n695 ) | ( ~n694 & n695 ) ;
  assign n698 = ~x76 & x204 ;
  assign n699 = ~x78 & x206 ;
  assign n700 = ( x207 & ~n696 ) | ( x207 & n699 ) | ( ~n696 & n699 ) ;
  assign n701 = ~x77 & x205 ;
  assign n702 = ( n698 & ~n700 ) | ( n698 & n701 ) | ( ~n700 & n701 ) ;
  assign n703 = n697 & ~n702 ;
  assign n704 = n700 & n703 ;
  assign n705 = x76 & ~x204 ;
  assign n706 = ( x77 & ~x205 ) | ( x77 & n705 ) | ( ~x205 & n705 ) ;
  assign n707 = ( x78 & ~x206 ) | ( x78 & n706 ) | ( ~x206 & n706 ) ;
  assign n708 = ( x79 & ~x207 ) | ( x79 & n707 ) | ( ~x207 & n707 ) ;
  assign n709 = ( n703 & ~n704 ) | ( n703 & n708 ) | ( ~n704 & n708 ) ;
  assign n710 = ~x81 & x209 ;
  assign n711 = x82 & x210 ;
  assign n712 = ( ~x83 & x211 ) | ( ~x83 & n710 ) | ( x211 & n710 ) ;
  assign n713 = ( x210 & n710 ) | ( x210 & ~n711 ) | ( n710 & ~n711 ) ;
  assign n714 = n709 & ~n713 ;
  assign n715 = ~n712 & n714 ;
  assign n716 = x80 & x208 ;
  assign n717 = ( ~x208 & n715 ) | ( ~x208 & n716 ) | ( n715 & n716 ) ;
  assign n718 = n628 | n717 ;
  assign n719 = ~x85 & x213 ;
  assign n720 = ~x86 & x214 ;
  assign n721 = x87 & x215 ;
  assign n722 = ( x215 & n720 ) | ( x215 & ~n721 ) | ( n720 & ~n721 ) ;
  assign n723 = ~x84 & x212 ;
  assign n724 = ( n719 & ~n722 ) | ( n719 & n723 ) | ( ~n722 & n723 ) ;
  assign n725 = n718 & ~n724 ;
  assign n726 = x91 & x219 ;
  assign n727 = x84 & ~x212 ;
  assign n728 = ( x85 & ~x213 ) | ( x85 & n727 ) | ( ~x213 & n727 ) ;
  assign n729 = ( x86 & ~x214 ) | ( x86 & n728 ) | ( ~x214 & n728 ) ;
  assign n730 = ( x87 & ~x215 ) | ( x87 & n729 ) | ( ~x215 & n729 ) ;
  assign n731 = n722 & n725 ;
  assign n732 = ( n725 & n730 ) | ( n725 & ~n731 ) | ( n730 & ~n731 ) ;
  assign n733 = ~x89 & x217 ;
  assign n734 = ~x90 & x218 ;
  assign n735 = ( x219 & ~n726 ) | ( x219 & n734 ) | ( ~n726 & n734 ) ;
  assign n736 = ~x88 & x216 ;
  assign n737 = ( n733 & ~n735 ) | ( n733 & n736 ) | ( ~n735 & n736 ) ;
  assign n738 = ( n732 & ~n735 ) | ( n732 & n737 ) | ( ~n735 & n737 ) ;
  assign n739 = x88 & ~x216 ;
  assign n740 = ( x89 & ~x217 ) | ( x89 & n739 ) | ( ~x217 & n739 ) ;
  assign n741 = ( x90 & ~x218 ) | ( x90 & n740 ) | ( ~x218 & n740 ) ;
  assign n742 = ( x91 & ~x219 ) | ( x91 & n741 ) | ( ~x219 & n741 ) ;
  assign n743 = n737 & n738 ;
  assign n744 = x95 & x223 ;
  assign n745 = ( n738 & n742 ) | ( n738 & ~n743 ) | ( n742 & ~n743 ) ;
  assign n746 = ~x94 & x222 ;
  assign n747 = ~x92 & x220 ;
  assign n748 = ( x223 & ~n744 ) | ( x223 & n746 ) | ( ~n744 & n746 ) ;
  assign n749 = ~x93 & x221 ;
  assign n750 = ( n747 & ~n748 ) | ( n747 & n749 ) | ( ~n748 & n749 ) ;
  assign n751 = x96 & x224 ;
  assign n752 = n745 & ~n750 ;
  assign n753 = x92 & ~x220 ;
  assign n754 = n748 & n752 ;
  assign n755 = ( x93 & ~x221 ) | ( x93 & n753 ) | ( ~x221 & n753 ) ;
  assign n756 = ( x94 & ~x222 ) | ( x94 & n755 ) | ( ~x222 & n755 ) ;
  assign n757 = ( x95 & ~x223 ) | ( x95 & n756 ) | ( ~x223 & n756 ) ;
  assign n758 = ( n752 & ~n754 ) | ( n752 & n757 ) | ( ~n754 & n757 ) ;
  assign n759 = ~x97 & x225 ;
  assign n760 = x98 & x226 ;
  assign n761 = ( x226 & n759 ) | ( x226 & ~n760 ) | ( n759 & ~n760 ) ;
  assign n762 = ( ~x99 & x227 ) | ( ~x99 & n759 ) | ( x227 & n759 ) ;
  assign n763 = n758 & ~n761 ;
  assign n764 = x96 & ~x224 ;
  assign n765 = ( x97 & ~x225 ) | ( x97 & n764 ) | ( ~x225 & n764 ) ;
  assign n766 = ( x98 & ~x226 ) | ( x98 & n765 ) | ( ~x226 & n765 ) ;
  assign n767 = ( x99 & ~x227 ) | ( x99 & n766 ) | ( ~x227 & n766 ) ;
  assign n768 = ~n762 & n763 ;
  assign n769 = ( ~x224 & n751 ) | ( ~x224 & n768 ) | ( n751 & n768 ) ;
  assign n770 = n767 | n769 ;
  assign n771 = ~x101 & x229 ;
  assign n772 = ~x102 & x230 ;
  assign n773 = x103 & x231 ;
  assign n774 = ( x231 & n772 ) | ( x231 & ~n773 ) | ( n772 & ~n773 ) ;
  assign n775 = ~x100 & x228 ;
  assign n776 = ( n771 & ~n774 ) | ( n771 & n775 ) | ( ~n774 & n775 ) ;
  assign n777 = n770 & ~n776 ;
  assign n778 = x107 & x235 ;
  assign n779 = x100 & ~x228 ;
  assign n780 = ( x101 & ~x229 ) | ( x101 & n779 ) | ( ~x229 & n779 ) ;
  assign n781 = ( x102 & ~x230 ) | ( x102 & n780 ) | ( ~x230 & n780 ) ;
  assign n782 = ( x103 & ~x231 ) | ( x103 & n781 ) | ( ~x231 & n781 ) ;
  assign n783 = n774 & n777 ;
  assign n784 = ( n777 & n782 ) | ( n777 & ~n783 ) | ( n782 & ~n783 ) ;
  assign n785 = ~x105 & x233 ;
  assign n786 = ~x106 & x234 ;
  assign n787 = ( x235 & ~n778 ) | ( x235 & n786 ) | ( ~n778 & n786 ) ;
  assign n788 = ~x104 & x232 ;
  assign n789 = ( n785 & ~n787 ) | ( n785 & n788 ) | ( ~n787 & n788 ) ;
  assign n790 = ( n784 & ~n787 ) | ( n784 & n789 ) | ( ~n787 & n789 ) ;
  assign n791 = x104 & ~x232 ;
  assign n792 = ( x105 & ~x233 ) | ( x105 & n791 ) | ( ~x233 & n791 ) ;
  assign n793 = ( x106 & ~x234 ) | ( x106 & n792 ) | ( ~x234 & n792 ) ;
  assign n794 = ( x107 & ~x235 ) | ( x107 & n793 ) | ( ~x235 & n793 ) ;
  assign n795 = n789 & n790 ;
  assign n796 = x111 & x239 ;
  assign n797 = ( n790 & n794 ) | ( n790 & ~n795 ) | ( n794 & ~n795 ) ;
  assign n798 = ~x110 & x238 ;
  assign n799 = ~x108 & x236 ;
  assign n800 = ( x239 & ~n796 ) | ( x239 & n798 ) | ( ~n796 & n798 ) ;
  assign n801 = ~x109 & x237 ;
  assign n802 = ( n799 & ~n800 ) | ( n799 & n801 ) | ( ~n800 & n801 ) ;
  assign n803 = x112 & x240 ;
  assign n804 = n797 & ~n802 ;
  assign n805 = x108 & ~x236 ;
  assign n806 = n800 & n804 ;
  assign n807 = ( x109 & ~x237 ) | ( x109 & n805 ) | ( ~x237 & n805 ) ;
  assign n808 = ( x110 & ~x238 ) | ( x110 & n807 ) | ( ~x238 & n807 ) ;
  assign n809 = ( x111 & ~x239 ) | ( x111 & n808 ) | ( ~x239 & n808 ) ;
  assign n810 = ( n804 & ~n806 ) | ( n804 & n809 ) | ( ~n806 & n809 ) ;
  assign n811 = ~x113 & x241 ;
  assign n812 = x114 & x242 ;
  assign n813 = ( x242 & n811 ) | ( x242 & ~n812 ) | ( n811 & ~n812 ) ;
  assign n814 = ( ~x115 & x243 ) | ( ~x115 & n811 ) | ( x243 & n811 ) ;
  assign n815 = n810 & ~n813 ;
  assign n816 = x112 & ~x240 ;
  assign n817 = ( x113 & ~x241 ) | ( x113 & n816 ) | ( ~x241 & n816 ) ;
  assign n818 = ( x114 & ~x242 ) | ( x114 & n817 ) | ( ~x242 & n817 ) ;
  assign n819 = ( x115 & ~x243 ) | ( x115 & n818 ) | ( ~x243 & n818 ) ;
  assign n820 = ~n814 & n815 ;
  assign n821 = ( ~x240 & n803 ) | ( ~x240 & n820 ) | ( n803 & n820 ) ;
  assign n822 = n819 | n821 ;
  assign n823 = x119 & x247 ;
  assign n824 = ~x117 & x245 ;
  assign n825 = ~x118 & x246 ;
  assign n826 = ( x247 & ~n823 ) | ( x247 & n825 ) | ( ~n823 & n825 ) ;
  assign n827 = ~x116 & x244 ;
  assign n828 = ( n824 & ~n826 ) | ( n824 & n827 ) | ( ~n826 & n827 ) ;
  assign n829 = ~x122 & x250 ;
  assign n830 = n822 & ~n828 ;
  assign n831 = x123 & x251 ;
  assign n832 = ( x251 & n829 ) | ( x251 & ~n831 ) | ( n829 & ~n831 ) ;
  assign n833 = n826 & n830 ;
  assign n834 = x116 & ~x244 ;
  assign n835 = ( x117 & ~x245 ) | ( x117 & n834 ) | ( ~x245 & n834 ) ;
  assign n836 = ( x118 & ~x246 ) | ( x118 & n835 ) | ( ~x246 & n835 ) ;
  assign n837 = ( x119 & ~x247 ) | ( x119 & n836 ) | ( ~x247 & n836 ) ;
  assign n838 = ( n830 & ~n833 ) | ( n830 & n837 ) | ( ~n833 & n837 ) ;
  assign n839 = ~x120 & x248 ;
  assign n840 = ~x121 & x249 ;
  assign n841 = ( ~n832 & n839 ) | ( ~n832 & n840 ) | ( n839 & n840 ) ;
  assign n842 = x256 & ~x384 ;
  assign n843 = ( x257 & ~x385 ) | ( x257 & n842 ) | ( ~x385 & n842 ) ;
  assign n844 = ( x258 & ~x386 ) | ( x258 & n843 ) | ( ~x386 & n843 ) ;
  assign n845 = ( x259 & ~x387 ) | ( x259 & n844 ) | ( ~x387 & n844 ) ;
  assign n846 = ( ~n832 & n838 ) | ( ~n832 & n841 ) | ( n838 & n841 ) ;
  assign n847 = x120 & ~x248 ;
  assign n848 = ( x260 & ~x388 ) | ( x260 & n845 ) | ( ~x388 & n845 ) ;
  assign n849 = ( x261 & ~x389 ) | ( x261 & n848 ) | ( ~x389 & n848 ) ;
  assign n850 = ( x262 & ~x390 ) | ( x262 & n849 ) | ( ~x390 & n849 ) ;
  assign n851 = ( x263 & ~x391 ) | ( x263 & n850 ) | ( ~x391 & n850 ) ;
  assign n852 = ( x264 & ~x392 ) | ( x264 & n851 ) | ( ~x392 & n851 ) ;
  assign n853 = ( x265 & ~x393 ) | ( x265 & n852 ) | ( ~x393 & n852 ) ;
  assign n854 = n841 & n846 ;
  assign n855 = ( x266 & ~x394 ) | ( x266 & n853 ) | ( ~x394 & n853 ) ;
  assign n856 = ( x267 & ~x395 ) | ( x267 & n855 ) | ( ~x395 & n855 ) ;
  assign n857 = ( x268 & ~x396 ) | ( x268 & n856 ) | ( ~x396 & n856 ) ;
  assign n858 = ( x269 & ~x397 ) | ( x269 & n857 ) | ( ~x397 & n857 ) ;
  assign n859 = ( x270 & ~x398 ) | ( x270 & n858 ) | ( ~x398 & n858 ) ;
  assign n860 = ( x271 & ~x399 ) | ( x271 & n859 ) | ( ~x399 & n859 ) ;
  assign n861 = ( x272 & ~x400 ) | ( x272 & n860 ) | ( ~x400 & n860 ) ;
  assign n862 = ( x121 & ~x249 ) | ( x121 & n847 ) | ( ~x249 & n847 ) ;
  assign n863 = ( x122 & ~x250 ) | ( x122 & n862 ) | ( ~x250 & n862 ) ;
  assign n864 = ( x123 & ~x251 ) | ( x123 & n863 ) | ( ~x251 & n863 ) ;
  assign n865 = ( n846 & ~n854 ) | ( n846 & n864 ) | ( ~n854 & n864 ) ;
  assign n866 = ( x273 & ~x401 ) | ( x273 & n861 ) | ( ~x401 & n861 ) ;
  assign n867 = ~x289 & x417 ;
  assign n868 = ~x295 & x423 ;
  assign n869 = ~x290 & x418 ;
  assign n870 = ~x291 & x419 ;
  assign n871 = ( ~n867 & n869 ) | ( ~n867 & n870 ) | ( n869 & n870 ) ;
  assign n872 = x294 & x422 ;
  assign n873 = ( x274 & ~x402 ) | ( x274 & n866 ) | ( ~x402 & n866 ) ;
  assign n874 = ( x275 & ~x403 ) | ( x275 & n873 ) | ( ~x403 & n873 ) ;
  assign n875 = ( x276 & ~x404 ) | ( x276 & n874 ) | ( ~x404 & n874 ) ;
  assign n876 = ( x277 & ~x405 ) | ( x277 & n875 ) | ( ~x405 & n875 ) ;
  assign n877 = ( x278 & ~x406 ) | ( x278 & n876 ) | ( ~x406 & n876 ) ;
  assign n878 = ( x279 & ~x407 ) | ( x279 & n877 ) | ( ~x407 & n877 ) ;
  assign n879 = ( x280 & ~x408 ) | ( x280 & n878 ) | ( ~x408 & n878 ) ;
  assign n880 = ( x281 & ~x409 ) | ( x281 & n879 ) | ( ~x409 & n879 ) ;
  assign n881 = ( x282 & ~x410 ) | ( x282 & n880 ) | ( ~x410 & n880 ) ;
  assign n882 = ( x283 & ~x411 ) | ( x283 & n881 ) | ( ~x411 & n881 ) ;
  assign n883 = ( x284 & ~x412 ) | ( x284 & n882 ) | ( ~x412 & n882 ) ;
  assign n884 = ( x422 & n868 ) | ( x422 & ~n872 ) | ( n868 & ~n872 ) ;
  assign n885 = ( x285 & ~x413 ) | ( x285 & n883 ) | ( ~x413 & n883 ) ;
  assign n886 = ( n867 & n871 ) | ( n867 & ~n884 ) | ( n871 & ~n884 ) ;
  assign n887 = ~x292 & x420 ;
  assign n888 = ( x286 & ~x414 ) | ( x286 & n885 ) | ( ~x414 & n885 ) ;
  assign n889 = ( x287 & ~x415 ) | ( x287 & n888 ) | ( ~x415 & n888 ) ;
  assign n890 = ~n886 & n889 ;
  assign n891 = ~x293 & x421 ;
  assign n892 = ( ~n884 & n887 ) | ( ~n884 & n891 ) | ( n887 & n891 ) ;
  assign n893 = n884 | n892 ;
  assign n894 = ( ~n884 & n890 ) | ( ~n884 & n892 ) | ( n890 & n892 ) ;
  assign n895 = ~n892 & n894 ;
  assign n896 = x288 & x416 ;
  assign n897 = ( ~x416 & n895 ) | ( ~x416 & n896 ) | ( n895 & n896 ) ;
  assign n898 = x288 & ~x416 ;
  assign n899 = ( x289 & ~x417 ) | ( x289 & n898 ) | ( ~x417 & n898 ) ;
  assign n900 = x292 & ~x420 ;
  assign n901 = ( x293 & ~x421 ) | ( x293 & n900 ) | ( ~x421 & n900 ) ;
  assign n902 = ( x294 & ~x422 ) | ( x294 & n901 ) | ( ~x422 & n901 ) ;
  assign n903 = ( x290 & ~x418 ) | ( x290 & n899 ) | ( ~x418 & n899 ) ;
  assign n904 = ( x291 & ~x419 ) | ( x291 & n903 ) | ( ~x419 & n903 ) ;
  assign n905 = n893 & n904 ;
  assign n906 = ~n868 & n902 ;
  assign n907 = ( n904 & ~n905 ) | ( n904 & n906 ) | ( ~n905 & n906 ) ;
  assign n908 = x295 & ~x423 ;
  assign n909 = ( ~n897 & n907 ) | ( ~n897 & n908 ) | ( n907 & n908 ) ;
  assign n910 = n897 | n909 ;
  assign n911 = ~x298 & x426 ;
  assign n912 = ~x296 & x424 ;
  assign n913 = x299 & x427 ;
  assign n914 = ( x427 & n911 ) | ( x427 & ~n913 ) | ( n911 & ~n913 ) ;
  assign n915 = ~x297 & x425 ;
  assign n916 = ~x303 & x431 ;
  assign n917 = ( n912 & ~n914 ) | ( n912 & n915 ) | ( ~n914 & n915 ) ;
  assign n918 = x302 & x430 ;
  assign n919 = ( x430 & n916 ) | ( x430 & ~n918 ) | ( n916 & ~n918 ) ;
  assign n920 = ( n914 & n917 ) | ( n914 & ~n919 ) | ( n917 & ~n919 ) ;
  assign n921 = n910 & ~n920 ;
  assign n922 = ~x301 & x429 ;
  assign n923 = ~x300 & x428 ;
  assign n924 = ( ~n919 & n922 ) | ( ~n919 & n923 ) | ( n922 & n923 ) ;
  assign n925 = ( ~n919 & n921 ) | ( ~n919 & n924 ) | ( n921 & n924 ) ;
  assign n926 = x300 & ~x428 ;
  assign n927 = ( x301 & ~x429 ) | ( x301 & n926 ) | ( ~x429 & n926 ) ;
  assign n928 = ( x302 & ~x430 ) | ( x302 & n927 ) | ( ~x430 & n927 ) ;
  assign n929 = n916 & n928 ;
  assign n930 = ~n924 & n925 ;
  assign n931 = ( n928 & ~n929 ) | ( n928 & n930 ) | ( ~n929 & n930 ) ;
  assign n932 = x296 & ~x424 ;
  assign n933 = ( x297 & ~x425 ) | ( x297 & n932 ) | ( ~x425 & n932 ) ;
  assign n934 = ( x298 & ~x426 ) | ( x298 & n933 ) | ( ~x426 & n933 ) ;
  assign n935 = ( x299 & ~x427 ) | ( x299 & n934 ) | ( ~x427 & n934 ) ;
  assign n936 = ( ~n919 & n924 ) | ( ~n919 & n935 ) | ( n924 & n935 ) ;
  assign n937 = ~n924 & n936 ;
  assign n938 = ~x305 & x433 ;
  assign n939 = ~x306 & x434 ;
  assign n940 = ~x307 & x435 ;
  assign n941 = ( ~n938 & n939 ) | ( ~n938 & n940 ) | ( n939 & n940 ) ;
  assign n942 = x303 & ~x431 ;
  assign n943 = ( ~n931 & n937 ) | ( ~n931 & n942 ) | ( n937 & n942 ) ;
  assign n944 = x311 & x439 ;
  assign n945 = n931 | n943 ;
  assign n946 = ~x310 & x438 ;
  assign n947 = ( x439 & ~n944 ) | ( x439 & n946 ) | ( ~n944 & n946 ) ;
  assign n948 = ( n938 & n941 ) | ( n938 & ~n947 ) | ( n941 & ~n947 ) ;
  assign n949 = ~x308 & x436 ;
  assign n950 = ~x309 & x437 ;
  assign n951 = ( ~n947 & n949 ) | ( ~n947 & n950 ) | ( n949 & n950 ) ;
  assign n952 = x304 & ~x432 ;
  assign n953 = ( x305 & ~x433 ) | ( x305 & n952 ) | ( ~x433 & n952 ) ;
  assign n954 = ( x306 & ~x434 ) | ( x306 & n953 ) | ( ~x434 & n953 ) ;
  assign n955 = ( x307 & ~x435 ) | ( x307 & n954 ) | ( ~x435 & n954 ) ;
  assign n956 = ( ~n947 & n948 ) | ( ~n947 & n951 ) | ( n948 & n951 ) ;
  assign n957 = n947 | n956 ;
  assign n958 = n947 | n951 ;
  assign n959 = x304 & x432 ;
  assign n960 = ( x432 & n957 ) | ( x432 & ~n959 ) | ( n957 & ~n959 ) ;
  assign n961 = x308 & ~x436 ;
  assign n962 = ( x309 & ~x437 ) | ( x309 & n961 ) | ( ~x437 & n961 ) ;
  assign n963 = ( x310 & ~x438 ) | ( x310 & n962 ) | ( ~x438 & n962 ) ;
  assign n964 = n945 & ~n960 ;
  assign n965 = x311 & ~x439 ;
  assign n966 = ( n955 & ~n958 ) | ( n955 & n965 ) | ( ~n958 & n965 ) ;
  assign n967 = ( x311 & ~x439 ) | ( x311 & n963 ) | ( ~x439 & n963 ) ;
  assign n968 = ( ~n964 & n966 ) | ( ~n964 & n967 ) | ( n966 & n967 ) ;
  assign n969 = n964 | n968 ;
  assign n970 = x318 & x446 ;
  assign n971 = ~x316 & x444 ;
  assign n972 = ~x319 & x447 ;
  assign n973 = ( x446 & ~n970 ) | ( x446 & n972 ) | ( ~n970 & n972 ) ;
  assign n974 = ~x317 & x445 ;
  assign n975 = ( ~n971 & n973 ) | ( ~n971 & n974 ) | ( n973 & n974 ) ;
  assign n976 = x312 & x440 ;
  assign n977 = n971 | n975 ;
  assign n978 = ( ~x313 & x441 ) | ( ~x313 & n977 ) | ( x441 & n977 ) ;
  assign n979 = ( x440 & ~n976 ) | ( x440 & n977 ) | ( ~n976 & n977 ) ;
  assign n980 = n978 | n979 ;
  assign n981 = ~x314 & x442 ;
  assign n982 = ~x315 & x443 ;
  assign n983 = ( n980 & n981 ) | ( n980 & ~n982 ) | ( n981 & ~n982 ) ;
  assign n984 = x316 & ~x444 ;
  assign n985 = ( x317 & ~x445 ) | ( x317 & n984 ) | ( ~x445 & n984 ) ;
  assign n986 = ( x318 & ~x446 ) | ( x318 & n985 ) | ( ~x446 & n985 ) ;
  assign n987 = n972 & n986 ;
  assign n988 = ( n969 & ~n982 ) | ( n969 & n983 ) | ( ~n982 & n983 ) ;
  assign n989 = ~n983 & n988 ;
  assign n990 = x331 & x459 ;
  assign n991 = ( n986 & ~n987 ) | ( n986 & n989 ) | ( ~n987 & n989 ) ;
  assign n992 = ~x330 & x458 ;
  assign n993 = ( x459 & ~n990 ) | ( x459 & n992 ) | ( ~n990 & n992 ) ;
  assign n994 = x312 & ~x440 ;
  assign n995 = ( x313 & ~x441 ) | ( x313 & n994 ) | ( ~x441 & n994 ) ;
  assign n996 = ( x314 & ~x442 ) | ( x314 & n995 ) | ( ~x442 & n995 ) ;
  assign n997 = ( x315 & ~x443 ) | ( x315 & n996 ) | ( ~x443 & n996 ) ;
  assign n998 = ~n977 & n997 ;
  assign n999 = ~x328 & x456 ;
  assign n1000 = x319 & ~x447 ;
  assign n1001 = ( ~n991 & n998 ) | ( ~n991 & n1000 ) | ( n998 & n1000 ) ;
  assign n1002 = x327 & x455 ;
  assign n1003 = ~x326 & x454 ;
  assign n1004 = n991 | n1001 ;
  assign n1005 = ( x455 & ~n1002 ) | ( x455 & n1003 ) | ( ~n1002 & n1003 ) ;
  assign n1006 = ~x325 & x453 ;
  assign n1007 = ~x324 & x452 ;
  assign n1008 = ( ~n1005 & n1006 ) | ( ~n1005 & n1007 ) | ( n1006 & n1007 ) ;
  assign n1009 = x328 & ~x456 ;
  assign n1010 = ( x320 & ~x448 ) | ( x320 & n1004 ) | ( ~x448 & n1004 ) ;
  assign n1011 = ( x321 & ~x449 ) | ( x321 & n1010 ) | ( ~x449 & n1010 ) ;
  assign n1012 = ( x329 & ~x457 ) | ( x329 & n1009 ) | ( ~x457 & n1009 ) ;
  assign n1013 = ( x330 & ~x458 ) | ( x330 & n1012 ) | ( ~x458 & n1012 ) ;
  assign n1014 = ( x322 & ~x450 ) | ( x322 & n1011 ) | ( ~x450 & n1011 ) ;
  assign n1015 = ( x323 & ~x451 ) | ( x323 & n1014 ) | ( ~x451 & n1014 ) ;
  assign n1016 = ~n1008 & n1015 ;
  assign n1017 = ~x329 & x457 ;
  assign n1018 = ( ~n993 & n999 ) | ( ~n993 & n1017 ) | ( n999 & n1017 ) ;
  assign n1019 = ( x331 & ~x459 ) | ( x331 & n1013 ) | ( ~x459 & n1013 ) ;
  assign n1020 = x324 & ~x452 ;
  assign n1021 = ( x325 & ~x453 ) | ( x325 & n1020 ) | ( ~x453 & n1020 ) ;
  assign n1022 = ( x326 & ~x454 ) | ( x326 & n1021 ) | ( ~x454 & n1021 ) ;
  assign n1023 = ( x327 & ~x455 ) | ( x327 & n1022 ) | ( ~x455 & n1022 ) ;
  assign n1024 = n1005 & n1016 ;
  assign n1025 = ( n1016 & n1023 ) | ( n1016 & ~n1024 ) | ( n1023 & ~n1024 ) ;
  assign n1026 = ( ~n993 & n1018 ) | ( ~n993 & n1025 ) | ( n1018 & n1025 ) ;
  assign n1027 = n1018 & n1026 ;
  assign n1028 = ( n1019 & n1026 ) | ( n1019 & ~n1027 ) | ( n1026 & ~n1027 ) ;
  assign n1029 = ~x333 & x461 ;
  assign n1030 = x335 & x463 ;
  assign n1031 = ~x334 & x462 ;
  assign n1032 = ( x463 & ~n1030 ) | ( x463 & n1031 ) | ( ~n1030 & n1031 ) ;
  assign n1033 = ~x332 & x460 ;
  assign n1034 = ( n1029 & ~n1032 ) | ( n1029 & n1033 ) | ( ~n1032 & n1033 ) ;
  assign n1035 = n1028 & ~n1034 ;
  assign n1036 = x338 & x466 ;
  assign n1037 = x332 & ~x460 ;
  assign n1038 = ( x333 & ~x461 ) | ( x333 & n1037 ) | ( ~x461 & n1037 ) ;
  assign n1039 = n1032 & n1035 ;
  assign n1040 = ( x334 & ~x462 ) | ( x334 & n1038 ) | ( ~x462 & n1038 ) ;
  assign n1041 = ( x335 & ~x463 ) | ( x335 & n1040 ) | ( ~x463 & n1040 ) ;
  assign n1042 = ( n1035 & ~n1039 ) | ( n1035 & n1041 ) | ( ~n1039 & n1041 ) ;
  assign n1043 = ~x337 & x465 ;
  assign n1044 = ( x466 & ~n1036 ) | ( x466 & n1043 ) | ( ~n1036 & n1043 ) ;
  assign n1045 = n1042 & ~n1044 ;
  assign n1046 = ( ~x339 & x467 ) | ( ~x339 & n1043 ) | ( x467 & n1043 ) ;
  assign n1047 = x336 & ~x464 ;
  assign n1048 = ( x337 & ~x465 ) | ( x337 & n1047 ) | ( ~x465 & n1047 ) ;
  assign n1049 = n1045 & ~n1046 ;
  assign n1050 = ( x338 & ~x466 ) | ( x338 & n1048 ) | ( ~x466 & n1048 ) ;
  assign n1051 = ( x339 & ~x467 ) | ( x339 & n1050 ) | ( ~x467 & n1050 ) ;
  assign n1052 = x336 & x464 ;
  assign n1053 = ( ~x464 & n1049 ) | ( ~x464 & n1052 ) | ( n1049 & n1052 ) ;
  assign n1054 = n1051 | n1053 ;
  assign n1055 = x343 & x471 ;
  assign n1056 = ~x340 & x468 ;
  assign n1057 = ~x342 & x470 ;
  assign n1058 = ( x471 & ~n1055 ) | ( x471 & n1057 ) | ( ~n1055 & n1057 ) ;
  assign n1059 = ~x341 & x469 ;
  assign n1060 = ( n1056 & ~n1058 ) | ( n1056 & n1059 ) | ( ~n1058 & n1059 ) ;
  assign n1061 = ~x346 & x474 ;
  assign n1062 = n1054 & ~n1060 ;
  assign n1063 = x347 & x475 ;
  assign n1064 = ( x475 & n1061 ) | ( x475 & ~n1063 ) | ( n1061 & ~n1063 ) ;
  assign n1065 = x340 & ~x468 ;
  assign n1066 = ( x341 & ~x469 ) | ( x341 & n1065 ) | ( ~x469 & n1065 ) ;
  assign n1067 = ( x342 & ~x470 ) | ( x342 & n1066 ) | ( ~x470 & n1066 ) ;
  assign n1068 = ( x343 & ~x471 ) | ( x343 & n1067 ) | ( ~x471 & n1067 ) ;
  assign n1069 = n1058 & n1062 ;
  assign n1070 = ( n1062 & n1068 ) | ( n1062 & ~n1069 ) | ( n1068 & ~n1069 ) ;
  assign n1071 = ~x345 & x473 ;
  assign n1072 = ~x344 & x472 ;
  assign n1073 = ( ~n1064 & n1071 ) | ( ~n1064 & n1072 ) | ( n1071 & n1072 ) ;
  assign n1074 = x344 & ~x472 ;
  assign n1075 = ( ~n1064 & n1070 ) | ( ~n1064 & n1073 ) | ( n1070 & n1073 ) ;
  assign n1076 = ( x345 & ~x473 ) | ( x345 & n1074 ) | ( ~x473 & n1074 ) ;
  assign n1077 = ( x346 & ~x474 ) | ( x346 & n1076 ) | ( ~x474 & n1076 ) ;
  assign n1078 = ( x347 & ~x475 ) | ( x347 & n1077 ) | ( ~x475 & n1077 ) ;
  assign n1079 = n1073 & n1075 ;
  assign n1080 = ( n1075 & n1078 ) | ( n1075 & ~n1079 ) | ( n1078 & ~n1079 ) ;
  assign n1081 = ~x349 & x477 ;
  assign n1082 = x351 & x479 ;
  assign n1083 = ~x350 & x478 ;
  assign n1084 = ( x479 & ~n1082 ) | ( x479 & n1083 ) | ( ~n1082 & n1083 ) ;
  assign n1085 = ~x348 & x476 ;
  assign n1086 = ( n1081 & ~n1084 ) | ( n1081 & n1085 ) | ( ~n1084 & n1085 ) ;
  assign n1087 = n1080 & ~n1086 ;
  assign n1088 = x354 & x482 ;
  assign n1089 = x348 & ~x476 ;
  assign n1090 = ( x349 & ~x477 ) | ( x349 & n1089 ) | ( ~x477 & n1089 ) ;
  assign n1091 = n1084 & n1087 ;
  assign n1092 = ( x350 & ~x478 ) | ( x350 & n1090 ) | ( ~x478 & n1090 ) ;
  assign n1093 = ( x351 & ~x479 ) | ( x351 & n1092 ) | ( ~x479 & n1092 ) ;
  assign n1094 = ( n1087 & ~n1091 ) | ( n1087 & n1093 ) | ( ~n1091 & n1093 ) ;
  assign n1095 = ~x353 & x481 ;
  assign n1096 = ( x482 & ~n1088 ) | ( x482 & n1095 ) | ( ~n1088 & n1095 ) ;
  assign n1097 = n1094 & ~n1096 ;
  assign n1098 = ( ~x355 & x483 ) | ( ~x355 & n1095 ) | ( x483 & n1095 ) ;
  assign n1099 = x352 & ~x480 ;
  assign n1100 = ( x353 & ~x481 ) | ( x353 & n1099 ) | ( ~x481 & n1099 ) ;
  assign n1101 = n1097 & ~n1098 ;
  assign n1102 = ( x354 & ~x482 ) | ( x354 & n1100 ) | ( ~x482 & n1100 ) ;
  assign n1103 = ( x355 & ~x483 ) | ( x355 & n1102 ) | ( ~x483 & n1102 ) ;
  assign n1104 = x352 & x480 ;
  assign n1105 = ( ~x480 & n1101 ) | ( ~x480 & n1104 ) | ( n1101 & n1104 ) ;
  assign n1106 = n1103 | n1105 ;
  assign n1107 = x359 & x487 ;
  assign n1108 = ~x356 & x484 ;
  assign n1109 = ~x358 & x486 ;
  assign n1110 = ( x487 & ~n1107 ) | ( x487 & n1109 ) | ( ~n1107 & n1109 ) ;
  assign n1111 = ~x357 & x485 ;
  assign n1112 = ( n1108 & ~n1110 ) | ( n1108 & n1111 ) | ( ~n1110 & n1111 ) ;
  assign n1113 = ~x362 & x490 ;
  assign n1114 = n1106 & ~n1112 ;
  assign n1115 = x363 & x491 ;
  assign n1116 = ( x491 & n1113 ) | ( x491 & ~n1115 ) | ( n1113 & ~n1115 ) ;
  assign n1117 = x356 & ~x484 ;
  assign n1118 = ( x357 & ~x485 ) | ( x357 & n1117 ) | ( ~x485 & n1117 ) ;
  assign n1119 = ( x358 & ~x486 ) | ( x358 & n1118 ) | ( ~x486 & n1118 ) ;
  assign n1120 = ( x359 & ~x487 ) | ( x359 & n1119 ) | ( ~x487 & n1119 ) ;
  assign n1121 = n1110 & n1114 ;
  assign n1122 = ( n1114 & n1120 ) | ( n1114 & ~n1121 ) | ( n1120 & ~n1121 ) ;
  assign n1123 = ~x361 & x489 ;
  assign n1124 = ~x360 & x488 ;
  assign n1125 = ( ~n1116 & n1123 ) | ( ~n1116 & n1124 ) | ( n1123 & n1124 ) ;
  assign n1126 = x360 & ~x488 ;
  assign n1127 = ( ~n1116 & n1122 ) | ( ~n1116 & n1125 ) | ( n1122 & n1125 ) ;
  assign n1128 = ( x361 & ~x489 ) | ( x361 & n1126 ) | ( ~x489 & n1126 ) ;
  assign n1129 = ( x362 & ~x490 ) | ( x362 & n1128 ) | ( ~x490 & n1128 ) ;
  assign n1130 = ( x363 & ~x491 ) | ( x363 & n1129 ) | ( ~x491 & n1129 ) ;
  assign n1131 = n1125 & n1127 ;
  assign n1132 = ( n1127 & n1130 ) | ( n1127 & ~n1131 ) | ( n1130 & ~n1131 ) ;
  assign n1133 = ~x366 & x494 ;
  assign n1134 = x367 & x495 ;
  assign n1135 = ( x495 & n1133 ) | ( x495 & ~n1134 ) | ( n1133 & ~n1134 ) ;
  assign n1136 = ~x365 & x493 ;
  assign n1137 = ~x364 & x492 ;
  assign n1138 = ( ~n1135 & n1136 ) | ( ~n1135 & n1137 ) | ( n1136 & n1137 ) ;
  assign n1139 = n1132 & ~n1138 ;
  assign n1140 = x364 & ~x492 ;
  assign n1141 = ( x365 & ~x493 ) | ( x365 & n1140 ) | ( ~x493 & n1140 ) ;
  assign n1142 = n1135 & n1139 ;
  assign n1143 = ( x366 & ~x494 ) | ( x366 & n1141 ) | ( ~x494 & n1141 ) ;
  assign n1144 = ( x367 & ~x495 ) | ( x367 & n1143 ) | ( ~x495 & n1143 ) ;
  assign n1145 = ( n1139 & ~n1142 ) | ( n1139 & n1144 ) | ( ~n1142 & n1144 ) ;
  assign n1146 = x375 & x503 ;
  assign n1147 = ~x374 & x502 ;
  assign n1148 = ( x503 & ~n1146 ) | ( x503 & n1147 ) | ( ~n1146 & n1147 ) ;
  assign n1149 = x370 & x498 ;
  assign n1150 = ~x369 & x497 ;
  assign n1151 = ( x498 & ~n1149 ) | ( x498 & n1150 ) | ( ~n1149 & n1150 ) ;
  assign n1152 = n1145 & ~n1151 ;
  assign n1153 = ( ~x371 & x499 ) | ( ~x371 & n1150 ) | ( x499 & n1150 ) ;
  assign n1154 = n1152 & ~n1153 ;
  assign n1155 = ~x372 & x500 ;
  assign n1156 = ~x373 & x501 ;
  assign n1157 = ( ~n1148 & n1155 ) | ( ~n1148 & n1156 ) | ( n1155 & n1156 ) ;
  assign n1158 = x368 & x496 ;
  assign n1159 = ( ~x496 & n1154 ) | ( ~x496 & n1158 ) | ( n1154 & n1158 ) ;
  assign n1160 = x368 & ~x496 ;
  assign n1161 = ( x369 & ~x497 ) | ( x369 & n1160 ) | ( ~x497 & n1160 ) ;
  assign n1162 = ( x370 & ~x498 ) | ( x370 & n1161 ) | ( ~x498 & n1161 ) ;
  assign n1163 = ( x371 & ~x499 ) | ( x371 & n1162 ) | ( ~x499 & n1162 ) ;
  assign n1164 = n1159 | n1163 ;
  assign n1165 = x372 & ~x500 ;
  assign n1166 = ( x373 & ~x501 ) | ( x373 & n1165 ) | ( ~x501 & n1165 ) ;
  assign n1167 = ( x374 & ~x502 ) | ( x374 & n1166 ) | ( ~x502 & n1166 ) ;
  assign n1168 = ~n1157 & n1164 ;
  assign n1169 = ( x375 & ~x503 ) | ( x375 & n1167 ) | ( ~x503 & n1167 ) ;
  assign n1170 = x379 & x507 ;
  assign n1171 = n1148 & n1168 ;
  assign n1172 = ( n1168 & n1169 ) | ( n1168 & ~n1171 ) | ( n1169 & ~n1171 ) ;
  assign n1173 = ~x378 & x506 ;
  assign n1174 = ( x507 & ~n1170 ) | ( x507 & n1173 ) | ( ~n1170 & n1173 ) ;
  assign n1175 = x376 & ~x504 ;
  assign n1176 = x126 & x254 ;
  assign n1177 = ( x377 & ~x505 ) | ( x377 & n1175 ) | ( ~x505 & n1175 ) ;
  assign n1178 = ~x377 & x505 ;
  assign n1179 = ~x124 & x252 ;
  assign n1180 = ~x376 & x504 ;
  assign n1181 = ( ~n1174 & n1178 ) | ( ~n1174 & n1180 ) | ( n1178 & n1180 ) ;
  assign n1182 = ( n1172 & ~n1174 ) | ( n1172 & n1181 ) | ( ~n1174 & n1181 ) ;
  assign n1183 = n1181 & n1182 ;
  assign n1184 = ( x378 & ~x506 ) | ( x378 & n1177 ) | ( ~x506 & n1177 ) ;
  assign n1185 = x380 & ~x508 ;
  assign n1186 = ( x381 & ~x509 ) | ( x381 & n1185 ) | ( ~x509 & n1185 ) ;
  assign n1187 = ~x381 & x509 ;
  assign n1188 = ( x379 & ~x507 ) | ( x379 & n1184 ) | ( ~x507 & n1184 ) ;
  assign n1189 = ( n1182 & ~n1183 ) | ( n1182 & n1188 ) | ( ~n1183 & n1188 ) ;
  assign n1190 = x382 & x510 ;
  assign n1191 = ~x380 & x508 ;
  assign n1192 = ( x510 & n1187 ) | ( x510 & ~n1190 ) | ( n1187 & ~n1190 ) ;
  assign n1193 = x383 & ~x511 ;
  assign n1194 = ( ~n1191 & n1192 ) | ( ~n1191 & n1193 ) | ( n1192 & n1193 ) ;
  assign n1195 = ~x125 & x253 ;
  assign n1196 = ( x382 & ~x510 ) | ( x382 & n1186 ) | ( ~x510 & n1186 ) ;
  assign n1197 = n1191 | n1194 ;
  assign n1198 = ( ~x383 & x511 ) | ( ~x383 & n1196 ) | ( x511 & n1196 ) ;
  assign n1199 = x383 & x511 ;
  assign n1200 = ( x254 & ~n1176 ) | ( x254 & n1195 ) | ( ~n1176 & n1195 ) ;
  assign n1201 = n1189 & n1197 ;
  assign n1202 = ( n1189 & n1198 ) | ( n1189 & ~n1201 ) | ( n1198 & ~n1201 ) ;
  assign n1203 = x127 & ~x255 ;
  assign n1204 = ( ~n1179 & n1200 ) | ( ~n1179 & n1203 ) | ( n1200 & n1203 ) ;
  assign n1205 = ( x383 & n1189 ) | ( x383 & n1199 ) | ( n1189 & n1199 ) ;
  assign n1206 = x127 & x255 ;
  assign n1207 = n1179 | n1204 ;
  assign n1208 = ( x127 & n865 ) | ( x127 & n1206 ) | ( n865 & n1206 ) ;
  assign n1209 = ( n1206 & ~n1207 ) | ( n1206 & n1208 ) | ( ~n1207 & n1208 ) ;
  assign n1210 = ( ~n1197 & n1199 ) | ( ~n1197 & n1205 ) | ( n1199 & n1205 ) ;
  assign n1211 = n1202 ^ x380 ^ 1'b0 ;
  assign n1212 = x124 & ~x252 ;
  assign n1213 = ( x125 & ~x253 ) | ( x125 & n1212 ) | ( ~x253 & n1212 ) ;
  assign n1214 = n1202 ^ x311 ^ 1'b0 ;
  assign n1215 = ( x311 & x439 ) | ( x311 & ~n1214 ) | ( x439 & ~n1214 ) ;
  assign n1216 = ( x380 & x508 ) | ( x380 & ~n1211 ) | ( x508 & ~n1211 ) ;
  assign n1217 = ( x126 & ~x254 ) | ( x126 & n1213 ) | ( ~x254 & n1213 ) ;
  assign n1218 = ( ~x127 & x255 ) | ( ~x127 & n1217 ) | ( x255 & n1217 ) ;
  assign n1219 = n865 & n1207 ;
  assign n1220 = ( n865 & n1218 ) | ( n865 & ~n1219 ) | ( n1218 & ~n1219 ) ;
  assign n1221 = n1220 ^ x55 ^ 1'b0 ;
  assign n1222 = ( x55 & x183 ) | ( x55 & ~n1221 ) | ( x183 & ~n1221 ) ;
  assign n1223 = n1220 ^ x52 ^ 1'b0 ;
  assign n1224 = ( x52 & x180 ) | ( x52 & ~n1223 ) | ( x180 & ~n1223 ) ;
  assign n1225 = n1202 ^ x309 ^ 1'b0 ;
  assign n1226 = n1202 ^ x308 ^ 1'b0 ;
  assign n1227 = ( x308 & x436 ) | ( x308 & ~n1226 ) | ( x436 & ~n1226 ) ;
  assign n1228 = n1220 ^ x53 ^ 1'b0 ;
  assign n1229 = n1202 ^ x310 ^ 1'b0 ;
  assign n1230 = n1220 ^ x50 ^ 1'b0 ;
  assign n1231 = n1220 ^ x54 ^ 1'b0 ;
  assign n1232 = ( x54 & x182 ) | ( x54 & ~n1231 ) | ( x182 & ~n1231 ) ;
  assign n1233 = n1202 ^ x306 ^ 1'b0 ;
  assign n1234 = ( x310 & x438 ) | ( x310 & ~n1229 ) | ( x438 & ~n1229 ) ;
  assign n1235 = ( x309 & x437 ) | ( x309 & ~n1225 ) | ( x437 & ~n1225 ) ;
  assign n1236 = ( x53 & x181 ) | ( x53 & ~n1228 ) | ( x181 & ~n1228 ) ;
  assign n1237 = n1220 ^ x49 ^ 1'b0 ;
  assign n1238 = ( x49 & x177 ) | ( x49 & ~n1237 ) | ( x177 & ~n1237 ) ;
  assign n1239 = n1235 & ~n1236 ;
  assign n1240 = ( x50 & x178 ) | ( x50 & ~n1230 ) | ( x178 & ~n1230 ) ;
  assign n1241 = n1202 ^ x307 ^ 1'b0 ;
  assign n1242 = ( x307 & x435 ) | ( x307 & ~n1241 ) | ( x435 & ~n1241 ) ;
  assign n1243 = n1220 ^ x51 ^ 1'b0 ;
  assign n1244 = n1232 & n1234 ;
  assign n1245 = n1215 & ~n1222 ;
  assign n1246 = ( x51 & x179 ) | ( x51 & ~n1243 ) | ( x179 & ~n1243 ) ;
  assign n1247 = ( n1234 & ~n1244 ) | ( n1234 & n1245 ) | ( ~n1244 & n1245 ) ;
  assign n1248 = n1220 ^ x48 ^ 1'b0 ;
  assign n1249 = ( x48 & x176 ) | ( x48 & ~n1248 ) | ( x176 & ~n1248 ) ;
  assign n1250 = n1202 ^ x305 ^ 1'b0 ;
  assign n1251 = ( x305 & x433 ) | ( x305 & ~n1250 ) | ( x433 & ~n1250 ) ;
  assign n1252 = ~n1238 & n1251 ;
  assign n1253 = n1242 | n1252 ;
  assign n1254 = ( x306 & x434 ) | ( x306 & ~n1233 ) | ( x434 & ~n1233 ) ;
  assign n1255 = ( ~n1240 & n1252 ) | ( ~n1240 & n1254 ) | ( n1252 & n1254 ) ;
  assign n1256 = ( ~n1246 & n1252 ) | ( ~n1246 & n1253 ) | ( n1252 & n1253 ) ;
  assign n1257 = ~n1224 & n1227 ;
  assign n1258 = ( ~n1239 & n1247 ) | ( ~n1239 & n1257 ) | ( n1247 & n1257 ) ;
  assign n1259 = n1239 | n1258 ;
  assign n1260 = n1202 ^ x304 ^ 1'b0 ;
  assign n1261 = ( x304 & x432 ) | ( x304 & ~n1260 ) | ( x432 & ~n1260 ) ;
  assign n1262 = ~n1215 & n1222 ;
  assign n1263 = n1255 | n1256 ;
  assign n1264 = n1249 & ~n1261 ;
  assign n1265 = ( n1238 & ~n1251 ) | ( n1238 & n1264 ) | ( ~n1251 & n1264 ) ;
  assign n1266 = ( n1240 & ~n1254 ) | ( n1240 & n1265 ) | ( ~n1254 & n1265 ) ;
  assign n1267 = ( ~n1242 & n1246 ) | ( ~n1242 & n1266 ) | ( n1246 & n1266 ) ;
  assign n1268 = ( ~n1259 & n1262 ) | ( ~n1259 & n1267 ) | ( n1262 & n1267 ) ;
  assign n1269 = ~n1249 & n1261 ;
  assign n1270 = ( n1259 & n1263 ) | ( n1259 & ~n1269 ) | ( n1263 & ~n1269 ) ;
  assign n1271 = n1224 & ~n1227 ;
  assign n1272 = ( ~n1235 & n1236 ) | ( ~n1235 & n1271 ) | ( n1236 & n1271 ) ;
  assign n1273 = ( n1232 & ~n1234 ) | ( n1232 & n1272 ) | ( ~n1234 & n1272 ) ;
  assign n1274 = ( ~n1215 & n1222 ) | ( ~n1215 & n1273 ) | ( n1222 & n1273 ) ;
  assign n1275 = n1220 ^ x63 ^ 1'b0 ;
  assign n1276 = ( x63 & x191 ) | ( x63 & ~n1275 ) | ( x191 & ~n1275 ) ;
  assign n1277 = n1202 ^ x317 ^ 1'b0 ;
  assign n1278 = n1202 ^ x318 ^ 1'b0 ;
  assign n1279 = n1220 ^ x61 ^ 1'b0 ;
  assign n1280 = n1202 ^ x319 ^ 1'b0 ;
  assign n1281 = ( x61 & x189 ) | ( x61 & ~n1279 ) | ( x189 & ~n1279 ) ;
  assign n1282 = n1202 ^ x316 ^ 1'b0 ;
  assign n1283 = ( x316 & x444 ) | ( x316 & ~n1282 ) | ( x444 & ~n1282 ) ;
  assign n1284 = n1220 ^ x125 ^ 1'b0 ;
  assign n1285 = n1202 ^ x382 ^ 1'b0 ;
  assign n1286 = ( x382 & x510 ) | ( x382 & ~n1285 ) | ( x510 & ~n1285 ) ;
  assign n1287 = ( x319 & x447 ) | ( x319 & ~n1280 ) | ( x447 & ~n1280 ) ;
  assign n1288 = n1220 ^ x62 ^ 1'b0 ;
  assign n1289 = ( x318 & x446 ) | ( x318 & ~n1278 ) | ( x446 & ~n1278 ) ;
  assign n1290 = ~n1276 & n1287 ;
  assign n1291 = ( x62 & x190 ) | ( x62 & ~n1288 ) | ( x190 & ~n1288 ) ;
  assign n1292 = n1289 & ~n1291 ;
  assign n1293 = ( x317 & x445 ) | ( x317 & ~n1277 ) | ( x445 & ~n1277 ) ;
  assign n1294 = n1220 ^ x60 ^ 1'b0 ;
  assign n1295 = ( x60 & x188 ) | ( x60 & ~n1294 ) | ( x188 & ~n1294 ) ;
  assign n1296 = ~n1281 & n1293 ;
  assign n1297 = n1290 | n1292 ;
  assign n1298 = n1283 & ~n1295 ;
  assign n1299 = n1202 ^ x381 ^ 1'b0 ;
  assign n1300 = n1220 ^ x43 ^ 1'b0 ;
  assign n1301 = n1220 ^ x42 ^ 1'b0 ;
  assign n1302 = ( x42 & x170 ) | ( x42 & ~n1301 ) | ( x170 & ~n1301 ) ;
  assign n1303 = ( x43 & x171 ) | ( x43 & ~n1300 ) | ( x171 & ~n1300 ) ;
  assign n1304 = n1220 ^ x126 ^ 1'b0 ;
  assign n1305 = n1220 ^ x124 ^ 1'b0 ;
  assign n1306 = n1202 ^ x298 ^ 1'b0 ;
  assign n1307 = n1209 & ~n1210 ;
  assign n1308 = ( x124 & x252 ) | ( x124 & ~n1305 ) | ( x252 & ~n1305 ) ;
  assign n1309 = n1202 ^ x299 ^ 1'b0 ;
  assign n1310 = ( x299 & x427 ) | ( x299 & ~n1309 ) | ( x427 & ~n1309 ) ;
  assign n1311 = ~n1303 & n1310 ;
  assign n1312 = ( x126 & x254 ) | ( x126 & ~n1304 ) | ( x254 & ~n1304 ) ;
  assign n1313 = ( n1296 & n1297 ) | ( n1296 & ~n1298 ) | ( n1297 & ~n1298 ) ;
  assign n1314 = n1298 | n1313 ;
  assign n1315 = ( x125 & x253 ) | ( x125 & ~n1284 ) | ( x253 & ~n1284 ) ;
  assign n1316 = n1286 & ~n1312 ;
  assign n1317 = ( x381 & x509 ) | ( x381 & ~n1299 ) | ( x509 & ~n1299 ) ;
  assign n1318 = n1315 & n1317 ;
  assign n1319 = ( n1316 & n1317 ) | ( n1316 & ~n1318 ) | ( n1317 & ~n1318 ) ;
  assign n1320 = n1216 & ~n1308 ;
  assign n1321 = ( n1307 & n1319 ) | ( n1307 & ~n1320 ) | ( n1319 & ~n1320 ) ;
  assign n1322 = ~n1216 & n1308 ;
  assign n1323 = n1320 | n1321 ;
  assign n1324 = ( x298 & x426 ) | ( x298 & ~n1306 ) | ( x426 & ~n1306 ) ;
  assign n1325 = n1311 | n1324 ;
  assign n1326 = ( ~n1302 & n1311 ) | ( ~n1302 & n1325 ) | ( n1311 & n1325 ) ;
  assign n1327 = ~n1283 & n1295 ;
  assign n1328 = ( n1315 & ~n1317 ) | ( n1315 & n1322 ) | ( ~n1317 & n1322 ) ;
  assign n1329 = ( ~n1286 & n1312 ) | ( ~n1286 & n1328 ) | ( n1312 & n1328 ) ;
  assign n1330 = ( n1281 & ~n1293 ) | ( n1281 & n1327 ) | ( ~n1293 & n1327 ) ;
  assign n1331 = ( ~n1289 & n1291 ) | ( ~n1289 & n1330 ) | ( n1291 & n1330 ) ;
  assign n1332 = n1290 & n1331 ;
  assign n1333 = ( ~n1209 & n1210 ) | ( ~n1209 & n1329 ) | ( n1210 & n1329 ) ;
  assign n1334 = n1202 ^ x288 ^ 1'b0 ;
  assign n1335 = ( x288 & x416 ) | ( x288 & ~n1334 ) | ( x416 & ~n1334 ) ;
  assign n1336 = n1220 ^ x36 ^ 1'b0 ;
  assign n1337 = ( x36 & x164 ) | ( x36 & ~n1336 ) | ( x164 & ~n1336 ) ;
  assign n1338 = n1202 ^ x292 ^ 1'b0 ;
  assign n1339 = ( x292 & x420 ) | ( x292 & ~n1338 ) | ( x420 & ~n1338 ) ;
  assign n1340 = ~n1337 & n1339 ;
  assign n1341 = n1220 ^ x37 ^ 1'b0 ;
  assign n1342 = ( x37 & x165 ) | ( x37 & ~n1341 ) | ( x165 & ~n1341 ) ;
  assign n1343 = n1202 ^ x293 ^ 1'b0 ;
  assign n1344 = ( x293 & x421 ) | ( x293 & ~n1343 ) | ( x421 & ~n1343 ) ;
  assign n1345 = ~n1342 & n1344 ;
  assign n1346 = n1220 ^ x39 ^ 1'b0 ;
  assign n1347 = ( x39 & x167 ) | ( x39 & ~n1346 ) | ( x167 & ~n1346 ) ;
  assign n1348 = n1202 ^ x295 ^ 1'b0 ;
  assign n1349 = ( x295 & x423 ) | ( x295 & ~n1348 ) | ( x423 & ~n1348 ) ;
  assign n1350 = ~n1347 & n1349 ;
  assign n1351 = n1220 ^ x38 ^ 1'b0 ;
  assign n1352 = ( x38 & x166 ) | ( x38 & ~n1351 ) | ( x166 & ~n1351 ) ;
  assign n1353 = n1202 ^ x294 ^ 1'b0 ;
  assign n1354 = ( x294 & x422 ) | ( x294 & ~n1353 ) | ( x422 & ~n1353 ) ;
  assign n1355 = n1350 | n1354 ;
  assign n1356 = ( n1350 & ~n1352 ) | ( n1350 & n1355 ) | ( ~n1352 & n1355 ) ;
  assign n1357 = ( n1340 & n1345 ) | ( n1340 & ~n1356 ) | ( n1345 & ~n1356 ) ;
  assign n1358 = n1220 ^ x33 ^ 1'b0 ;
  assign n1359 = ( x33 & x161 ) | ( x33 & ~n1358 ) | ( x161 & ~n1358 ) ;
  assign n1360 = n1202 ^ x289 ^ 1'b0 ;
  assign n1361 = ( x289 & x417 ) | ( x289 & ~n1360 ) | ( x417 & ~n1360 ) ;
  assign n1362 = n1220 ^ x35 ^ 1'b0 ;
  assign n1363 = ( x35 & x163 ) | ( x35 & ~n1362 ) | ( x163 & ~n1362 ) ;
  assign n1364 = n1202 ^ x291 ^ 1'b0 ;
  assign n1365 = ( x291 & x419 ) | ( x291 & ~n1364 ) | ( x419 & ~n1364 ) ;
  assign n1366 = n1202 ^ x290 ^ 1'b0 ;
  assign n1367 = ( x290 & x418 ) | ( x290 & ~n1366 ) | ( x418 & ~n1366 ) ;
  assign n1368 = n1220 ^ x34 ^ 1'b0 ;
  assign n1369 = ( x34 & x162 ) | ( x34 & ~n1368 ) | ( x162 & ~n1368 ) ;
  assign n1370 = n1220 ^ x32 ^ 1'b0 ;
  assign n1371 = ( x32 & x160 ) | ( x32 & ~n1370 ) | ( x160 & ~n1370 ) ;
  assign n1372 = ~n1335 & n1371 ;
  assign n1373 = ( n1359 & ~n1361 ) | ( n1359 & n1372 ) | ( ~n1361 & n1372 ) ;
  assign n1374 = ( ~n1367 & n1369 ) | ( ~n1367 & n1373 ) | ( n1369 & n1373 ) ;
  assign n1375 = ( n1363 & ~n1365 ) | ( n1363 & n1374 ) | ( ~n1365 & n1374 ) ;
  assign n1376 = n1337 & ~n1339 ;
  assign n1377 = ( n1342 & ~n1344 ) | ( n1342 & n1376 ) | ( ~n1344 & n1376 ) ;
  assign n1378 = ( n1352 & ~n1354 ) | ( n1352 & n1377 ) | ( ~n1354 & n1377 ) ;
  assign n1379 = ~n1350 & n1378 ;
  assign n1380 = n1356 | n1357 ;
  assign n1381 = n1375 & n1380 ;
  assign n1382 = ( n1375 & n1379 ) | ( n1375 & ~n1381 ) | ( n1379 & ~n1381 ) ;
  assign n1383 = n1220 ^ x5 ^ 1'b0 ;
  assign n1384 = n1202 ^ x262 ^ 1'b0 ;
  assign n1385 = n1220 ^ x1 ^ 1'b0 ;
  assign n1386 = n1202 ^ x264 ^ 1'b0 ;
  assign n1387 = n1202 ^ x257 ^ 1'b0 ;
  assign n1388 = n1202 ^ x259 ^ 1'b0 ;
  assign n1389 = n1202 ^ x260 ^ 1'b0 ;
  assign n1390 = n1220 ^ x6 ^ 1'b0 ;
  assign n1391 = n1202 ^ x263 ^ 1'b0 ;
  assign n1392 = n1220 ^ x3 ^ 1'b0 ;
  assign n1393 = n1202 ^ x256 ^ 1'b0 ;
  assign n1394 = n1220 ^ x2 ^ 1'b0 ;
  assign n1395 = ( x256 & x384 ) | ( x256 & ~n1393 ) | ( x384 & ~n1393 ) ;
  assign n1396 = n1202 ^ x266 ^ 1'b0 ;
  assign n1397 = n1202 ^ x265 ^ 1'b0 ;
  assign n1398 = n1220 ^ x4 ^ 1'b0 ;
  assign n1399 = n1220 ^ x7 ^ 1'b0 ;
  assign n1400 = n1220 ^ x0 ^ 1'b0 ;
  assign n1401 = ( x259 & x387 ) | ( x259 & ~n1388 ) | ( x387 & ~n1388 ) ;
  assign n1402 = ( x4 & x132 ) | ( x4 & ~n1398 ) | ( x132 & ~n1398 ) ;
  assign n1403 = n1220 ^ x9 ^ 1'b0 ;
  assign n1404 = ( x2 & x130 ) | ( x2 & ~n1394 ) | ( x130 & ~n1394 ) ;
  assign n1405 = ( x1 & x129 ) | ( x1 & ~n1385 ) | ( x129 & ~n1385 ) ;
  assign n1406 = ( x0 & x128 ) | ( x0 & ~n1400 ) | ( x128 & ~n1400 ) ;
  assign n1407 = ( x3 & x131 ) | ( x3 & ~n1392 ) | ( x131 & ~n1392 ) ;
  assign n1408 = ~n1395 & n1406 ;
  assign n1409 = ( x5 & x133 ) | ( x5 & ~n1383 ) | ( x133 & ~n1383 ) ;
  assign n1410 = n1220 ^ x8 ^ 1'b0 ;
  assign n1411 = n1202 ^ x258 ^ 1'b0 ;
  assign n1412 = ( x258 & x386 ) | ( x258 & ~n1411 ) | ( x386 & ~n1411 ) ;
  assign n1413 = ( x257 & x385 ) | ( x257 & ~n1387 ) | ( x385 & ~n1387 ) ;
  assign n1414 = ( n1405 & n1408 ) | ( n1405 & ~n1413 ) | ( n1408 & ~n1413 ) ;
  assign n1415 = ( n1404 & ~n1412 ) | ( n1404 & n1414 ) | ( ~n1412 & n1414 ) ;
  assign n1416 = n1202 ^ x261 ^ 1'b0 ;
  assign n1417 = ( x261 & x389 ) | ( x261 & ~n1416 ) | ( x389 & ~n1416 ) ;
  assign n1418 = ( x262 & x390 ) | ( x262 & ~n1384 ) | ( x390 & ~n1384 ) ;
  assign n1419 = ( x265 & x393 ) | ( x265 & ~n1397 ) | ( x393 & ~n1397 ) ;
  assign n1420 = ( ~n1401 & n1407 ) | ( ~n1401 & n1415 ) | ( n1407 & n1415 ) ;
  assign n1421 = ( x260 & x388 ) | ( x260 & ~n1389 ) | ( x388 & ~n1389 ) ;
  assign n1422 = ( n1402 & n1420 ) | ( n1402 & ~n1421 ) | ( n1420 & ~n1421 ) ;
  assign n1423 = ( x7 & x135 ) | ( x7 & ~n1399 ) | ( x135 & ~n1399 ) ;
  assign n1424 = ( x263 & x391 ) | ( x263 & ~n1391 ) | ( x391 & ~n1391 ) ;
  assign n1425 = ( x8 & x136 ) | ( x8 & ~n1410 ) | ( x136 & ~n1410 ) ;
  assign n1426 = ( x6 & x134 ) | ( x6 & ~n1390 ) | ( x134 & ~n1390 ) ;
  assign n1427 = ( x264 & x392 ) | ( x264 & ~n1386 ) | ( x392 & ~n1386 ) ;
  assign n1428 = ( n1409 & ~n1417 ) | ( n1409 & n1422 ) | ( ~n1417 & n1422 ) ;
  assign n1429 = ( x9 & x137 ) | ( x9 & ~n1403 ) | ( x137 & ~n1403 ) ;
  assign n1430 = ( ~n1418 & n1426 ) | ( ~n1418 & n1428 ) | ( n1426 & n1428 ) ;
  assign n1431 = ( n1423 & ~n1424 ) | ( n1423 & n1430 ) | ( ~n1424 & n1430 ) ;
  assign n1432 = ( n1425 & ~n1427 ) | ( n1425 & n1431 ) | ( ~n1427 & n1431 ) ;
  assign n1433 = ( x266 & x394 ) | ( x266 & ~n1396 ) | ( x394 & ~n1396 ) ;
  assign n1434 = n1220 ^ x16 ^ 1'b0 ;
  assign n1435 = n1220 ^ x10 ^ 1'b0 ;
  assign n1436 = n1220 ^ x18 ^ 1'b0 ;
  assign n1437 = ( x10 & x138 ) | ( x10 & ~n1435 ) | ( x138 & ~n1435 ) ;
  assign n1438 = n1202 ^ x272 ^ 1'b0 ;
  assign n1439 = n1220 ^ x15 ^ 1'b0 ;
  assign n1440 = n1202 ^ x275 ^ 1'b0 ;
  assign n1441 = n1202 ^ x271 ^ 1'b0 ;
  assign n1442 = ( x275 & x403 ) | ( x275 & ~n1440 ) | ( x403 & ~n1440 ) ;
  assign n1443 = n1202 ^ x273 ^ 1'b0 ;
  assign n1444 = n1202 ^ x276 ^ 1'b0 ;
  assign n1445 = n1202 ^ x269 ^ 1'b0 ;
  assign n1446 = ( x269 & x397 ) | ( x269 & ~n1445 ) | ( x397 & ~n1445 ) ;
  assign n1447 = ( x273 & x401 ) | ( x273 & ~n1443 ) | ( x401 & ~n1443 ) ;
  assign n1448 = n1202 ^ x270 ^ 1'b0 ;
  assign n1449 = n1220 ^ x14 ^ 1'b0 ;
  assign n1450 = ( x14 & x142 ) | ( x14 & ~n1449 ) | ( x142 & ~n1449 ) ;
  assign n1451 = ( x270 & x398 ) | ( x270 & ~n1448 ) | ( x398 & ~n1448 ) ;
  assign n1452 = ( x15 & x143 ) | ( x15 & ~n1439 ) | ( x143 & ~n1439 ) ;
  assign n1453 = n1220 ^ x17 ^ 1'b0 ;
  assign n1454 = ( x18 & x146 ) | ( x18 & ~n1436 ) | ( x146 & ~n1436 ) ;
  assign n1455 = n1202 ^ x268 ^ 1'b0 ;
  assign n1456 = n1202 ^ x267 ^ 1'b0 ;
  assign n1457 = ( x267 & x395 ) | ( x267 & ~n1456 ) | ( x395 & ~n1456 ) ;
  assign n1458 = n1220 ^ x19 ^ 1'b0 ;
  assign n1459 = n1220 ^ x11 ^ 1'b0 ;
  assign n1460 = ( x17 & x145 ) | ( x17 & ~n1453 ) | ( x145 & ~n1453 ) ;
  assign n1461 = ( x19 & x147 ) | ( x19 & ~n1458 ) | ( x147 & ~n1458 ) ;
  assign n1462 = n1220 ^ x20 ^ 1'b0 ;
  assign n1463 = ( x268 & x396 ) | ( x268 & ~n1455 ) | ( x396 & ~n1455 ) ;
  assign n1464 = ( x276 & x404 ) | ( x276 & ~n1444 ) | ( x404 & ~n1444 ) ;
  assign n1465 = ( ~n1419 & n1429 ) | ( ~n1419 & n1432 ) | ( n1429 & n1432 ) ;
  assign n1466 = ( x11 & x139 ) | ( x11 & ~n1459 ) | ( x139 & ~n1459 ) ;
  assign n1467 = ( ~n1433 & n1437 ) | ( ~n1433 & n1465 ) | ( n1437 & n1465 ) ;
  assign n1468 = ( x16 & x144 ) | ( x16 & ~n1434 ) | ( x144 & ~n1434 ) ;
  assign n1469 = n1220 ^ x13 ^ 1'b0 ;
  assign n1470 = n1220 ^ x12 ^ 1'b0 ;
  assign n1471 = ( x12 & x140 ) | ( x12 & ~n1470 ) | ( x140 & ~n1470 ) ;
  assign n1472 = ( x13 & x141 ) | ( x13 & ~n1469 ) | ( x141 & ~n1469 ) ;
  assign n1473 = ( ~n1457 & n1466 ) | ( ~n1457 & n1467 ) | ( n1466 & n1467 ) ;
  assign n1474 = ( ~n1463 & n1471 ) | ( ~n1463 & n1473 ) | ( n1471 & n1473 ) ;
  assign n1475 = ( x271 & x399 ) | ( x271 & ~n1441 ) | ( x399 & ~n1441 ) ;
  assign n1476 = ( x20 & x148 ) | ( x20 & ~n1462 ) | ( x148 & ~n1462 ) ;
  assign n1477 = n1202 ^ x274 ^ 1'b0 ;
  assign n1478 = ( x274 & x402 ) | ( x274 & ~n1477 ) | ( x402 & ~n1477 ) ;
  assign n1479 = ( ~n1446 & n1472 ) | ( ~n1446 & n1474 ) | ( n1472 & n1474 ) ;
  assign n1480 = ( n1450 & ~n1451 ) | ( n1450 & n1479 ) | ( ~n1451 & n1479 ) ;
  assign n1481 = ( n1452 & ~n1475 ) | ( n1452 & n1480 ) | ( ~n1475 & n1480 ) ;
  assign n1482 = ( x272 & x400 ) | ( x272 & ~n1438 ) | ( x400 & ~n1438 ) ;
  assign n1483 = ( n1468 & n1481 ) | ( n1468 & ~n1482 ) | ( n1481 & ~n1482 ) ;
  assign n1484 = ( ~n1447 & n1460 ) | ( ~n1447 & n1483 ) | ( n1460 & n1483 ) ;
  assign n1485 = ( n1454 & ~n1478 ) | ( n1454 & n1484 ) | ( ~n1478 & n1484 ) ;
  assign n1486 = ( ~n1442 & n1461 ) | ( ~n1442 & n1485 ) | ( n1461 & n1485 ) ;
  assign n1487 = n1220 ^ x22 ^ 1'b0 ;
  assign n1488 = ( ~n1464 & n1476 ) | ( ~n1464 & n1486 ) | ( n1476 & n1486 ) ;
  assign n1489 = n1202 ^ x282 ^ 1'b0 ;
  assign n1490 = n1202 ^ x278 ^ 1'b0 ;
  assign n1491 = n1202 ^ x281 ^ 1'b0 ;
  assign n1492 = n1220 ^ x21 ^ 1'b0 ;
  assign n1493 = ( x281 & x409 ) | ( x281 & ~n1491 ) | ( x409 & ~n1491 ) ;
  assign n1494 = n1202 ^ x279 ^ 1'b0 ;
  assign n1495 = n1202 ^ x280 ^ 1'b0 ;
  assign n1496 = ( x279 & x407 ) | ( x279 & ~n1494 ) | ( x407 & ~n1494 ) ;
  assign n1497 = n1202 ^ x277 ^ 1'b0 ;
  assign n1498 = n1220 ^ x30 ^ 1'b0 ;
  assign n1499 = n1202 ^ x283 ^ 1'b0 ;
  assign n1500 = n1220 ^ x24 ^ 1'b0 ;
  assign n1501 = ( x21 & x149 ) | ( x21 & ~n1492 ) | ( x149 & ~n1492 ) ;
  assign n1502 = ( x283 & x411 ) | ( x283 & ~n1499 ) | ( x411 & ~n1499 ) ;
  assign n1503 = ( x24 & x152 ) | ( x24 & ~n1500 ) | ( x152 & ~n1500 ) ;
  assign n1504 = ( x278 & x406 ) | ( x278 & ~n1490 ) | ( x406 & ~n1490 ) ;
  assign n1505 = n1202 ^ x284 ^ 1'b0 ;
  assign n1506 = ( x22 & x150 ) | ( x22 & ~n1487 ) | ( x150 & ~n1487 ) ;
  assign n1507 = ~n1363 & n1365 ;
  assign n1508 = n1202 ^ x287 ^ 1'b0 ;
  assign n1509 = ( x277 & x405 ) | ( x277 & ~n1497 ) | ( x405 & ~n1497 ) ;
  assign n1510 = ( n1488 & n1501 ) | ( n1488 & ~n1509 ) | ( n1501 & ~n1509 ) ;
  assign n1511 = ( x284 & x412 ) | ( x284 & ~n1505 ) | ( x412 & ~n1505 ) ;
  assign n1512 = ~n1359 & n1361 ;
  assign n1513 = n1202 ^ x285 ^ 1'b0 ;
  assign n1514 = n1220 ^ x28 ^ 1'b0 ;
  assign n1515 = ( x28 & x156 ) | ( x28 & ~n1514 ) | ( x156 & ~n1514 ) ;
  assign n1516 = ( ~n1504 & n1506 ) | ( ~n1504 & n1510 ) | ( n1506 & n1510 ) ;
  assign n1517 = ( x282 & x410 ) | ( x282 & ~n1489 ) | ( x410 & ~n1489 ) ;
  assign n1518 = n1220 ^ x23 ^ 1'b0 ;
  assign n1519 = ( x23 & x151 ) | ( x23 & ~n1518 ) | ( x151 & ~n1518 ) ;
  assign n1520 = ( ~n1496 & n1516 ) | ( ~n1496 & n1519 ) | ( n1516 & n1519 ) ;
  assign n1521 = ( x280 & x408 ) | ( x280 & ~n1495 ) | ( x408 & ~n1495 ) ;
  assign n1522 = ( n1503 & n1520 ) | ( n1503 & ~n1521 ) | ( n1520 & ~n1521 ) ;
  assign n1523 = n1367 & ~n1369 ;
  assign n1524 = ( n1507 & ~n1512 ) | ( n1507 & n1523 ) | ( ~n1512 & n1523 ) ;
  assign n1525 = n1220 ^ x25 ^ 1'b0 ;
  assign n1526 = ( x25 & x153 ) | ( x25 & ~n1525 ) | ( x153 & ~n1525 ) ;
  assign n1527 = ( ~n1493 & n1522 ) | ( ~n1493 & n1526 ) | ( n1522 & n1526 ) ;
  assign n1528 = n1220 ^ x26 ^ 1'b0 ;
  assign n1529 = ( x26 & x154 ) | ( x26 & ~n1528 ) | ( x154 & ~n1528 ) ;
  assign n1530 = n1220 ^ x27 ^ 1'b0 ;
  assign n1531 = ( x27 & x155 ) | ( x27 & ~n1530 ) | ( x155 & ~n1530 ) ;
  assign n1532 = n1202 ^ x286 ^ 1'b0 ;
  assign n1533 = ( x30 & x158 ) | ( x30 & ~n1498 ) | ( x158 & ~n1498 ) ;
  assign n1534 = ( x286 & x414 ) | ( x286 & ~n1532 ) | ( x414 & ~n1532 ) ;
  assign n1535 = ( x287 & x415 ) | ( x287 & ~n1508 ) | ( x415 & ~n1508 ) ;
  assign n1536 = n1220 ^ x29 ^ 1'b0 ;
  assign n1537 = ( x29 & x157 ) | ( x29 & ~n1536 ) | ( x157 & ~n1536 ) ;
  assign n1538 = ( x285 & x413 ) | ( x285 & ~n1513 ) | ( x413 & ~n1513 ) ;
  assign n1539 = ( ~n1517 & n1527 ) | ( ~n1517 & n1529 ) | ( n1527 & n1529 ) ;
  assign n1540 = ( ~n1502 & n1531 ) | ( ~n1502 & n1539 ) | ( n1531 & n1539 ) ;
  assign n1541 = ( ~n1511 & n1515 ) | ( ~n1511 & n1540 ) | ( n1515 & n1540 ) ;
  assign n1542 = ( n1537 & ~n1538 ) | ( n1537 & n1541 ) | ( ~n1538 & n1541 ) ;
  assign n1543 = n1220 ^ x31 ^ 1'b0 ;
  assign n1544 = ( x31 & x159 ) | ( x31 & ~n1543 ) | ( x159 & ~n1543 ) ;
  assign n1545 = ( n1533 & ~n1534 ) | ( n1533 & n1542 ) | ( ~n1534 & n1542 ) ;
  assign n1546 = ( ~n1535 & n1544 ) | ( ~n1535 & n1545 ) | ( n1544 & n1545 ) ;
  assign n1547 = ~n1524 & n1546 ;
  assign n1548 = ~n1512 & n1547 ;
  assign n1549 = ( ~n1356 & n1357 ) | ( ~n1356 & n1548 ) | ( n1357 & n1548 ) ;
  assign n1550 = ~n1357 & n1549 ;
  assign n1551 = n1347 & ~n1349 ;
  assign n1552 = n1335 & n1371 ;
  assign n1553 = ( ~n1335 & n1550 ) | ( ~n1335 & n1552 ) | ( n1550 & n1552 ) ;
  assign n1554 = ( n1382 & n1551 ) | ( n1382 & ~n1553 ) | ( n1551 & ~n1553 ) ;
  assign n1555 = n1553 | n1554 ;
  assign n1556 = n1220 ^ x47 ^ 1'b0 ;
  assign n1557 = n1202 ^ x302 ^ 1'b0 ;
  assign n1558 = n1220 ^ x46 ^ 1'b0 ;
  assign n1559 = ( x302 & x430 ) | ( x302 & ~n1557 ) | ( x430 & ~n1557 ) ;
  assign n1560 = ( x46 & x174 ) | ( x46 & ~n1558 ) | ( x174 & ~n1558 ) ;
  assign n1561 = n1559 & ~n1560 ;
  assign n1562 = n1202 ^ x296 ^ 1'b0 ;
  assign n1563 = ( x296 & x424 ) | ( x296 & ~n1562 ) | ( x424 & ~n1562 ) ;
  assign n1564 = ( x47 & x175 ) | ( x47 & ~n1556 ) | ( x175 & ~n1556 ) ;
  assign n1565 = n1202 ^ x297 ^ 1'b0 ;
  assign n1566 = n1202 ^ x303 ^ 1'b0 ;
  assign n1567 = n1220 ^ x40 ^ 1'b0 ;
  assign n1568 = ( x303 & x431 ) | ( x303 & ~n1566 ) | ( x431 & ~n1566 ) ;
  assign n1569 = ( x297 & x425 ) | ( x297 & ~n1565 ) | ( x425 & ~n1565 ) ;
  assign n1570 = ( x40 & x168 ) | ( x40 & ~n1567 ) | ( x168 & ~n1567 ) ;
  assign n1571 = ~n1564 & n1568 ;
  assign n1572 = n1202 ^ x301 ^ 1'b0 ;
  assign n1573 = ( x301 & x429 ) | ( x301 & ~n1572 ) | ( x429 & ~n1572 ) ;
  assign n1574 = n1220 ^ x44 ^ 1'b0 ;
  assign n1575 = n1561 | n1571 ;
  assign n1576 = n1202 ^ x300 ^ 1'b0 ;
  assign n1577 = n1563 & ~n1570 ;
  assign n1578 = n1220 ^ x41 ^ 1'b0 ;
  assign n1579 = ( x41 & x169 ) | ( x41 & ~n1578 ) | ( x169 & ~n1578 ) ;
  assign n1580 = n1569 & ~n1579 ;
  assign n1581 = ( ~n1326 & n1577 ) | ( ~n1326 & n1580 ) | ( n1577 & n1580 ) ;
  assign n1582 = ( x300 & x428 ) | ( x300 & ~n1576 ) | ( x428 & ~n1576 ) ;
  assign n1583 = ( x44 & x172 ) | ( x44 & ~n1574 ) | ( x172 & ~n1574 ) ;
  assign n1584 = n1220 ^ x45 ^ 1'b0 ;
  assign n1585 = ( x45 & x173 ) | ( x45 & ~n1584 ) | ( x173 & ~n1584 ) ;
  assign n1586 = ( n1326 & ~n1575 ) | ( n1326 & n1581 ) | ( ~n1575 & n1581 ) ;
  assign n1587 = n1582 & ~n1583 ;
  assign n1588 = n1555 & ~n1586 ;
  assign n1589 = n1573 & ~n1585 ;
  assign n1590 = ( ~n1575 & n1587 ) | ( ~n1575 & n1589 ) | ( n1587 & n1589 ) ;
  assign n1591 = ~n1563 & n1570 ;
  assign n1592 = ( ~n1569 & n1579 ) | ( ~n1569 & n1591 ) | ( n1579 & n1591 ) ;
  assign n1593 = ( n1302 & ~n1324 ) | ( n1302 & n1592 ) | ( ~n1324 & n1592 ) ;
  assign n1594 = ( n1303 & ~n1310 ) | ( n1303 & n1593 ) | ( ~n1310 & n1593 ) ;
  assign n1595 = ( ~n1575 & n1590 ) | ( ~n1575 & n1594 ) | ( n1590 & n1594 ) ;
  assign n1596 = ~n1590 & n1595 ;
  assign n1597 = ~n1575 & n1588 ;
  assign n1598 = ~n1582 & n1583 ;
  assign n1599 = ( ~n1573 & n1585 ) | ( ~n1573 & n1598 ) | ( n1585 & n1598 ) ;
  assign n1600 = ( ~n1559 & n1560 ) | ( ~n1559 & n1599 ) | ( n1560 & n1599 ) ;
  assign n1601 = ~n1590 & n1597 ;
  assign n1602 = n1571 & n1600 ;
  assign n1603 = ( n1600 & n1601 ) | ( n1600 & ~n1602 ) | ( n1601 & ~n1602 ) ;
  assign n1604 = n1564 & ~n1568 ;
  assign n1605 = ( n1596 & ~n1603 ) | ( n1596 & n1604 ) | ( ~n1603 & n1604 ) ;
  assign n1606 = n1603 | n1605 ;
  assign n1607 = ( ~n1269 & n1270 ) | ( ~n1269 & n1606 ) | ( n1270 & n1606 ) ;
  assign n1608 = ~n1270 & n1607 ;
  assign n1609 = ( n1268 & n1274 ) | ( n1268 & ~n1608 ) | ( n1274 & ~n1608 ) ;
  assign n1610 = n1608 | n1609 ;
  assign n1611 = n1202 ^ x312 ^ 1'b0 ;
  assign n1612 = n1220 ^ x58 ^ 1'b0 ;
  assign n1613 = n1220 ^ x57 ^ 1'b0 ;
  assign n1614 = ( x57 & x185 ) | ( x57 & ~n1613 ) | ( x185 & ~n1613 ) ;
  assign n1615 = n1220 ^ x56 ^ 1'b0 ;
  assign n1616 = ( x56 & x184 ) | ( x56 & ~n1615 ) | ( x184 & ~n1615 ) ;
  assign n1617 = n1202 ^ x313 ^ 1'b0 ;
  assign n1618 = ( x313 & x441 ) | ( x313 & ~n1617 ) | ( x441 & ~n1617 ) ;
  assign n1619 = ( x312 & x440 ) | ( x312 & ~n1611 ) | ( x440 & ~n1611 ) ;
  assign n1620 = ( n1314 & ~n1614 ) | ( n1314 & n1618 ) | ( ~n1614 & n1618 ) ;
  assign n1621 = n1314 | n1619 ;
  assign n1622 = ( n1314 & ~n1616 ) | ( n1314 & n1621 ) | ( ~n1616 & n1621 ) ;
  assign n1623 = n1202 ^ x315 ^ 1'b0 ;
  assign n1624 = n1202 ^ x314 ^ 1'b0 ;
  assign n1625 = ( x314 & x442 ) | ( x314 & ~n1624 ) | ( x442 & ~n1624 ) ;
  assign n1626 = n1616 & ~n1619 ;
  assign n1627 = n1220 ^ x59 ^ 1'b0 ;
  assign n1628 = ( x59 & x187 ) | ( x59 & ~n1627 ) | ( x187 & ~n1627 ) ;
  assign n1629 = ( x315 & x443 ) | ( x315 & ~n1623 ) | ( x443 & ~n1623 ) ;
  assign n1630 = n1620 | n1622 ;
  assign n1631 = ( n1614 & ~n1618 ) | ( n1614 & n1626 ) | ( ~n1618 & n1626 ) ;
  assign n1632 = ~n1628 & n1629 ;
  assign n1633 = ( x58 & x186 ) | ( x58 & ~n1612 ) | ( x186 & ~n1612 ) ;
  assign n1634 = ( ~n1625 & n1631 ) | ( ~n1625 & n1633 ) | ( n1631 & n1633 ) ;
  assign n1635 = ( n1628 & ~n1629 ) | ( n1628 & n1634 ) | ( ~n1629 & n1634 ) ;
  assign n1636 = ~n1314 & n1635 ;
  assign n1637 = n1625 & ~n1633 ;
  assign n1638 = ( n1630 & ~n1632 ) | ( n1630 & n1637 ) | ( ~n1632 & n1637 ) ;
  assign n1639 = ( n1610 & ~n1632 ) | ( n1610 & n1638 ) | ( ~n1632 & n1638 ) ;
  assign n1640 = ~n1638 & n1639 ;
  assign n1641 = ( n1331 & ~n1332 ) | ( n1331 & n1640 ) | ( ~n1332 & n1640 ) ;
  assign n1642 = n1202 ^ x320 ^ 1'b0 ;
  assign n1643 = n1276 & ~n1287 ;
  assign n1644 = n1202 ^ x321 ^ 1'b0 ;
  assign n1645 = ( x321 & x449 ) | ( x321 & ~n1644 ) | ( x449 & ~n1644 ) ;
  assign n1646 = n1220 ^ x65 ^ 1'b0 ;
  assign n1647 = ( n1636 & ~n1641 ) | ( n1636 & n1643 ) | ( ~n1641 & n1643 ) ;
  assign n1648 = n1220 ^ x64 ^ 1'b0 ;
  assign n1649 = n1641 | n1647 ;
  assign n1650 = ( x320 & x448 ) | ( x320 & ~n1642 ) | ( x448 & ~n1642 ) ;
  assign n1651 = ( x65 & x193 ) | ( x65 & ~n1646 ) | ( x193 & ~n1646 ) ;
  assign n1652 = ( ~n1645 & n1649 ) | ( ~n1645 & n1651 ) | ( n1649 & n1651 ) ;
  assign n1653 = ( x64 & x192 ) | ( x64 & ~n1648 ) | ( x192 & ~n1648 ) ;
  assign n1654 = n1649 & n1652 ;
  assign n1655 = ~n1650 & n1653 ;
  assign n1656 = n1650 & n1653 ;
  assign n1657 = ( ~n1650 & n1654 ) | ( ~n1650 & n1656 ) | ( n1654 & n1656 ) ;
  assign n1658 = ( ~n1645 & n1651 ) | ( ~n1645 & n1655 ) | ( n1651 & n1655 ) ;
  assign n1659 = n1657 | n1658 ;
  assign n1660 = n1220 ^ x75 ^ 1'b0 ;
  assign n1661 = n1202 ^ x323 ^ 1'b0 ;
  assign n1662 = n1202 ^ x326 ^ 1'b0 ;
  assign n1663 = ( x326 & x454 ) | ( x326 & ~n1662 ) | ( x454 & ~n1662 ) ;
  assign n1664 = n1220 ^ x68 ^ 1'b0 ;
  assign n1665 = ( x68 & x196 ) | ( x68 & ~n1664 ) | ( x196 & ~n1664 ) ;
  assign n1666 = n1202 ^ x324 ^ 1'b0 ;
  assign n1667 = ( x324 & x452 ) | ( x324 & ~n1666 ) | ( x452 & ~n1666 ) ;
  assign n1668 = n1202 ^ x329 ^ 1'b0 ;
  assign n1669 = n1665 & ~n1667 ;
  assign n1670 = ( x329 & x457 ) | ( x329 & ~n1668 ) | ( x457 & ~n1668 ) ;
  assign n1671 = n1220 ^ x74 ^ 1'b0 ;
  assign n1672 = ( x75 & x203 ) | ( x75 & ~n1660 ) | ( x203 & ~n1660 ) ;
  assign n1673 = n1202 ^ x327 ^ 1'b0 ;
  assign n1674 = n1220 ^ x71 ^ 1'b0 ;
  assign n1675 = ( x327 & x455 ) | ( x327 & ~n1673 ) | ( x455 & ~n1673 ) ;
  assign n1676 = ( x71 & x199 ) | ( x71 & ~n1674 ) | ( x199 & ~n1674 ) ;
  assign n1677 = n1675 & ~n1676 ;
  assign n1678 = n1663 | n1677 ;
  assign n1679 = n1220 ^ x69 ^ 1'b0 ;
  assign n1680 = n1202 ^ x325 ^ 1'b0 ;
  assign n1681 = ( x325 & x453 ) | ( x325 & ~n1680 ) | ( x453 & ~n1680 ) ;
  assign n1682 = ( x69 & x197 ) | ( x69 & ~n1679 ) | ( x197 & ~n1679 ) ;
  assign n1683 = ( n1669 & ~n1681 ) | ( n1669 & n1682 ) | ( ~n1681 & n1682 ) ;
  assign n1684 = n1220 ^ x70 ^ 1'b0 ;
  assign n1685 = ( x70 & x198 ) | ( x70 & ~n1684 ) | ( x198 & ~n1684 ) ;
  assign n1686 = n1202 ^ x322 ^ 1'b0 ;
  assign n1687 = ( x322 & x450 ) | ( x322 & ~n1686 ) | ( x450 & ~n1686 ) ;
  assign n1688 = ( n1677 & n1678 ) | ( n1677 & ~n1685 ) | ( n1678 & ~n1685 ) ;
  assign n1689 = n1202 ^ x331 ^ 1'b0 ;
  assign n1690 = ( x74 & x202 ) | ( x74 & ~n1671 ) | ( x202 & ~n1671 ) ;
  assign n1691 = n1220 ^ x66 ^ 1'b0 ;
  assign n1692 = ( ~n1663 & n1683 ) | ( ~n1663 & n1685 ) | ( n1683 & n1685 ) ;
  assign n1693 = ( x66 & x194 ) | ( x66 & ~n1691 ) | ( x194 & ~n1691 ) ;
  assign n1694 = n1220 ^ x73 ^ 1'b0 ;
  assign n1695 = ( x331 & x459 ) | ( x331 & ~n1689 ) | ( x459 & ~n1689 ) ;
  assign n1696 = n1202 ^ x330 ^ 1'b0 ;
  assign n1697 = ( x73 & x201 ) | ( x73 & ~n1694 ) | ( x201 & ~n1694 ) ;
  assign n1698 = ~n1672 & n1695 ;
  assign n1699 = ( x330 & x458 ) | ( x330 & ~n1696 ) | ( x458 & ~n1696 ) ;
  assign n1700 = ( x323 & x451 ) | ( x323 & ~n1661 ) | ( x451 & ~n1661 ) ;
  assign n1701 = n1690 & n1699 ;
  assign n1702 = ( n1659 & ~n1687 ) | ( n1659 & n1693 ) | ( ~n1687 & n1693 ) ;
  assign n1703 = ~n1665 & n1667 ;
  assign n1704 = ( n1698 & n1699 ) | ( n1698 & ~n1701 ) | ( n1699 & ~n1701 ) ;
  assign n1705 = n1220 ^ x67 ^ 1'b0 ;
  assign n1706 = ( x67 & x195 ) | ( x67 & ~n1705 ) | ( x195 & ~n1705 ) ;
  assign n1707 = ( ~n1700 & n1702 ) | ( ~n1700 & n1706 ) | ( n1702 & n1706 ) ;
  assign n1708 = ( ~n1675 & n1676 ) | ( ~n1675 & n1692 ) | ( n1676 & n1692 ) ;
  assign n1709 = n1681 & ~n1682 ;
  assign n1710 = ( ~n1688 & n1703 ) | ( ~n1688 & n1709 ) | ( n1703 & n1709 ) ;
  assign n1711 = n1707 & ~n1710 ;
  assign n1712 = n1220 ^ x72 ^ 1'b0 ;
  assign n1713 = ( x72 & x200 ) | ( x72 & ~n1712 ) | ( x200 & ~n1712 ) ;
  assign n1714 = n1688 & n1711 ;
  assign n1715 = ( n1708 & n1711 ) | ( n1708 & ~n1714 ) | ( n1711 & ~n1714 ) ;
  assign n1716 = n1202 ^ x328 ^ 1'b0 ;
  assign n1717 = ( x328 & x456 ) | ( x328 & ~n1716 ) | ( x456 & ~n1716 ) ;
  assign n1718 = ~n1713 & n1717 ;
  assign n1719 = n1670 & ~n1697 ;
  assign n1720 = ( ~n1704 & n1718 ) | ( ~n1704 & n1719 ) | ( n1718 & n1719 ) ;
  assign n1721 = n1713 & ~n1717 ;
  assign n1722 = ( ~n1670 & n1697 ) | ( ~n1670 & n1721 ) | ( n1697 & n1721 ) ;
  assign n1723 = ( n1690 & ~n1699 ) | ( n1690 & n1722 ) | ( ~n1699 & n1722 ) ;
  assign n1724 = ( n1672 & ~n1695 ) | ( n1672 & n1723 ) | ( ~n1695 & n1723 ) ;
  assign n1725 = ( ~n1704 & n1715 ) | ( ~n1704 & n1720 ) | ( n1715 & n1720 ) ;
  assign n1726 = n1720 & n1725 ;
  assign n1727 = ( n1724 & n1725 ) | ( n1724 & ~n1726 ) | ( n1725 & ~n1726 ) ;
  assign n1728 = n1202 ^ x332 ^ 1'b0 ;
  assign n1729 = n1202 ^ x333 ^ 1'b0 ;
  assign n1730 = n1220 ^ x78 ^ 1'b0 ;
  assign n1731 = n1202 ^ x336 ^ 1'b0 ;
  assign n1732 = n1202 ^ x339 ^ 1'b0 ;
  assign n1733 = n1220 ^ x79 ^ 1'b0 ;
  assign n1734 = ( x79 & x207 ) | ( x79 & ~n1733 ) | ( x207 & ~n1733 ) ;
  assign n1735 = n1220 ^ x77 ^ 1'b0 ;
  assign n1736 = ( x336 & x464 ) | ( x336 & ~n1731 ) | ( x464 & ~n1731 ) ;
  assign n1737 = n1220 ^ x76 ^ 1'b0 ;
  assign n1738 = n1220 ^ x82 ^ 1'b0 ;
  assign n1739 = n1202 ^ x335 ^ 1'b0 ;
  assign n1740 = ( x76 & x204 ) | ( x76 & ~n1737 ) | ( x204 & ~n1737 ) ;
  assign n1741 = n1202 ^ x338 ^ 1'b0 ;
  assign n1742 = ( x78 & x206 ) | ( x78 & ~n1730 ) | ( x206 & ~n1730 ) ;
  assign n1743 = n1202 ^ x334 ^ 1'b0 ;
  assign n1744 = ( x334 & x462 ) | ( x334 & ~n1743 ) | ( x462 & ~n1743 ) ;
  assign n1745 = ( x335 & x463 ) | ( x335 & ~n1739 ) | ( x463 & ~n1739 ) ;
  assign n1746 = ~n1734 & n1745 ;
  assign n1747 = n1744 | n1746 ;
  assign n1748 = ( ~n1742 & n1746 ) | ( ~n1742 & n1747 ) | ( n1746 & n1747 ) ;
  assign n1749 = ( x77 & x205 ) | ( x77 & ~n1735 ) | ( x205 & ~n1735 ) ;
  assign n1750 = ( x332 & x460 ) | ( x332 & ~n1728 ) | ( x460 & ~n1728 ) ;
  assign n1751 = ( x82 & x210 ) | ( x82 & ~n1738 ) | ( x210 & ~n1738 ) ;
  assign n1752 = n1220 ^ x80 ^ 1'b0 ;
  assign n1753 = ( x80 & x208 ) | ( x80 & ~n1752 ) | ( x208 & ~n1752 ) ;
  assign n1754 = ~n1740 & n1750 ;
  assign n1755 = n1740 & ~n1750 ;
  assign n1756 = ( x333 & x461 ) | ( x333 & ~n1729 ) | ( x461 & ~n1729 ) ;
  assign n1757 = ~n1749 & n1756 ;
  assign n1758 = ( ~n1748 & n1754 ) | ( ~n1748 & n1757 ) | ( n1754 & n1757 ) ;
  assign n1759 = n1727 & ~n1758 ;
  assign n1760 = n1748 & n1759 ;
  assign n1761 = ( n1749 & n1755 ) | ( n1749 & ~n1756 ) | ( n1755 & ~n1756 ) ;
  assign n1762 = ( n1742 & ~n1744 ) | ( n1742 & n1761 ) | ( ~n1744 & n1761 ) ;
  assign n1763 = ( n1734 & ~n1745 ) | ( n1734 & n1762 ) | ( ~n1745 & n1762 ) ;
  assign n1764 = n1202 ^ x337 ^ 1'b0 ;
  assign n1765 = ( x337 & x465 ) | ( x337 & ~n1764 ) | ( x465 & ~n1764 ) ;
  assign n1766 = ( x339 & x467 ) | ( x339 & ~n1732 ) | ( x467 & ~n1732 ) ;
  assign n1767 = n1220 ^ x83 ^ 1'b0 ;
  assign n1768 = ( x83 & x211 ) | ( x83 & ~n1767 ) | ( x211 & ~n1767 ) ;
  assign n1769 = ( x338 & x466 ) | ( x338 & ~n1741 ) | ( x466 & ~n1741 ) ;
  assign n1770 = ( n1759 & ~n1760 ) | ( n1759 & n1763 ) | ( ~n1760 & n1763 ) ;
  assign n1771 = n1751 & n1769 ;
  assign n1772 = n1766 & ~n1768 ;
  assign n1773 = ( n1769 & ~n1771 ) | ( n1769 & n1772 ) | ( ~n1771 & n1772 ) ;
  assign n1774 = n1220 ^ x81 ^ 1'b0 ;
  assign n1775 = ( x81 & x209 ) | ( x81 & ~n1774 ) | ( x209 & ~n1774 ) ;
  assign n1776 = n1770 & ~n1773 ;
  assign n1777 = n1765 & n1775 ;
  assign n1778 = ( ~n1765 & n1776 ) | ( ~n1765 & n1777 ) | ( n1776 & n1777 ) ;
  assign n1779 = n1736 & n1753 ;
  assign n1780 = ( ~n1736 & n1778 ) | ( ~n1736 & n1779 ) | ( n1778 & n1779 ) ;
  assign n1781 = ~n1736 & n1753 ;
  assign n1782 = ( ~n1765 & n1775 ) | ( ~n1765 & n1781 ) | ( n1775 & n1781 ) ;
  assign n1783 = ( n1751 & ~n1769 ) | ( n1751 & n1782 ) | ( ~n1769 & n1782 ) ;
  assign n1784 = ( ~n1766 & n1768 ) | ( ~n1766 & n1783 ) | ( n1768 & n1783 ) ;
  assign n1785 = n1780 | n1784 ;
  assign n1786 = n1202 ^ x343 ^ 1'b0 ;
  assign n1787 = n1220 ^ x85 ^ 1'b0 ;
  assign n1788 = n1202 ^ x342 ^ 1'b0 ;
  assign n1789 = n1202 ^ x346 ^ 1'b0 ;
  assign n1790 = ( x343 & x471 ) | ( x343 & ~n1786 ) | ( x471 & ~n1786 ) ;
  assign n1791 = n1220 ^ x90 ^ 1'b0 ;
  assign n1792 = n1202 ^ x344 ^ 1'b0 ;
  assign n1793 = ( x342 & x470 ) | ( x342 & ~n1788 ) | ( x470 & ~n1788 ) ;
  assign n1794 = n1220 ^ x87 ^ 1'b0 ;
  assign n1795 = ( x87 & x215 ) | ( x87 & ~n1794 ) | ( x215 & ~n1794 ) ;
  assign n1796 = ( x346 & x474 ) | ( x346 & ~n1789 ) | ( x474 & ~n1789 ) ;
  assign n1797 = n1790 & ~n1795 ;
  assign n1798 = n1202 ^ x345 ^ 1'b0 ;
  assign n1799 = ( x90 & x218 ) | ( x90 & ~n1791 ) | ( x218 & ~n1791 ) ;
  assign n1800 = n1202 ^ x347 ^ 1'b0 ;
  assign n1801 = n1793 | n1797 ;
  assign n1802 = n1220 ^ x86 ^ 1'b0 ;
  assign n1803 = n1220 ^ x84 ^ 1'b0 ;
  assign n1804 = ( x85 & x213 ) | ( x85 & ~n1787 ) | ( x213 & ~n1787 ) ;
  assign n1805 = n1202 ^ x341 ^ 1'b0 ;
  assign n1806 = n1796 & n1799 ;
  assign n1807 = n1202 ^ x340 ^ 1'b0 ;
  assign n1808 = ( x84 & x212 ) | ( x84 & ~n1803 ) | ( x212 & ~n1803 ) ;
  assign n1809 = ( x340 & x468 ) | ( x340 & ~n1807 ) | ( x468 & ~n1807 ) ;
  assign n1810 = ~n1808 & n1809 ;
  assign n1811 = ( x341 & x469 ) | ( x341 & ~n1805 ) | ( x469 & ~n1805 ) ;
  assign n1812 = ~n1804 & n1811 ;
  assign n1813 = ( x86 & x214 ) | ( x86 & ~n1802 ) | ( x214 & ~n1802 ) ;
  assign n1814 = ( n1797 & n1801 ) | ( n1797 & ~n1813 ) | ( n1801 & ~n1813 ) ;
  assign n1815 = n1220 ^ x91 ^ 1'b0 ;
  assign n1816 = n1220 ^ x88 ^ 1'b0 ;
  assign n1817 = ( x344 & x472 ) | ( x344 & ~n1792 ) | ( x472 & ~n1792 ) ;
  assign n1818 = ( x91 & x219 ) | ( x91 & ~n1815 ) | ( x219 & ~n1815 ) ;
  assign n1819 = ( n1810 & n1812 ) | ( n1810 & ~n1814 ) | ( n1812 & ~n1814 ) ;
  assign n1820 = n1785 & ~n1819 ;
  assign n1821 = n1808 & ~n1809 ;
  assign n1822 = n1814 & n1820 ;
  assign n1823 = ( x347 & x475 ) | ( x347 & ~n1800 ) | ( x475 & ~n1800 ) ;
  assign n1824 = ( x88 & x216 ) | ( x88 & ~n1816 ) | ( x216 & ~n1816 ) ;
  assign n1825 = ~n1818 & n1823 ;
  assign n1826 = ( n1796 & ~n1806 ) | ( n1796 & n1825 ) | ( ~n1806 & n1825 ) ;
  assign n1827 = ( n1804 & ~n1811 ) | ( n1804 & n1821 ) | ( ~n1811 & n1821 ) ;
  assign n1828 = n1220 ^ x89 ^ 1'b0 ;
  assign n1829 = ( x89 & x217 ) | ( x89 & ~n1828 ) | ( x217 & ~n1828 ) ;
  assign n1830 = ( x345 & x473 ) | ( x345 & ~n1798 ) | ( x473 & ~n1798 ) ;
  assign n1831 = ( ~n1793 & n1813 ) | ( ~n1793 & n1827 ) | ( n1813 & n1827 ) ;
  assign n1832 = ( ~n1790 & n1795 ) | ( ~n1790 & n1831 ) | ( n1795 & n1831 ) ;
  assign n1833 = ( n1820 & ~n1822 ) | ( n1820 & n1832 ) | ( ~n1822 & n1832 ) ;
  assign n1834 = n1817 & ~n1824 ;
  assign n1835 = ~n1829 & n1830 ;
  assign n1836 = ( ~n1826 & n1834 ) | ( ~n1826 & n1835 ) | ( n1834 & n1835 ) ;
  assign n1837 = ~n1817 & n1824 ;
  assign n1838 = ( n1829 & ~n1830 ) | ( n1829 & n1837 ) | ( ~n1830 & n1837 ) ;
  assign n1839 = ( ~n1826 & n1833 ) | ( ~n1826 & n1836 ) | ( n1833 & n1836 ) ;
  assign n1840 = n1836 & n1839 ;
  assign n1841 = ( ~n1796 & n1799 ) | ( ~n1796 & n1838 ) | ( n1799 & n1838 ) ;
  assign n1842 = ( n1818 & ~n1823 ) | ( n1818 & n1841 ) | ( ~n1823 & n1841 ) ;
  assign n1843 = ( n1839 & ~n1840 ) | ( n1839 & n1842 ) | ( ~n1840 & n1842 ) ;
  assign n1844 = n1220 ^ x99 ^ 1'b0 ;
  assign n1845 = ( x99 & x227 ) | ( x99 & ~n1844 ) | ( x227 & ~n1844 ) ;
  assign n1846 = n1220 ^ x97 ^ 1'b0 ;
  assign n1847 = n1220 ^ x93 ^ 1'b0 ;
  assign n1848 = n1202 ^ x348 ^ 1'b0 ;
  assign n1849 = ( x93 & x221 ) | ( x93 & ~n1847 ) | ( x221 & ~n1847 ) ;
  assign n1850 = n1202 ^ x354 ^ 1'b0 ;
  assign n1851 = ( x348 & x476 ) | ( x348 & ~n1848 ) | ( x476 & ~n1848 ) ;
  assign n1852 = n1202 ^ x355 ^ 1'b0 ;
  assign n1853 = n1202 ^ x351 ^ 1'b0 ;
  assign n1854 = n1220 ^ x95 ^ 1'b0 ;
  assign n1855 = n1220 ^ x92 ^ 1'b0 ;
  assign n1856 = n1202 ^ x349 ^ 1'b0 ;
  assign n1857 = ( x92 & x220 ) | ( x92 & ~n1855 ) | ( x220 & ~n1855 ) ;
  assign n1858 = n1220 ^ x98 ^ 1'b0 ;
  assign n1859 = ( x98 & x226 ) | ( x98 & ~n1858 ) | ( x226 & ~n1858 ) ;
  assign n1860 = ( x355 & x483 ) | ( x355 & ~n1852 ) | ( x483 & ~n1852 ) ;
  assign n1861 = ( x354 & x482 ) | ( x354 & ~n1850 ) | ( x482 & ~n1850 ) ;
  assign n1862 = n1220 ^ x94 ^ 1'b0 ;
  assign n1863 = n1859 & n1861 ;
  assign n1864 = n1202 ^ x350 ^ 1'b0 ;
  assign n1865 = ( x349 & x477 ) | ( x349 & ~n1856 ) | ( x477 & ~n1856 ) ;
  assign n1866 = ( x350 & x478 ) | ( x350 & ~n1864 ) | ( x478 & ~n1864 ) ;
  assign n1867 = ( x94 & x222 ) | ( x94 & ~n1862 ) | ( x222 & ~n1862 ) ;
  assign n1868 = ( x351 & x479 ) | ( x351 & ~n1853 ) | ( x479 & ~n1853 ) ;
  assign n1869 = ( x95 & x223 ) | ( x95 & ~n1854 ) | ( x223 & ~n1854 ) ;
  assign n1870 = n1868 & ~n1869 ;
  assign n1871 = n1866 | n1870 ;
  assign n1872 = ( ~n1867 & n1870 ) | ( ~n1867 & n1871 ) | ( n1870 & n1871 ) ;
  assign n1873 = ~n1849 & n1865 ;
  assign n1874 = n1851 & ~n1857 ;
  assign n1875 = ( ~n1872 & n1873 ) | ( ~n1872 & n1874 ) | ( n1873 & n1874 ) ;
  assign n1876 = n1843 & ~n1875 ;
  assign n1877 = ~n1845 & n1860 ;
  assign n1878 = ( n1861 & ~n1863 ) | ( n1861 & n1877 ) | ( ~n1863 & n1877 ) ;
  assign n1879 = n1220 ^ x96 ^ 1'b0 ;
  assign n1880 = ( x97 & x225 ) | ( x97 & ~n1846 ) | ( x225 & ~n1846 ) ;
  assign n1881 = n1872 & n1876 ;
  assign n1882 = ~n1851 & n1857 ;
  assign n1883 = ( n1849 & ~n1865 ) | ( n1849 & n1882 ) | ( ~n1865 & n1882 ) ;
  assign n1884 = ( ~n1866 & n1867 ) | ( ~n1866 & n1883 ) | ( n1867 & n1883 ) ;
  assign n1885 = ( ~n1868 & n1869 ) | ( ~n1868 & n1884 ) | ( n1869 & n1884 ) ;
  assign n1886 = ( n1876 & ~n1881 ) | ( n1876 & n1885 ) | ( ~n1881 & n1885 ) ;
  assign n1887 = n1202 ^ x353 ^ 1'b0 ;
  assign n1888 = ~n1878 & n1886 ;
  assign n1889 = ( x96 & x224 ) | ( x96 & ~n1879 ) | ( x224 & ~n1879 ) ;
  assign n1890 = n1202 ^ x352 ^ 1'b0 ;
  assign n1891 = ( x352 & x480 ) | ( x352 & ~n1890 ) | ( x480 & ~n1890 ) ;
  assign n1892 = ( x353 & x481 ) | ( x353 & ~n1887 ) | ( x481 & ~n1887 ) ;
  assign n1893 = n1880 & n1892 ;
  assign n1894 = ( n1888 & ~n1892 ) | ( n1888 & n1893 ) | ( ~n1892 & n1893 ) ;
  assign n1895 = n1889 & n1891 ;
  assign n1896 = ( ~n1891 & n1894 ) | ( ~n1891 & n1895 ) | ( n1894 & n1895 ) ;
  assign n1897 = n1889 & ~n1891 ;
  assign n1898 = ( n1880 & ~n1892 ) | ( n1880 & n1897 ) | ( ~n1892 & n1897 ) ;
  assign n1899 = ( n1859 & ~n1861 ) | ( n1859 & n1898 ) | ( ~n1861 & n1898 ) ;
  assign n1900 = ( n1845 & ~n1860 ) | ( n1845 & n1899 ) | ( ~n1860 & n1899 ) ;
  assign n1901 = n1896 | n1900 ;
  assign n1902 = n1202 ^ x362 ^ 1'b0 ;
  assign n1903 = ( x362 & x490 ) | ( x362 & ~n1902 ) | ( x490 & ~n1902 ) ;
  assign n1904 = n1220 ^ x107 ^ 1'b0 ;
  assign n1905 = ( x107 & x235 ) | ( x107 & ~n1904 ) | ( x235 & ~n1904 ) ;
  assign n1906 = n1202 ^ x363 ^ 1'b0 ;
  assign n1907 = ( x363 & x491 ) | ( x363 & ~n1906 ) | ( x491 & ~n1906 ) ;
  assign n1908 = ~n1905 & n1907 ;
  assign n1909 = n1220 ^ x106 ^ 1'b0 ;
  assign n1910 = ( x106 & x234 ) | ( x106 & ~n1909 ) | ( x234 & ~n1909 ) ;
  assign n1911 = n1903 & n1910 ;
  assign n1912 = ( n1903 & n1908 ) | ( n1903 & ~n1911 ) | ( n1908 & ~n1911 ) ;
  assign n1913 = n1220 ^ x105 ^ 1'b0 ;
  assign n1914 = ( x105 & x233 ) | ( x105 & ~n1913 ) | ( x233 & ~n1913 ) ;
  assign n1915 = n1202 ^ x361 ^ 1'b0 ;
  assign n1916 = ( x361 & x489 ) | ( x361 & ~n1915 ) | ( x489 & ~n1915 ) ;
  assign n1917 = ~n1914 & n1916 ;
  assign n1918 = n1202 ^ x360 ^ 1'b0 ;
  assign n1919 = ( x360 & x488 ) | ( x360 & ~n1918 ) | ( x488 & ~n1918 ) ;
  assign n1920 = n1220 ^ x104 ^ 1'b0 ;
  assign n1921 = ( x104 & x232 ) | ( x104 & ~n1920 ) | ( x232 & ~n1920 ) ;
  assign n1922 = n1919 & ~n1921 ;
  assign n1923 = ( ~n1912 & n1917 ) | ( ~n1912 & n1922 ) | ( n1917 & n1922 ) ;
  assign n1924 = n1220 ^ x101 ^ 1'b0 ;
  assign n1925 = ( x101 & x229 ) | ( x101 & ~n1924 ) | ( x229 & ~n1924 ) ;
  assign n1926 = n1202 ^ x357 ^ 1'b0 ;
  assign n1927 = ( x357 & x485 ) | ( x357 & ~n1926 ) | ( x485 & ~n1926 ) ;
  assign n1928 = ~n1925 & n1927 ;
  assign n1929 = n1220 ^ x100 ^ 1'b0 ;
  assign n1930 = ( x100 & x228 ) | ( x100 & ~n1929 ) | ( x228 & ~n1929 ) ;
  assign n1931 = n1202 ^ x356 ^ 1'b0 ;
  assign n1932 = ( x356 & x484 ) | ( x356 & ~n1931 ) | ( x484 & ~n1931 ) ;
  assign n1933 = ~n1930 & n1932 ;
  assign n1934 = n1220 ^ x103 ^ 1'b0 ;
  assign n1935 = ( x103 & x231 ) | ( x103 & ~n1934 ) | ( x231 & ~n1934 ) ;
  assign n1936 = n1202 ^ x359 ^ 1'b0 ;
  assign n1937 = ( x359 & x487 ) | ( x359 & ~n1936 ) | ( x487 & ~n1936 ) ;
  assign n1938 = ~n1935 & n1937 ;
  assign n1939 = n1220 ^ x102 ^ 1'b0 ;
  assign n1940 = ( x102 & x230 ) | ( x102 & ~n1939 ) | ( x230 & ~n1939 ) ;
  assign n1941 = n1202 ^ x358 ^ 1'b0 ;
  assign n1942 = ( x358 & x486 ) | ( x358 & ~n1941 ) | ( x486 & ~n1941 ) ;
  assign n1943 = n1938 | n1942 ;
  assign n1944 = ( n1938 & ~n1940 ) | ( n1938 & n1943 ) | ( ~n1940 & n1943 ) ;
  assign n1945 = ( n1928 & n1933 ) | ( n1928 & ~n1944 ) | ( n1933 & ~n1944 ) ;
  assign n1946 = n1901 & ~n1945 ;
  assign n1947 = n1930 & ~n1932 ;
  assign n1948 = ( n1925 & ~n1927 ) | ( n1925 & n1947 ) | ( ~n1927 & n1947 ) ;
  assign n1949 = ( n1940 & ~n1942 ) | ( n1940 & n1948 ) | ( ~n1942 & n1948 ) ;
  assign n1950 = ( n1935 & ~n1937 ) | ( n1935 & n1949 ) | ( ~n1937 & n1949 ) ;
  assign n1951 = n1944 & n1946 ;
  assign n1952 = ( n1946 & n1950 ) | ( n1946 & ~n1951 ) | ( n1950 & ~n1951 ) ;
  assign n1953 = ( ~n1912 & n1923 ) | ( ~n1912 & n1952 ) | ( n1923 & n1952 ) ;
  assign n1954 = ~n1919 & n1921 ;
  assign n1955 = ( n1914 & ~n1916 ) | ( n1914 & n1954 ) | ( ~n1916 & n1954 ) ;
  assign n1956 = ( ~n1903 & n1910 ) | ( ~n1903 & n1955 ) | ( n1910 & n1955 ) ;
  assign n1957 = ( n1905 & ~n1907 ) | ( n1905 & n1956 ) | ( ~n1907 & n1956 ) ;
  assign n1958 = n1923 & n1953 ;
  assign n1959 = ( n1953 & n1957 ) | ( n1953 & ~n1958 ) | ( n1957 & ~n1958 ) ;
  assign n1960 = n1220 ^ x111 ^ 1'b0 ;
  assign n1961 = ( x111 & x239 ) | ( x111 & ~n1960 ) | ( x239 & ~n1960 ) ;
  assign n1962 = n1202 ^ x367 ^ 1'b0 ;
  assign n1963 = ( x367 & x495 ) | ( x367 & ~n1962 ) | ( x495 & ~n1962 ) ;
  assign n1964 = ~n1961 & n1963 ;
  assign n1965 = n1220 ^ x110 ^ 1'b0 ;
  assign n1966 = ( x110 & x238 ) | ( x110 & ~n1965 ) | ( x238 & ~n1965 ) ;
  assign n1967 = n1202 ^ x366 ^ 1'b0 ;
  assign n1968 = ( x366 & x494 ) | ( x366 & ~n1967 ) | ( x494 & ~n1967 ) ;
  assign n1969 = n1964 | n1968 ;
  assign n1970 = ( n1964 & ~n1966 ) | ( n1964 & n1969 ) | ( ~n1966 & n1969 ) ;
  assign n1971 = n1220 ^ x116 ^ 1'b0 ;
  assign n1972 = ( x116 & x244 ) | ( x116 & ~n1971 ) | ( x244 & ~n1971 ) ;
  assign n1973 = n1220 ^ x119 ^ 1'b0 ;
  assign n1974 = n1202 ^ x371 ^ 1'b0 ;
  assign n1975 = ( x371 & x499 ) | ( x371 & ~n1974 ) | ( x499 & ~n1974 ) ;
  assign n1976 = n1220 ^ x114 ^ 1'b0 ;
  assign n1977 = n1220 ^ x115 ^ 1'b0 ;
  assign n1978 = n1202 ^ x372 ^ 1'b0 ;
  assign n1979 = ( x115 & x243 ) | ( x115 & ~n1977 ) | ( x243 & ~n1977 ) ;
  assign n1980 = n1202 ^ x370 ^ 1'b0 ;
  assign n1981 = ( x114 & x242 ) | ( x114 & ~n1976 ) | ( x242 & ~n1976 ) ;
  assign n1982 = ( x119 & x247 ) | ( x119 & ~n1973 ) | ( x247 & ~n1973 ) ;
  assign n1983 = ( x372 & x500 ) | ( x372 & ~n1978 ) | ( x500 & ~n1978 ) ;
  assign n1984 = ( x370 & x498 ) | ( x370 & ~n1980 ) | ( x498 & ~n1980 ) ;
  assign n1985 = n1975 & ~n1979 ;
  assign n1986 = n1202 ^ x365 ^ 1'b0 ;
  assign n1987 = n1220 ^ x109 ^ 1'b0 ;
  assign n1988 = ( x365 & x493 ) | ( x365 & ~n1986 ) | ( x493 & ~n1986 ) ;
  assign n1989 = n1202 ^ x375 ^ 1'b0 ;
  assign n1990 = ( x109 & x237 ) | ( x109 & ~n1987 ) | ( x237 & ~n1987 ) ;
  assign n1991 = ( x375 & x503 ) | ( x375 & ~n1989 ) | ( x503 & ~n1989 ) ;
  assign n1992 = n1220 ^ x113 ^ 1'b0 ;
  assign n1993 = ( x113 & x241 ) | ( x113 & ~n1992 ) | ( x241 & ~n1992 ) ;
  assign n1994 = n1202 ^ x369 ^ 1'b0 ;
  assign n1995 = ~n1982 & n1991 ;
  assign n1996 = ( x369 & x497 ) | ( x369 & ~n1994 ) | ( x497 & ~n1994 ) ;
  assign n1997 = n1993 & n1996 ;
  assign n1998 = n1988 & ~n1990 ;
  assign n1999 = n1202 ^ x374 ^ 1'b0 ;
  assign n2000 = n1202 ^ x364 ^ 1'b0 ;
  assign n2001 = n1220 ^ x108 ^ 1'b0 ;
  assign n2002 = ( x364 & x492 ) | ( x364 & ~n2000 ) | ( x492 & ~n2000 ) ;
  assign n2003 = ( x374 & x502 ) | ( x374 & ~n1999 ) | ( x502 & ~n1999 ) ;
  assign n2004 = ( x108 & x236 ) | ( x108 & ~n2001 ) | ( x236 & ~n2001 ) ;
  assign n2005 = n2002 & ~n2004 ;
  assign n2006 = ~n2002 & n2004 ;
  assign n2007 = ( ~n1970 & n1998 ) | ( ~n1970 & n2005 ) | ( n1998 & n2005 ) ;
  assign n2008 = ( ~n1988 & n1990 ) | ( ~n1988 & n2006 ) | ( n1990 & n2006 ) ;
  assign n2009 = n1959 & ~n2007 ;
  assign n2010 = ( n1966 & ~n1968 ) | ( n1966 & n2008 ) | ( ~n1968 & n2008 ) ;
  assign n2011 = n1970 & n2009 ;
  assign n2012 = ( n1961 & ~n1963 ) | ( n1961 & n2010 ) | ( ~n1963 & n2010 ) ;
  assign n2013 = ( n2009 & ~n2011 ) | ( n2009 & n2012 ) | ( ~n2011 & n2012 ) ;
  assign n2014 = n1202 ^ x368 ^ 1'b0 ;
  assign n2015 = n1995 | n2003 ;
  assign n2016 = n1981 & n1984 ;
  assign n2017 = ( n1984 & n1985 ) | ( n1984 & ~n2016 ) | ( n1985 & ~n2016 ) ;
  assign n2018 = n1202 ^ x373 ^ 1'b0 ;
  assign n2019 = n2013 & ~n2017 ;
  assign n2020 = ( x368 & x496 ) | ( x368 & ~n2014 ) | ( x496 & ~n2014 ) ;
  assign n2021 = ( ~n1996 & n1997 ) | ( ~n1996 & n2019 ) | ( n1997 & n2019 ) ;
  assign n2022 = n1220 ^ x112 ^ 1'b0 ;
  assign n2023 = ( x112 & x240 ) | ( x112 & ~n2022 ) | ( x240 & ~n2022 ) ;
  assign n2024 = n2020 & n2023 ;
  assign n2025 = ( ~n2020 & n2021 ) | ( ~n2020 & n2024 ) | ( n2021 & n2024 ) ;
  assign n2026 = ~n2020 & n2023 ;
  assign n2027 = ( n1993 & ~n1996 ) | ( n1993 & n2026 ) | ( ~n1996 & n2026 ) ;
  assign n2028 = n1220 ^ x118 ^ 1'b0 ;
  assign n2029 = ( x373 & x501 ) | ( x373 & ~n2018 ) | ( x501 & ~n2018 ) ;
  assign n2030 = ( x118 & x246 ) | ( x118 & ~n2028 ) | ( x246 & ~n2028 ) ;
  assign n2031 = ( n1995 & n2015 ) | ( n1995 & ~n2030 ) | ( n2015 & ~n2030 ) ;
  assign n2032 = n1220 ^ x117 ^ 1'b0 ;
  assign n2033 = ( n1981 & ~n1984 ) | ( n1981 & n2027 ) | ( ~n1984 & n2027 ) ;
  assign n2034 = ( ~n1975 & n1979 ) | ( ~n1975 & n2033 ) | ( n1979 & n2033 ) ;
  assign n2035 = ( x117 & x245 ) | ( x117 & ~n2032 ) | ( x245 & ~n2032 ) ;
  assign n2036 = n2025 | n2034 ;
  assign n2037 = n2029 & ~n2035 ;
  assign n2038 = ~n1972 & n1983 ;
  assign n2039 = ( ~n2031 & n2037 ) | ( ~n2031 & n2038 ) | ( n2037 & n2038 ) ;
  assign n2040 = n1972 & ~n1983 ;
  assign n2041 = n2036 & ~n2039 ;
  assign n2042 = n2031 & n2041 ;
  assign n2043 = ( ~n2029 & n2035 ) | ( ~n2029 & n2040 ) | ( n2035 & n2040 ) ;
  assign n2044 = ( ~n2003 & n2030 ) | ( ~n2003 & n2043 ) | ( n2030 & n2043 ) ;
  assign n2045 = ( n1982 & ~n1991 ) | ( n1982 & n2044 ) | ( ~n1991 & n2044 ) ;
  assign n2046 = ( n2041 & ~n2042 ) | ( n2041 & n2045 ) | ( ~n2042 & n2045 ) ;
  assign n2047 = n1220 ^ x123 ^ 1'b0 ;
  assign n2048 = ( x123 & x251 ) | ( x123 & ~n2047 ) | ( x251 & ~n2047 ) ;
  assign n2049 = n1202 ^ x379 ^ 1'b0 ;
  assign n2050 = ( x379 & x507 ) | ( x379 & ~n2049 ) | ( x507 & ~n2049 ) ;
  assign n2051 = ~n2048 & n2050 ;
  assign n2052 = n1202 ^ x378 ^ 1'b0 ;
  assign n2053 = ( x378 & x506 ) | ( x378 & ~n2052 ) | ( x506 & ~n2052 ) ;
  assign n2054 = n1220 ^ x122 ^ 1'b0 ;
  assign n2055 = ( x122 & x250 ) | ( x122 & ~n2054 ) | ( x250 & ~n2054 ) ;
  assign n2056 = n2053 & n2055 ;
  assign n2057 = ( n2051 & n2053 ) | ( n2051 & ~n2056 ) | ( n2053 & ~n2056 ) ;
  assign n2058 = n1220 ^ x121 ^ 1'b0 ;
  assign n2059 = ( x121 & x249 ) | ( x121 & ~n2058 ) | ( x249 & ~n2058 ) ;
  assign n2060 = n1202 ^ x377 ^ 1'b0 ;
  assign n2061 = ( x377 & x505 ) | ( x377 & ~n2060 ) | ( x505 & ~n2060 ) ;
  assign n2062 = ~n2059 & n2061 ;
  assign n2063 = n1202 ^ x376 ^ 1'b0 ;
  assign n2064 = ( x376 & x504 ) | ( x376 & ~n2063 ) | ( x504 & ~n2063 ) ;
  assign n2065 = n1220 ^ x120 ^ 1'b0 ;
  assign n2066 = ( x120 & x248 ) | ( x120 & ~n2065 ) | ( x248 & ~n2065 ) ;
  assign n2067 = n2064 & ~n2066 ;
  assign n2068 = ( ~n2057 & n2062 ) | ( ~n2057 & n2067 ) | ( n2062 & n2067 ) ;
  assign n2069 = ( n2046 & ~n2057 ) | ( n2046 & n2068 ) | ( ~n2057 & n2068 ) ;
  assign n2070 = ~n2064 & n2066 ;
  assign n2071 = ( n2059 & ~n2061 ) | ( n2059 & n2070 ) | ( ~n2061 & n2070 ) ;
  assign n2072 = ( ~n2053 & n2055 ) | ( ~n2053 & n2071 ) | ( n2055 & n2071 ) ;
  assign n2073 = ( n2048 & ~n2050 ) | ( n2048 & n2072 ) | ( ~n2050 & n2072 ) ;
  assign n2074 = n2068 & n2069 ;
  assign n2075 = ( n2069 & n2073 ) | ( n2069 & ~n2074 ) | ( n2073 & ~n2074 ) ;
  assign n2076 = n1323 & n2075 ;
  assign n2077 = ( n1333 & n2075 ) | ( n1333 & ~n2076 ) | ( n2075 & ~n2076 ) ;
  assign n2078 = n2077 ^ n1406 ^ 1'b0 ;
  assign n2079 = ( n1395 & n1406 ) | ( n1395 & ~n2078 ) | ( n1406 & ~n2078 ) ;
  assign n2080 = n2077 ^ n1405 ^ 1'b0 ;
  assign n2081 = ( n1405 & n1413 ) | ( n1405 & ~n2080 ) | ( n1413 & ~n2080 ) ;
  assign n2082 = n2077 ^ n1404 ^ 1'b0 ;
  assign n2083 = ( n1404 & n1412 ) | ( n1404 & ~n2082 ) | ( n1412 & ~n2082 ) ;
  assign n2084 = n2077 ^ n1775 ^ 1'b0 ;
  assign n2085 = ( n1765 & n1775 ) | ( n1765 & ~n2084 ) | ( n1775 & ~n2084 ) ;
  assign n2086 = n2077 ^ n2059 ^ 1'b0 ;
  assign n2087 = ( n2059 & n2061 ) | ( n2059 & ~n2086 ) | ( n2061 & ~n2086 ) ;
  assign n2088 = n2077 ^ n2048 ^ 1'b0 ;
  assign n2089 = ( n2048 & n2050 ) | ( n2048 & ~n2088 ) | ( n2050 & ~n2088 ) ;
  assign n2090 = ( n1210 & ~n1323 ) | ( n1210 & n2075 ) | ( ~n1323 & n2075 ) ;
  assign n2091 = n1209 & n1210 ;
  assign n2092 = ( n1209 & n2090 ) | ( n1209 & n2091 ) | ( n2090 & n2091 ) ;
  assign n2093 = n2077 ^ n1407 ^ 1'b0 ;
  assign n2094 = ( n1401 & n1407 ) | ( n1401 & ~n2093 ) | ( n1407 & ~n2093 ) ;
  assign n2095 = n2077 ^ n1402 ^ 1'b0 ;
  assign n2096 = n2077 ^ n1409 ^ 1'b0 ;
  assign n2097 = ( n1409 & n1417 ) | ( n1409 & ~n2096 ) | ( n1417 & ~n2096 ) ;
  assign n2098 = n2077 ^ n1426 ^ 1'b0 ;
  assign n2099 = ( n1418 & n1426 ) | ( n1418 & ~n2098 ) | ( n1426 & ~n2098 ) ;
  assign n2100 = n2077 ^ n1423 ^ 1'b0 ;
  assign n2101 = ( n1423 & n1424 ) | ( n1423 & ~n2100 ) | ( n1424 & ~n2100 ) ;
  assign n2102 = n2077 ^ n1425 ^ 1'b0 ;
  assign n2103 = ( n1425 & n1427 ) | ( n1425 & ~n2102 ) | ( n1427 & ~n2102 ) ;
  assign n2104 = n2077 ^ n1437 ^ 1'b0 ;
  assign n2105 = ( n1433 & n1437 ) | ( n1433 & ~n2104 ) | ( n1437 & ~n2104 ) ;
  assign n2106 = n2077 ^ n1471 ^ 1'b0 ;
  assign n2107 = ( n1402 & n1421 ) | ( n1402 & ~n2095 ) | ( n1421 & ~n2095 ) ;
  assign n2108 = ( n1463 & n1471 ) | ( n1463 & ~n2106 ) | ( n1471 & ~n2106 ) ;
  assign n2109 = n2077 ^ n1461 ^ 1'b0 ;
  assign n2110 = ( n1442 & n1461 ) | ( n1442 & ~n2109 ) | ( n1461 & ~n2109 ) ;
  assign n2111 = n2077 ^ n1506 ^ 1'b0 ;
  assign n2112 = ( n1504 & n1506 ) | ( n1504 & ~n2111 ) | ( n1506 & ~n2111 ) ;
  assign n2113 = n2077 ^ n1529 ^ 1'b0 ;
  assign n2114 = ( n1517 & n1529 ) | ( n1517 & ~n2113 ) | ( n1529 & ~n2113 ) ;
  assign n2115 = n2077 ^ n1337 ^ 1'b0 ;
  assign n2116 = ( n1337 & n1339 ) | ( n1337 & ~n2115 ) | ( n1339 & ~n2115 ) ;
  assign n2117 = n2077 ^ n1570 ^ 1'b0 ;
  assign n2118 = ( n1563 & n1570 ) | ( n1563 & ~n2117 ) | ( n1570 & ~n2117 ) ;
  assign n2119 = n2077 ^ n1749 ^ 1'b0 ;
  assign n2120 = ( n1749 & n1756 ) | ( n1749 & ~n2119 ) | ( n1756 & ~n2119 ) ;
  assign n2121 = n2077 ^ n1804 ^ 1'b0 ;
  assign n2122 = ( n1804 & n1811 ) | ( n1804 & ~n2121 ) | ( n1811 & ~n2121 ) ;
  assign n2123 = n2077 ^ n1829 ^ 1'b0 ;
  assign n2124 = ( n1829 & n1830 ) | ( n1829 & ~n2123 ) | ( n1830 & ~n2123 ) ;
  assign n2125 = n2077 ^ n1849 ^ 1'b0 ;
  assign n2126 = ( n1849 & n1865 ) | ( n1849 & ~n2125 ) | ( n1865 & ~n2125 ) ;
  assign n2127 = n2077 ^ n1880 ^ 1'b0 ;
  assign n2128 = ( n1880 & n1892 ) | ( n1880 & ~n2127 ) | ( n1892 & ~n2127 ) ;
  assign n2129 = n2077 ^ n1925 ^ 1'b0 ;
  assign n2130 = ( n1925 & n1927 ) | ( n1925 & ~n2129 ) | ( n1927 & ~n2129 ) ;
  assign n2131 = n2077 ^ n1914 ^ 1'b0 ;
  assign n2132 = ( n1914 & n1916 ) | ( n1914 & ~n2131 ) | ( n1916 & ~n2131 ) ;
  assign n2133 = n2077 ^ n1429 ^ 1'b0 ;
  assign n2134 = ( n1419 & n1429 ) | ( n1419 & ~n2133 ) | ( n1429 & ~n2133 ) ;
  assign n2135 = n2077 ^ n1466 ^ 1'b0 ;
  assign n2136 = ( n1457 & n1466 ) | ( n1457 & ~n2135 ) | ( n1466 & ~n2135 ) ;
  assign n2137 = n2077 ^ n1472 ^ 1'b0 ;
  assign n2138 = n2077 ^ n1450 ^ 1'b0 ;
  assign n2139 = ( n1450 & n1451 ) | ( n1450 & ~n2138 ) | ( n1451 & ~n2138 ) ;
  assign n2140 = n2077 ^ n1452 ^ 1'b0 ;
  assign n2141 = ( n1452 & n1475 ) | ( n1452 & ~n2140 ) | ( n1475 & ~n2140 ) ;
  assign n2142 = n2077 ^ n1468 ^ 1'b0 ;
  assign n2143 = ( n1468 & n1482 ) | ( n1468 & ~n2142 ) | ( n1482 & ~n2142 ) ;
  assign n2144 = n2077 ^ n1460 ^ 1'b0 ;
  assign n2145 = ( n1447 & n1460 ) | ( n1447 & ~n2144 ) | ( n1460 & ~n2144 ) ;
  assign n2146 = n2077 ^ n1454 ^ 1'b0 ;
  assign n2147 = ( n1454 & n1478 ) | ( n1454 & ~n2146 ) | ( n1478 & ~n2146 ) ;
  assign n2148 = n2077 ^ n1476 ^ 1'b0 ;
  assign n2149 = ( n1464 & n1476 ) | ( n1464 & ~n2148 ) | ( n1476 & ~n2148 ) ;
  assign n2150 = n2077 ^ n1503 ^ 1'b0 ;
  assign n2151 = ( n1503 & n1521 ) | ( n1503 & ~n2150 ) | ( n1521 & ~n2150 ) ;
  assign n2152 = n2077 ^ n1369 ^ 1'b0 ;
  assign n2153 = ( n1367 & n1369 ) | ( n1367 & ~n2152 ) | ( n1369 & ~n2152 ) ;
  assign n2154 = n2077 ^ n1352 ^ 1'b0 ;
  assign n2155 = ( n1352 & n1354 ) | ( n1352 & ~n2154 ) | ( n1354 & ~n2154 ) ;
  assign n2156 = n2077 ^ n1302 ^ 1'b0 ;
  assign n2157 = ( n1446 & n1472 ) | ( n1446 & ~n2137 ) | ( n1472 & ~n2137 ) ;
  assign n2158 = ( n1302 & n1324 ) | ( n1302 & ~n2156 ) | ( n1324 & ~n2156 ) ;
  assign n2159 = n2077 ^ n1583 ^ 1'b0 ;
  assign n2160 = ( n1582 & n1583 ) | ( n1582 & ~n2159 ) | ( n1583 & ~n2159 ) ;
  assign n2161 = n2077 ^ n1560 ^ 1'b0 ;
  assign n2162 = ( n1559 & n1560 ) | ( n1559 & ~n2161 ) | ( n1560 & ~n2161 ) ;
  assign n2163 = n2077 ^ n1249 ^ 1'b0 ;
  assign n2164 = ( n1249 & n1261 ) | ( n1249 & ~n2163 ) | ( n1261 & ~n2163 ) ;
  assign n2165 = n2077 ^ n1240 ^ 1'b0 ;
  assign n2166 = ( n1240 & n1254 ) | ( n1240 & ~n2165 ) | ( n1254 & ~n2165 ) ;
  assign n2167 = n2077 ^ n1224 ^ 1'b0 ;
  assign n2168 = ( n1224 & n1227 ) | ( n1224 & ~n2167 ) | ( n1227 & ~n2167 ) ;
  assign n2169 = n2077 ^ n1232 ^ 1'b0 ;
  assign n2170 = ( n1232 & n1234 ) | ( n1232 & ~n2169 ) | ( n1234 & ~n2169 ) ;
  assign n2171 = n2077 ^ n1616 ^ 1'b0 ;
  assign n2172 = ( n1616 & n1619 ) | ( n1616 & ~n2171 ) | ( n1619 & ~n2171 ) ;
  assign n2173 = n2077 ^ n1682 ^ 1'b0 ;
  assign n2174 = ( n1681 & n1682 ) | ( n1681 & ~n2173 ) | ( n1682 & ~n2173 ) ;
  assign n2175 = n2077 ^ n1676 ^ 1'b0 ;
  assign n2176 = ( n1675 & n1676 ) | ( n1675 & ~n2175 ) | ( n1676 & ~n2175 ) ;
  assign n2177 = n2077 ^ n1697 ^ 1'b0 ;
  assign n2178 = ( n1670 & n1697 ) | ( n1670 & ~n2177 ) | ( n1697 & ~n2177 ) ;
  assign n2179 = n2077 ^ n1672 ^ 1'b0 ;
  assign n2180 = ( n1672 & n1695 ) | ( n1672 & ~n2179 ) | ( n1695 & ~n2179 ) ;
  assign n2181 = n2077 ^ n1734 ^ 1'b0 ;
  assign n2182 = ( n1734 & n1745 ) | ( n1734 & ~n2181 ) | ( n1745 & ~n2181 ) ;
  assign n2183 = n2077 ^ n1768 ^ 1'b0 ;
  assign n2184 = ( n1766 & n1768 ) | ( n1766 & ~n2183 ) | ( n1768 & ~n2183 ) ;
  assign n2185 = n2077 ^ n1795 ^ 1'b0 ;
  assign n2186 = ( n1790 & n1795 ) | ( n1790 & ~n2185 ) | ( n1795 & ~n2185 ) ;
  assign n2187 = n2077 ^ n1818 ^ 1'b0 ;
  assign n2188 = ( n1818 & n1823 ) | ( n1818 & ~n2187 ) | ( n1823 & ~n2187 ) ;
  assign n2189 = n2077 ^ n1869 ^ 1'b0 ;
  assign n2190 = ( n1868 & n1869 ) | ( n1868 & ~n2189 ) | ( n1869 & ~n2189 ) ;
  assign n2191 = n2077 ^ n1845 ^ 1'b0 ;
  assign n2192 = ( n1845 & n1860 ) | ( n1845 & ~n2191 ) | ( n1860 & ~n2191 ) ;
  assign n2193 = n2077 ^ n1935 ^ 1'b0 ;
  assign n2194 = ( n1935 & n1937 ) | ( n1935 & ~n2193 ) | ( n1937 & ~n2193 ) ;
  assign n2195 = n2077 ^ n1905 ^ 1'b0 ;
  assign n2196 = ( n1905 & n1907 ) | ( n1905 & ~n2195 ) | ( n1907 & ~n2195 ) ;
  assign n2197 = n2077 ^ n1990 ^ 1'b0 ;
  assign n2198 = ( n1988 & n1990 ) | ( n1988 & ~n2197 ) | ( n1990 & ~n2197 ) ;
  assign n2199 = n2077 ^ n1961 ^ 1'b0 ;
  assign n2200 = ( n1961 & n1963 ) | ( n1961 & ~n2199 ) | ( n1963 & ~n2199 ) ;
  assign n2201 = n2077 ^ n1993 ^ 1'b0 ;
  assign n2202 = ( n1993 & n1996 ) | ( n1993 & ~n2201 ) | ( n1996 & ~n2201 ) ;
  assign n2203 = n2077 ^ n2055 ^ 1'b0 ;
  assign n2204 = ( n2053 & n2055 ) | ( n2053 & ~n2203 ) | ( n2055 & ~n2203 ) ;
  assign n2205 = n2077 ^ n1501 ^ 1'b0 ;
  assign n2206 = ( n1501 & n1509 ) | ( n1501 & ~n2205 ) | ( n1509 & ~n2205 ) ;
  assign n2207 = n2077 ^ n1519 ^ 1'b0 ;
  assign n2208 = ( n1496 & n1519 ) | ( n1496 & ~n2207 ) | ( n1519 & ~n2207 ) ;
  assign n2209 = n2077 ^ n1526 ^ 1'b0 ;
  assign n2210 = n2077 ^ n1531 ^ 1'b0 ;
  assign n2211 = ( n1502 & n1531 ) | ( n1502 & ~n2210 ) | ( n1531 & ~n2210 ) ;
  assign n2212 = n2077 ^ n1515 ^ 1'b0 ;
  assign n2213 = ( n1511 & n1515 ) | ( n1511 & ~n2212 ) | ( n1515 & ~n2212 ) ;
  assign n2214 = n2077 ^ n1537 ^ 1'b0 ;
  assign n2215 = ( n1537 & n1538 ) | ( n1537 & ~n2214 ) | ( n1538 & ~n2214 ) ;
  assign n2216 = n2077 ^ n1533 ^ 1'b0 ;
  assign n2217 = ( n1533 & n1534 ) | ( n1533 & ~n2216 ) | ( n1534 & ~n2216 ) ;
  assign n2218 = n2077 ^ n1544 ^ 1'b0 ;
  assign n2219 = ( n1535 & n1544 ) | ( n1535 & ~n2218 ) | ( n1544 & ~n2218 ) ;
  assign n2220 = n2077 ^ n1371 ^ 1'b0 ;
  assign n2221 = ( n1335 & n1371 ) | ( n1335 & ~n2220 ) | ( n1371 & ~n2220 ) ;
  assign n2222 = n2077 ^ n1359 ^ 1'b0 ;
  assign n2223 = ( n1359 & n1361 ) | ( n1359 & ~n2222 ) | ( n1361 & ~n2222 ) ;
  assign n2224 = n2077 ^ n1363 ^ 1'b0 ;
  assign n2225 = ( n1363 & n1365 ) | ( n1363 & ~n2224 ) | ( n1365 & ~n2224 ) ;
  assign n2226 = n2077 ^ n1347 ^ 1'b0 ;
  assign n2227 = ( n1347 & n1349 ) | ( n1347 & ~n2226 ) | ( n1349 & ~n2226 ) ;
  assign n2228 = n2077 ^ n1238 ^ 1'b0 ;
  assign n2229 = ( n1493 & n1526 ) | ( n1493 & ~n2209 ) | ( n1526 & ~n2209 ) ;
  assign n2230 = ( n1238 & n1251 ) | ( n1238 & ~n2228 ) | ( n1251 & ~n2228 ) ;
  assign n2231 = n2077 ^ n1236 ^ 1'b0 ;
  assign n2232 = ( n1235 & n1236 ) | ( n1235 & ~n2231 ) | ( n1236 & ~n2231 ) ;
  assign n2233 = n2077 ^ n1614 ^ 1'b0 ;
  assign n2234 = ( n1614 & n1618 ) | ( n1614 & ~n2233 ) | ( n1618 & ~n2233 ) ;
  assign n2235 = n2077 ^ n1628 ^ 1'b0 ;
  assign n2236 = ( n1628 & n1629 ) | ( n1628 & ~n2235 ) | ( n1629 & ~n2235 ) ;
  assign n2237 = n2077 ^ n1281 ^ 1'b0 ;
  assign n2238 = ( n1281 & n1293 ) | ( n1281 & ~n2237 ) | ( n1293 & ~n2237 ) ;
  assign n2239 = n2077 ^ n1276 ^ 1'b0 ;
  assign n2240 = ( n1276 & n1287 ) | ( n1276 & ~n2239 ) | ( n1287 & ~n2239 ) ;
  assign n2241 = n2077 ^ n1685 ^ 1'b0 ;
  assign n2242 = ( n1663 & n1685 ) | ( n1663 & ~n2241 ) | ( n1685 & ~n2241 ) ;
  assign n2243 = n2077 ^ n1690 ^ 1'b0 ;
  assign n2244 = ( n1690 & n1699 ) | ( n1690 & ~n2243 ) | ( n1699 & ~n2243 ) ;
  assign n2245 = n2077 ^ n1742 ^ 1'b0 ;
  assign n2246 = ( n1742 & n1744 ) | ( n1742 & ~n2245 ) | ( n1744 & ~n2245 ) ;
  assign n2247 = n2077 ^ n1751 ^ 1'b0 ;
  assign n2248 = ( n1751 & n1769 ) | ( n1751 & ~n2247 ) | ( n1769 & ~n2247 ) ;
  assign n2249 = n2077 ^ n1813 ^ 1'b0 ;
  assign n2250 = ( n1793 & n1813 ) | ( n1793 & ~n2249 ) | ( n1813 & ~n2249 ) ;
  assign n2251 = n2077 ^ n1799 ^ 1'b0 ;
  assign n2252 = ( n1796 & n1799 ) | ( n1796 & ~n2251 ) | ( n1799 & ~n2251 ) ;
  assign n2253 = n2077 ^ n1867 ^ 1'b0 ;
  assign n2254 = ( n1866 & n1867 ) | ( n1866 & ~n2253 ) | ( n1867 & ~n2253 ) ;
  assign n2255 = n2077 ^ n1859 ^ 1'b0 ;
  assign n2256 = ( n1859 & n1861 ) | ( n1859 & ~n2255 ) | ( n1861 & ~n2255 ) ;
  assign n2257 = n2077 ^ n1940 ^ 1'b0 ;
  assign n2258 = ( n1940 & n1942 ) | ( n1940 & ~n2257 ) | ( n1942 & ~n2257 ) ;
  assign n2259 = n2077 ^ n1910 ^ 1'b0 ;
  assign n2260 = ( n1903 & n1910 ) | ( n1903 & ~n2259 ) | ( n1910 & ~n2259 ) ;
  assign n2261 = n2077 ^ n1966 ^ 1'b0 ;
  assign n2262 = ( n1966 & n1968 ) | ( n1966 & ~n2261 ) | ( n1968 & ~n2261 ) ;
  assign n2263 = n2077 ^ n1981 ^ 1'b0 ;
  assign n2264 = ( n1981 & n1984 ) | ( n1981 & ~n2263 ) | ( n1984 & ~n2263 ) ;
  assign n2265 = n2077 ^ n1982 ^ 1'b0 ;
  assign n2266 = ( n1982 & n1991 ) | ( n1982 & ~n2265 ) | ( n1991 & ~n2265 ) ;
  assign n2267 = n2077 ^ n2066 ^ 1'b0 ;
  assign n2268 = ( n2064 & n2066 ) | ( n2064 & ~n2267 ) | ( n2066 & ~n2267 ) ;
  assign n2269 = n2077 ^ n1308 ^ 1'b0 ;
  assign n2270 = ( n1216 & n1308 ) | ( n1216 & ~n2269 ) | ( n1308 & ~n2269 ) ;
  assign n2271 = n2077 ^ n1315 ^ 1'b0 ;
  assign n2272 = ( n1315 & n1317 ) | ( n1315 & ~n2271 ) | ( n1317 & ~n2271 ) ;
  assign n2273 = n2077 ^ n1312 ^ 1'b0 ;
  assign n2274 = ( n1286 & n1312 ) | ( n1286 & ~n2273 ) | ( n1312 & ~n2273 ) ;
  assign n2275 = n2077 ^ n1220 ^ 1'b0 ;
  assign n2276 = ( n1202 & n1220 ) | ( n1202 & ~n2275 ) | ( n1220 & ~n2275 ) ;
  assign n2277 = n2077 ^ n1342 ^ 1'b0 ;
  assign n2278 = ( n1342 & n1344 ) | ( n1342 & ~n2277 ) | ( n1344 & ~n2277 ) ;
  assign n2279 = n2077 ^ n1579 ^ 1'b0 ;
  assign n2280 = ( n1569 & n1579 ) | ( n1569 & ~n2279 ) | ( n1579 & ~n2279 ) ;
  assign n2281 = n2077 ^ n1303 ^ 1'b0 ;
  assign n2282 = ( n1303 & n1310 ) | ( n1303 & ~n2281 ) | ( n1310 & ~n2281 ) ;
  assign n2283 = n2077 ^ n1585 ^ 1'b0 ;
  assign n2284 = ( n1573 & n1585 ) | ( n1573 & ~n2283 ) | ( n1585 & ~n2283 ) ;
  assign n2285 = n2077 ^ n1564 ^ 1'b0 ;
  assign n2286 = ( n1564 & n1568 ) | ( n1564 & ~n2285 ) | ( n1568 & ~n2285 ) ;
  assign n2287 = n2077 ^ n1246 ^ 1'b0 ;
  assign n2288 = ( n1242 & n1246 ) | ( n1242 & ~n2287 ) | ( n1246 & ~n2287 ) ;
  assign n2289 = n2077 ^ n1222 ^ 1'b0 ;
  assign n2290 = ( n1215 & n1222 ) | ( n1215 & ~n2289 ) | ( n1222 & ~n2289 ) ;
  assign n2291 = n2077 ^ n1633 ^ 1'b0 ;
  assign n2292 = ( n1625 & n1633 ) | ( n1625 & ~n2291 ) | ( n1633 & ~n2291 ) ;
  assign n2293 = n2077 ^ n1295 ^ 1'b0 ;
  assign n2294 = ( n1283 & n1295 ) | ( n1283 & ~n2293 ) | ( n1295 & ~n2293 ) ;
  assign n2295 = n2077 ^ n1291 ^ 1'b0 ;
  assign n2296 = ( n1289 & n1291 ) | ( n1289 & ~n2295 ) | ( n1291 & ~n2295 ) ;
  assign n2297 = n2077 ^ n1653 ^ 1'b0 ;
  assign n2298 = ( n1650 & n1653 ) | ( n1650 & ~n2297 ) | ( n1653 & ~n2297 ) ;
  assign n2299 = n2077 ^ n1651 ^ 1'b0 ;
  assign n2300 = ( n1645 & n1651 ) | ( n1645 & ~n2299 ) | ( n1651 & ~n2299 ) ;
  assign n2301 = n2077 ^ n1693 ^ 1'b0 ;
  assign n2302 = ( n1687 & n1693 ) | ( n1687 & ~n2301 ) | ( n1693 & ~n2301 ) ;
  assign n2303 = n2077 ^ n1706 ^ 1'b0 ;
  assign n2304 = ( n1700 & n1706 ) | ( n1700 & ~n2303 ) | ( n1706 & ~n2303 ) ;
  assign n2305 = n2077 ^ n1665 ^ 1'b0 ;
  assign n2306 = ( n1665 & n1667 ) | ( n1665 & ~n2305 ) | ( n1667 & ~n2305 ) ;
  assign n2307 = n2077 ^ n1713 ^ 1'b0 ;
  assign n2308 = ( n1713 & n1717 ) | ( n1713 & ~n2307 ) | ( n1717 & ~n2307 ) ;
  assign n2309 = n2077 ^ n1740 ^ 1'b0 ;
  assign n2310 = ( n1740 & n1750 ) | ( n1740 & ~n2309 ) | ( n1750 & ~n2309 ) ;
  assign n2311 = n2077 ^ n1753 ^ 1'b0 ;
  assign n2312 = ( n1736 & n1753 ) | ( n1736 & ~n2311 ) | ( n1753 & ~n2311 ) ;
  assign n2313 = n2077 ^ n1808 ^ 1'b0 ;
  assign n2314 = ( n1808 & n1809 ) | ( n1808 & ~n2313 ) | ( n1809 & ~n2313 ) ;
  assign n2315 = n2077 ^ n1824 ^ 1'b0 ;
  assign n2316 = ( n1817 & n1824 ) | ( n1817 & ~n2315 ) | ( n1824 & ~n2315 ) ;
  assign n2317 = n2077 ^ n1857 ^ 1'b0 ;
  assign n2318 = ( n1851 & n1857 ) | ( n1851 & ~n2317 ) | ( n1857 & ~n2317 ) ;
  assign n2319 = n2077 ^ n1889 ^ 1'b0 ;
  assign n2320 = ( n1889 & n1891 ) | ( n1889 & ~n2319 ) | ( n1891 & ~n2319 ) ;
  assign n2321 = n2077 ^ n1930 ^ 1'b0 ;
  assign n2322 = ( n1930 & n1932 ) | ( n1930 & ~n2321 ) | ( n1932 & ~n2321 ) ;
  assign n2323 = n2077 ^ n1921 ^ 1'b0 ;
  assign n2324 = ( n1919 & n1921 ) | ( n1919 & ~n2323 ) | ( n1921 & ~n2323 ) ;
  assign n2325 = n2077 ^ n2004 ^ 1'b0 ;
  assign n2326 = ( n2002 & n2004 ) | ( n2002 & ~n2325 ) | ( n2004 & ~n2325 ) ;
  assign n2327 = n2077 ^ n2023 ^ 1'b0 ;
  assign n2328 = ( n2020 & n2023 ) | ( n2020 & ~n2327 ) | ( n2023 & ~n2327 ) ;
  assign n2329 = n2077 ^ n1979 ^ 1'b0 ;
  assign n2330 = ( n1975 & n1979 ) | ( n1975 & ~n2329 ) | ( n1979 & ~n2329 ) ;
  assign n2331 = n2077 ^ n1972 ^ 1'b0 ;
  assign n2332 = ( n1972 & n1983 ) | ( n1972 & ~n2331 ) | ( n1983 & ~n2331 ) ;
  assign n2333 = n2077 ^ n2035 ^ 1'b0 ;
  assign n2334 = ( n2029 & n2035 ) | ( n2029 & ~n2333 ) | ( n2035 & ~n2333 ) ;
  assign n2335 = n2077 ^ n2030 ^ 1'b0 ;
  assign n2336 = ( n2003 & n2030 ) | ( n2003 & ~n2335 ) | ( n2030 & ~n2335 ) ;
  assign y0 = n2079 ;
  assign y1 = n2081 ;
  assign y2 = n2083 ;
  assign y3 = n2094 ;
  assign y4 = n2107 ;
  assign y5 = n2097 ;
  assign y6 = n2099 ;
  assign y7 = n2101 ;
  assign y8 = n2103 ;
  assign y9 = n2134 ;
  assign y10 = n2105 ;
  assign y11 = n2136 ;
  assign y12 = n2108 ;
  assign y13 = n2157 ;
  assign y14 = n2139 ;
  assign y15 = n2141 ;
  assign y16 = n2143 ;
  assign y17 = n2145 ;
  assign y18 = n2147 ;
  assign y19 = n2110 ;
  assign y20 = n2149 ;
  assign y21 = n2206 ;
  assign y22 = n2112 ;
  assign y23 = n2208 ;
  assign y24 = n2151 ;
  assign y25 = n2229 ;
  assign y26 = n2114 ;
  assign y27 = n2211 ;
  assign y28 = n2213 ;
  assign y29 = n2215 ;
  assign y30 = n2217 ;
  assign y31 = n2219 ;
  assign y32 = n2221 ;
  assign y33 = n2223 ;
  assign y34 = n2153 ;
  assign y35 = n2225 ;
  assign y36 = n2116 ;
  assign y37 = n2278 ;
  assign y38 = n2155 ;
  assign y39 = n2227 ;
  assign y40 = n2118 ;
  assign y41 = n2280 ;
  assign y42 = n2158 ;
  assign y43 = n2282 ;
  assign y44 = n2160 ;
  assign y45 = n2284 ;
  assign y46 = n2162 ;
  assign y47 = n2286 ;
  assign y48 = n2164 ;
  assign y49 = n2230 ;
  assign y50 = n2166 ;
  assign y51 = n2288 ;
  assign y52 = n2168 ;
  assign y53 = n2232 ;
  assign y54 = n2170 ;
  assign y55 = n2290 ;
  assign y56 = n2172 ;
  assign y57 = n2234 ;
  assign y58 = n2292 ;
  assign y59 = n2236 ;
  assign y60 = n2294 ;
  assign y61 = n2238 ;
  assign y62 = n2296 ;
  assign y63 = n2240 ;
  assign y64 = n2298 ;
  assign y65 = n2300 ;
  assign y66 = n2302 ;
  assign y67 = n2304 ;
  assign y68 = n2306 ;
  assign y69 = n2174 ;
  assign y70 = n2242 ;
  assign y71 = n2176 ;
  assign y72 = n2308 ;
  assign y73 = n2178 ;
  assign y74 = n2244 ;
  assign y75 = n2180 ;
  assign y76 = n2310 ;
  assign y77 = n2120 ;
  assign y78 = n2246 ;
  assign y79 = n2182 ;
  assign y80 = n2312 ;
  assign y81 = n2085 ;
  assign y82 = n2248 ;
  assign y83 = n2184 ;
  assign y84 = n2314 ;
  assign y85 = n2122 ;
  assign y86 = n2250 ;
  assign y87 = n2186 ;
  assign y88 = n2316 ;
  assign y89 = n2124 ;
  assign y90 = n2252 ;
  assign y91 = n2188 ;
  assign y92 = n2318 ;
  assign y93 = n2126 ;
  assign y94 = n2254 ;
  assign y95 = n2190 ;
  assign y96 = n2320 ;
  assign y97 = n2128 ;
  assign y98 = n2256 ;
  assign y99 = n2192 ;
  assign y100 = n2322 ;
  assign y101 = n2130 ;
  assign y102 = n2258 ;
  assign y103 = n2194 ;
  assign y104 = n2324 ;
  assign y105 = n2132 ;
  assign y106 = n2260 ;
  assign y107 = n2196 ;
  assign y108 = n2326 ;
  assign y109 = n2198 ;
  assign y110 = n2262 ;
  assign y111 = n2200 ;
  assign y112 = n2328 ;
  assign y113 = n2202 ;
  assign y114 = n2264 ;
  assign y115 = n2330 ;
  assign y116 = n2332 ;
  assign y117 = n2334 ;
  assign y118 = n2336 ;
  assign y119 = n2266 ;
  assign y120 = n2268 ;
  assign y121 = n2087 ;
  assign y122 = n2204 ;
  assign y123 = n2089 ;
  assign y124 = n2270 ;
  assign y125 = n2272 ;
  assign y126 = n2274 ;
  assign y127 = n2092 ;
  assign y128 = ~n2276 ;
  assign y129 = ~n2077 ;
endmodule
