module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 ;
  assign n129 = x124 | x125 ;
  assign n130 = x122 | x123 ;
  assign n131 = x126 | x127 ;
  assign n132 = ~n129 & n130 ;
  assign n133 = n131 | n132 ;
  assign n134 = ( x122 & ~x123 ) | ( x122 & x124 ) | ( ~x123 & x124 ) ;
  assign n135 = ( x124 & ~x125 ) | ( x124 & n134 ) | ( ~x125 & n134 ) ;
  assign n136 = x126 & ~x127 ;
  assign n137 = ( ~x125 & x126 ) | ( ~x125 & n135 ) | ( x126 & n135 ) ;
  assign n138 = ( x121 & n129 ) | ( x121 & ~n132 ) | ( n129 & ~n132 ) ;
  assign n139 = ~n131 & n138 ;
  assign n140 = ( ~x127 & n136 ) | ( ~x127 & n137 ) | ( n136 & n137 ) ;
  assign n141 = n140 ^ n139 ^ n133 ;
  assign n142 = ( x120 & ~n133 ) | ( x120 & n139 ) | ( ~n133 & n139 ) ;
  assign n143 = n141 ^ x119 ^ 1'b0 ;
  assign n144 = n142 ^ n141 ^ n133 ;
  assign n145 = ( n141 & n143 ) | ( n141 & ~n144 ) | ( n143 & ~n144 ) ;
  assign n146 = x118 | x119 ;
  assign n147 = ( n133 & ~n142 ) | ( n133 & n146 ) | ( ~n142 & n146 ) ;
  assign n148 = x116 | x117 ;
  assign n149 = ( n142 & ~n147 ) | ( n142 & n148 ) | ( ~n147 & n148 ) ;
  assign n150 = x114 | x115 ;
  assign n151 = n146 | n148 ;
  assign n152 = n150 ^ n149 ^ 1'b0 ;
  assign n153 = ( n147 & ~n149 ) | ( n147 & n152 ) | ( ~n149 & n152 ) ;
  assign n154 = n147 ^ n145 ^ n142 ;
  assign n155 = n129 | n131 ;
  assign n156 = n145 ^ x117 ^ 1'b0 ;
  assign n157 = ( n145 & ~n154 ) | ( n145 & n156 ) | ( ~n154 & n156 ) ;
  assign n158 = n157 ^ n149 ^ n147 ;
  assign n159 = x112 | x113 ;
  assign n160 = ( ~x120 & x121 ) | ( ~x120 & n130 ) | ( x121 & n130 ) ;
  assign n161 = x120 | n160 ;
  assign n162 = n157 ^ x115 ^ 1'b0 ;
  assign n163 = ( n157 & ~n158 ) | ( n157 & n162 ) | ( ~n158 & n162 ) ;
  assign n164 = n159 ^ n153 ^ 1'b0 ;
  assign n165 = ( n149 & ~n153 ) | ( n149 & n164 ) | ( ~n153 & n164 ) ;
  assign n166 = n163 ^ n153 ^ n149 ;
  assign n167 = n163 ^ x113 ^ 1'b0 ;
  assign n168 = ( n163 & ~n166 ) | ( n163 & n167 ) | ( ~n166 & n167 ) ;
  assign n169 = n151 & ~n161 ;
  assign n170 = ( ~n150 & n151 ) | ( ~n150 & n159 ) | ( n151 & n159 ) ;
  assign n171 = ( x115 & n161 ) | ( x115 & ~n169 ) | ( n161 & ~n169 ) ;
  assign n172 = n155 | n161 ;
  assign n173 = x114 | n159 ;
  assign n174 = n155 | n169 ;
  assign n175 = n150 | n170 ;
  assign n176 = ~n155 & n171 ;
  assign n177 = n168 ^ x111 ^ 1'b0 ;
  assign n178 = n168 ^ n165 ^ n153 ;
  assign n179 = n174 ^ n173 ^ 1'b0 ;
  assign n180 = ( n168 & n177 ) | ( n168 & ~n178 ) | ( n177 & ~n178 ) ;
  assign n181 = n180 ^ x109 ^ 1'b0 ;
  assign n182 = x110 | x111 ;
  assign n183 = ( ~n174 & n176 ) | ( ~n174 & n179 ) | ( n176 & n179 ) ;
  assign n184 = n182 ^ n165 ^ 1'b0 ;
  assign n185 = ( n153 & ~n165 ) | ( n153 & n184 ) | ( ~n165 & n184 ) ;
  assign n186 = n185 ^ n180 ^ n165 ;
  assign n187 = ( n180 & n181 ) | ( n180 & ~n186 ) | ( n181 & ~n186 ) ;
  assign n188 = x108 | x109 ;
  assign n189 = x106 | x107 ;
  assign n190 = n188 ^ n185 ^ 1'b0 ;
  assign n191 = ( n165 & ~n185 ) | ( n165 & n190 ) | ( ~n185 & n190 ) ;
  assign n192 = n191 ^ n189 ^ 1'b0 ;
  assign n193 = ( n185 & ~n191 ) | ( n185 & n192 ) | ( ~n191 & n192 ) ;
  assign n194 = n187 ^ x107 ^ 1'b0 ;
  assign n195 = n191 ^ n187 ^ n185 ;
  assign n196 = x104 | x105 ;
  assign n197 = n189 | n196 ;
  assign n198 = n196 ^ n193 ^ 1'b0 ;
  assign n199 = ( n187 & n194 ) | ( n187 & ~n195 ) | ( n194 & ~n195 ) ;
  assign n200 = n199 ^ n193 ^ n191 ;
  assign n201 = n199 ^ x105 ^ 1'b0 ;
  assign n202 = ( n191 & ~n193 ) | ( n191 & n198 ) | ( ~n193 & n198 ) ;
  assign n203 = x102 | x103 ;
  assign n204 = ( n199 & ~n200 ) | ( n199 & n201 ) | ( ~n200 & n201 ) ;
  assign n205 = x100 | x101 ;
  assign n206 = n203 ^ n202 ^ 1'b0 ;
  assign n207 = ( n193 & ~n202 ) | ( n193 & n206 ) | ( ~n202 & n206 ) ;
  assign n208 = n204 ^ n202 ^ n193 ;
  assign n209 = n182 | n188 ;
  assign n210 = n204 ^ x103 ^ 1'b0 ;
  assign n211 = ( n204 & ~n208 ) | ( n204 & n210 ) | ( ~n208 & n210 ) ;
  assign n212 = n211 ^ x101 ^ 1'b0 ;
  assign n213 = n211 ^ n207 ^ n202 ;
  assign n214 = ( n211 & n212 ) | ( n211 & ~n213 ) | ( n212 & ~n213 ) ;
  assign n215 = n207 ^ n205 ^ 1'b0 ;
  assign n216 = ( n202 & ~n207 ) | ( n202 & n215 ) | ( ~n207 & n215 ) ;
  assign n217 = n214 ^ x99 ^ 1'b0 ;
  assign n218 = ( n174 & ~n183 ) | ( n174 & n209 ) | ( ~n183 & n209 ) ;
  assign n219 = n197 | n209 ;
  assign n220 = x98 | x99 ;
  assign n221 = ( n183 & n197 ) | ( n183 & ~n218 ) | ( n197 & ~n218 ) ;
  assign n222 = n216 ^ n214 ^ n207 ;
  assign n223 = ( n214 & n217 ) | ( n214 & ~n222 ) | ( n217 & ~n222 ) ;
  assign n224 = x96 | x97 ;
  assign n225 = n220 ^ n216 ^ 1'b0 ;
  assign n226 = ( n207 & ~n216 ) | ( n207 & n225 ) | ( ~n216 & n225 ) ;
  assign n227 = n226 ^ n224 ^ 1'b0 ;
  assign n228 = n203 | n205 ;
  assign n229 = n220 | n224 ;
  assign n230 = ( n216 & ~n226 ) | ( n216 & n227 ) | ( ~n226 & n227 ) ;
  assign n231 = ( ~x102 & n205 ) | ( ~x102 & n229 ) | ( n205 & n229 ) ;
  assign n232 = x102 | n231 ;
  assign n233 = n223 ^ x97 ^ 1'b0 ;
  assign n234 = n226 ^ n223 ^ n216 ;
  assign n235 = ( n223 & n233 ) | ( n223 & ~n234 ) | ( n233 & ~n234 ) ;
  assign n236 = n228 ^ n221 ^ 1'b0 ;
  assign n237 = ( n218 & ~n221 ) | ( n218 & n236 ) | ( ~n221 & n236 ) ;
  assign n238 = ~n175 & n219 ;
  assign n239 = ( n219 & ~n228 ) | ( n219 & n229 ) | ( ~n228 & n229 ) ;
  assign n240 = n228 | n239 ;
  assign n241 = n237 ^ n229 ^ 1'b0 ;
  assign n242 = n235 ^ n230 ^ n226 ;
  assign n243 = x94 | x95 ;
  assign n244 = ( n221 & ~n237 ) | ( n221 & n241 ) | ( ~n237 & n241 ) ;
  assign n245 = n235 ^ x95 ^ 1'b0 ;
  assign n246 = ( n235 & ~n242 ) | ( n235 & n245 ) | ( ~n242 & n245 ) ;
  assign n247 = n172 | n238 ;
  assign n248 = n243 ^ n230 ^ 1'b0 ;
  assign n249 = ( n226 & ~n230 ) | ( n226 & n248 ) | ( ~n230 & n248 ) ;
  assign n250 = n172 & ~n238 ;
  assign n251 = n250 ^ n238 ^ n232 ;
  assign n252 = ( x103 & n175 ) | ( x103 & ~n238 ) | ( n175 & ~n238 ) ;
  assign n253 = n172 | n175 ;
  assign n254 = ( ~n238 & n251 ) | ( ~n238 & n252 ) | ( n251 & n252 ) ;
  assign n255 = ~n172 & n254 ;
  assign n256 = n246 ^ x93 ^ 1'b0 ;
  assign n257 = n249 ^ n246 ^ n230 ;
  assign n258 = ( n246 & n256 ) | ( n246 & ~n257 ) | ( n256 & ~n257 ) ;
  assign n259 = x92 | x93 ;
  assign n260 = n259 ^ n249 ^ 1'b0 ;
  assign n261 = n258 ^ x91 ^ 1'b0 ;
  assign n262 = ( n230 & ~n249 ) | ( n230 & n260 ) | ( ~n249 & n260 ) ;
  assign n263 = n262 ^ n258 ^ n249 ;
  assign n264 = ( n258 & n261 ) | ( n258 & ~n263 ) | ( n261 & ~n263 ) ;
  assign n265 = n243 | n259 ;
  assign n266 = x90 | x91 ;
  assign n267 = n266 ^ n262 ^ 1'b0 ;
  assign n268 = ( n249 & ~n262 ) | ( n249 & n267 ) | ( ~n262 & n267 ) ;
  assign n269 = x88 | x89 ;
  assign n270 = n269 ^ n268 ^ 1'b0 ;
  assign n271 = n266 | n269 ;
  assign n272 = ( n262 & ~n268 ) | ( n262 & n270 ) | ( ~n268 & n270 ) ;
  assign n273 = n264 ^ x89 ^ 1'b0 ;
  assign n274 = n268 ^ n264 ^ n262 ;
  assign n275 = ( n264 & n273 ) | ( n264 & ~n274 ) | ( n273 & ~n274 ) ;
  assign n276 = n275 ^ n272 ^ n268 ;
  assign n277 = n275 ^ x87 ^ 1'b0 ;
  assign n278 = ( n275 & ~n276 ) | ( n275 & n277 ) | ( ~n276 & n277 ) ;
  assign n279 = x86 | x87 ;
  assign n280 = n279 ^ n272 ^ 1'b0 ;
  assign n281 = ( n268 & ~n272 ) | ( n268 & n280 ) | ( ~n272 & n280 ) ;
  assign n282 = n265 | n271 ;
  assign n283 = n265 ^ n244 ^ 1'b0 ;
  assign n284 = ( n247 & ~n255 ) | ( n247 & n282 ) | ( ~n255 & n282 ) ;
  assign n285 = ( n237 & ~n244 ) | ( n237 & n283 ) | ( ~n244 & n283 ) ;
  assign n286 = x84 | x85 ;
  assign n287 = n279 | n286 ;
  assign n288 = n286 ^ n281 ^ 1'b0 ;
  assign n289 = n285 ^ n271 ^ 1'b0 ;
  assign n290 = ( n244 & ~n285 ) | ( n244 & n289 ) | ( ~n285 & n289 ) ;
  assign n291 = ( n272 & ~n281 ) | ( n272 & n288 ) | ( ~n281 & n288 ) ;
  assign n292 = n278 ^ x85 ^ 1'b0 ;
  assign n293 = n281 ^ n278 ^ n272 ;
  assign n294 = ( n278 & n292 ) | ( n278 & ~n293 ) | ( n292 & ~n293 ) ;
  assign n295 = n294 ^ n291 ^ n281 ;
  assign n296 = n294 ^ x83 ^ 1'b0 ;
  assign n297 = ( n294 & ~n295 ) | ( n294 & n296 ) | ( ~n295 & n296 ) ;
  assign n298 = n290 ^ n287 ^ 1'b0 ;
  assign n299 = x82 | x83 ;
  assign n300 = ( n285 & ~n290 ) | ( n285 & n298 ) | ( ~n290 & n298 ) ;
  assign n301 = n299 ^ n291 ^ 1'b0 ;
  assign n302 = ( n281 & ~n291 ) | ( n281 & n301 ) | ( ~n291 & n301 ) ;
  assign n303 = x80 | x81 ;
  assign n304 = n299 | n303 ;
  assign n305 = n303 ^ n302 ^ 1'b0 ;
  assign n306 = ( n291 & ~n302 ) | ( n291 & n305 ) | ( ~n302 & n305 ) ;
  assign n307 = n287 | n304 ;
  assign n308 = ( n255 & ~n284 ) | ( n255 & n307 ) | ( ~n284 & n307 ) ;
  assign n309 = n304 ^ n300 ^ 1'b0 ;
  assign n310 = n302 ^ n297 ^ n291 ;
  assign n311 = n282 | n307 ;
  assign n312 = n297 ^ x81 ^ 1'b0 ;
  assign n313 = ( n297 & ~n310 ) | ( n297 & n312 ) | ( ~n310 & n312 ) ;
  assign n314 = n313 ^ x79 ^ 1'b0 ;
  assign n315 = n313 ^ n306 ^ n302 ;
  assign n316 = ( n313 & n314 ) | ( n313 & ~n315 ) | ( n314 & ~n315 ) ;
  assign n317 = x78 | x79 ;
  assign n318 = n317 ^ n306 ^ 1'b0 ;
  assign n319 = ( n302 & ~n306 ) | ( n302 & n318 ) | ( ~n306 & n318 ) ;
  assign n320 = n316 ^ x77 ^ 1'b0 ;
  assign n321 = ( n290 & ~n300 ) | ( n290 & n309 ) | ( ~n300 & n309 ) ;
  assign n322 = n319 ^ n316 ^ n306 ;
  assign n323 = ( n316 & n320 ) | ( n316 & ~n322 ) | ( n320 & ~n322 ) ;
  assign n324 = ( ~x67 & x68 ) | ( ~x67 & n311 ) | ( x68 & n311 ) ;
  assign n325 = ~n240 & n311 ;
  assign n326 = x67 | n324 ;
  assign n327 = ( ~x69 & x70 ) | ( ~x69 & n326 ) | ( x70 & n326 ) ;
  assign n328 = x69 | n327 ;
  assign n329 = ( ~x65 & x66 ) | ( ~x65 & n328 ) | ( x66 & n328 ) ;
  assign n330 = x65 | n329 ;
  assign n331 = x76 | x77 ;
  assign n332 = n323 ^ x75 ^ 1'b0 ;
  assign n333 = n331 ^ n319 ^ 1'b0 ;
  assign n334 = ( n306 & ~n319 ) | ( n306 & n333 ) | ( ~n319 & n333 ) ;
  assign n335 = n334 ^ n323 ^ n319 ;
  assign n336 = ( n323 & n332 ) | ( n323 & ~n335 ) | ( n332 & ~n335 ) ;
  assign n337 = x74 | x75 ;
  assign n338 = n337 ^ n334 ^ 1'b0 ;
  assign n339 = ( n319 & ~n334 ) | ( n319 & n338 ) | ( ~n334 & n338 ) ;
  assign n340 = ( ~x73 & x74 ) | ( ~x73 & n331 ) | ( x74 & n331 ) ;
  assign n341 = x73 | n340 ;
  assign n342 = ( ~x75 & x78 ) | ( ~x75 & n341 ) | ( x78 & n341 ) ;
  assign n343 = n317 | n331 ;
  assign n344 = n343 ^ n321 ^ 1'b0 ;
  assign n345 = ( n300 & ~n321 ) | ( n300 & n344 ) | ( ~n321 & n344 ) ;
  assign n346 = x72 | x73 ;
  assign n347 = n337 | n346 ;
  assign n348 = n346 ^ n339 ^ 1'b0 ;
  assign n349 = ( n334 & ~n339 ) | ( n334 & n348 ) | ( ~n339 & n348 ) ;
  assign n350 = x75 | n342 ;
  assign n351 = ( ~x71 & x72 ) | ( ~x71 & n350 ) | ( x72 & n350 ) ;
  assign n352 = n339 ^ n336 ^ n334 ;
  assign n353 = x71 | n351 ;
  assign n354 = n343 | n347 ;
  assign n355 = n347 ^ n345 ^ 1'b0 ;
  assign n356 = ( n321 & ~n345 ) | ( n321 & n355 ) | ( ~n345 & n355 ) ;
  assign n357 = x71 | n354 ;
  assign n358 = ( ~x69 & x70 ) | ( ~x69 & n353 ) | ( x70 & n353 ) ;
  assign n359 = x69 | n358 ;
  assign n360 = ( ~x64 & n330 ) | ( ~x64 & n357 ) | ( n330 & n357 ) ;
  assign n361 = n354 ^ n308 ^ 1'b0 ;
  assign n362 = x64 | n360 ;
  assign n363 = ( n284 & ~n308 ) | ( n284 & n361 ) | ( ~n308 & n361 ) ;
  assign n364 = n336 ^ x73 ^ 1'b0 ;
  assign n365 = ( ~x67 & x68 ) | ( ~x67 & n359 ) | ( x68 & n359 ) ;
  assign n366 = ( n336 & ~n352 ) | ( n336 & n364 ) | ( ~n352 & n364 ) ;
  assign n367 = x67 | n365 ;
  assign n368 = x64 | x65 ;
  assign n369 = n253 & ~n325 ;
  assign n370 = ( ~x66 & n367 ) | ( ~x66 & n368 ) | ( n367 & n368 ) ;
  assign n371 = x66 | n370 ;
  assign n372 = n371 ^ n369 ^ n325 ;
  assign n373 = ( x79 & n240 ) | ( x79 & ~n325 ) | ( n240 & ~n325 ) ;
  assign n374 = x70 | x71 ;
  assign n375 = ( ~n325 & n372 ) | ( ~n325 & n373 ) | ( n372 & n373 ) ;
  assign n376 = n374 ^ n349 ^ 1'b0 ;
  assign n377 = ( n339 & ~n349 ) | ( n339 & n376 ) | ( ~n349 & n376 ) ;
  assign n378 = n240 | n253 ;
  assign n379 = n366 ^ n349 ^ n339 ;
  assign n380 = ~n253 & n375 ;
  assign n381 = n253 | n325 ;
  assign n382 = n366 ^ x71 ^ 1'b0 ;
  assign n383 = ( n366 & ~n379 ) | ( n366 & n382 ) | ( ~n379 & n382 ) ;
  assign n384 = n383 ^ n377 ^ n349 ;
  assign n385 = n383 ^ x69 ^ 1'b0 ;
  assign n386 = ( n383 & ~n384 ) | ( n383 & n385 ) | ( ~n384 & n385 ) ;
  assign n387 = x68 | x69 ;
  assign n388 = n374 | n387 ;
  assign n389 = n387 ^ n377 ^ 1'b0 ;
  assign n390 = ( n349 & ~n377 ) | ( n349 & n389 ) | ( ~n377 & n389 ) ;
  assign n391 = n388 ^ n356 ^ 1'b0 ;
  assign n392 = ( n345 & ~n356 ) | ( n345 & n391 ) | ( ~n356 & n391 ) ;
  assign n393 = n386 ^ x67 ^ 1'b0 ;
  assign n394 = n390 ^ n386 ^ n377 ;
  assign n395 = ( n386 & n393 ) | ( n386 & ~n394 ) | ( n393 & ~n394 ) ;
  assign n396 = x66 | x67 ;
  assign n397 = n396 ^ n390 ^ 1'b0 ;
  assign n398 = ( n377 & ~n390 ) | ( n377 & n397 ) | ( ~n390 & n397 ) ;
  assign n399 = n398 ^ n368 ^ 1'b0 ;
  assign n400 = n368 | n396 ;
  assign n401 = n400 ^ n392 ^ 1'b0 ;
  assign n402 = n388 | n400 ;
  assign n403 = ( n356 & ~n392 ) | ( n356 & n401 ) | ( ~n392 & n401 ) ;
  assign n404 = n398 ^ n395 ^ n390 ;
  assign n405 = ( n390 & ~n398 ) | ( n390 & n399 ) | ( ~n398 & n399 ) ;
  assign n406 = n402 ^ n363 ^ 1'b0 ;
  assign n407 = ( n308 & ~n363 ) | ( n308 & n406 ) | ( ~n363 & n406 ) ;
  assign n408 = n395 ^ x65 ^ 1'b0 ;
  assign n409 = ( n395 & ~n404 ) | ( n395 & n408 ) | ( ~n404 & n408 ) ;
  assign n410 = n409 ^ n405 ^ n398 ;
  assign n411 = n409 ^ x63 ^ 1'b0 ;
  assign n412 = ( n409 & ~n410 ) | ( n409 & n411 ) | ( ~n410 & n411 ) ;
  assign n413 = x62 | x63 ;
  assign n414 = n413 ^ n405 ^ 1'b0 ;
  assign n415 = x60 | x61 ;
  assign n416 = ( n398 & ~n405 ) | ( n398 & n414 ) | ( ~n405 & n414 ) ;
  assign n417 = n416 ^ n415 ^ 1'b0 ;
  assign n418 = n412 ^ x61 ^ 1'b0 ;
  assign n419 = ( n405 & ~n416 ) | ( n405 & n417 ) | ( ~n416 & n417 ) ;
  assign n420 = n416 ^ n412 ^ n405 ;
  assign n421 = ( n412 & n418 ) | ( n412 & ~n420 ) | ( n418 & ~n420 ) ;
  assign n422 = n421 ^ x59 ^ 1'b0 ;
  assign n423 = n421 ^ n419 ^ n416 ;
  assign n424 = ( n421 & n422 ) | ( n421 & ~n423 ) | ( n422 & ~n423 ) ;
  assign n425 = x58 | x59 ;
  assign n426 = n425 ^ n419 ^ 1'b0 ;
  assign n427 = ( n416 & ~n419 ) | ( n416 & n426 ) | ( ~n419 & n426 ) ;
  assign n428 = n413 | n415 ;
  assign n429 = n424 ^ x57 ^ 1'b0 ;
  assign n430 = n428 ^ n403 ^ 1'b0 ;
  assign n431 = ( n392 & ~n403 ) | ( n392 & n430 ) | ( ~n403 & n430 ) ;
  assign n432 = n427 ^ n424 ^ n419 ;
  assign n433 = ( n424 & n429 ) | ( n424 & ~n432 ) | ( n429 & ~n432 ) ;
  assign n434 = x56 | x57 ;
  assign n435 = n434 ^ n427 ^ 1'b0 ;
  assign n436 = n425 | n434 ;
  assign n437 = ( n419 & ~n427 ) | ( n419 & n435 ) | ( ~n427 & n435 ) ;
  assign n438 = n437 ^ n433 ^ n427 ;
  assign n439 = n433 ^ x55 ^ 1'b0 ;
  assign n440 = ( n433 & ~n438 ) | ( n433 & n439 ) | ( ~n438 & n439 ) ;
  assign n441 = x54 | x55 ;
  assign n442 = n441 ^ n437 ^ 1'b0 ;
  assign n443 = ( n427 & ~n437 ) | ( n427 & n442 ) | ( ~n437 & n442 ) ;
  assign n444 = n428 | n436 ;
  assign n445 = n444 ^ n407 ^ 1'b0 ;
  assign n446 = ( n363 & ~n407 ) | ( n363 & n445 ) | ( ~n407 & n445 ) ;
  assign n447 = x52 | x53 ;
  assign n448 = n441 | n447 ;
  assign n449 = n447 ^ n443 ^ 1'b0 ;
  assign n450 = n436 ^ n431 ^ 1'b0 ;
  assign n451 = ( n437 & ~n443 ) | ( n437 & n449 ) | ( ~n443 & n449 ) ;
  assign n452 = n443 ^ n440 ^ n437 ;
  assign n453 = ( n403 & ~n431 ) | ( n403 & n450 ) | ( ~n431 & n450 ) ;
  assign n454 = n453 ^ n448 ^ 1'b0 ;
  assign n455 = ( n431 & ~n453 ) | ( n431 & n454 ) | ( ~n453 & n454 ) ;
  assign n456 = n440 ^ x53 ^ 1'b0 ;
  assign n457 = ( n440 & ~n452 ) | ( n440 & n456 ) | ( ~n452 & n456 ) ;
  assign n458 = n457 ^ x51 ^ 1'b0 ;
  assign n459 = n457 ^ n451 ^ n443 ;
  assign n460 = ( n457 & n458 ) | ( n457 & ~n459 ) | ( n458 & ~n459 ) ;
  assign n461 = x50 | x51 ;
  assign n462 = n461 ^ n451 ^ 1'b0 ;
  assign n463 = ( n443 & ~n451 ) | ( n443 & n462 ) | ( ~n451 & n462 ) ;
  assign n464 = x48 | x49 ;
  assign n465 = n461 | n464 ;
  assign n466 = n464 ^ n463 ^ 1'b0 ;
  assign n467 = n448 | n465 ;
  assign n468 = ( n451 & ~n463 ) | ( n451 & n466 ) | ( ~n463 & n466 ) ;
  assign n469 = n465 ^ n455 ^ 1'b0 ;
  assign n470 = n463 ^ n460 ^ n451 ;
  assign n471 = n444 | n467 ;
  assign n472 = n467 ^ n446 ^ 1'b0 ;
  assign n473 = ( n407 & ~n446 ) | ( n407 & n472 ) | ( ~n446 & n472 ) ;
  assign n474 = n460 ^ x49 ^ 1'b0 ;
  assign n475 = ( n460 & ~n470 ) | ( n460 & n474 ) | ( ~n470 & n474 ) ;
  assign n476 = ( n453 & ~n455 ) | ( n453 & n469 ) | ( ~n455 & n469 ) ;
  assign n477 = n475 ^ x47 ^ 1'b0 ;
  assign n478 = n475 ^ n468 ^ n463 ;
  assign n479 = ( n475 & n477 ) | ( n475 & ~n478 ) | ( n477 & ~n478 ) ;
  assign n480 = ( ~n380 & n381 ) | ( ~n380 & n471 ) | ( n381 & n471 ) ;
  assign n481 = x46 | x47 ;
  assign n482 = x44 | x45 ;
  assign n483 = n479 ^ x45 ^ 1'b0 ;
  assign n484 = n481 ^ n468 ^ 1'b0 ;
  assign n485 = ( n463 & ~n468 ) | ( n463 & n484 ) | ( ~n468 & n484 ) ;
  assign n486 = n485 ^ n482 ^ 1'b0 ;
  assign n487 = ( n468 & ~n485 ) | ( n468 & n486 ) | ( ~n485 & n486 ) ;
  assign n488 = n485 ^ n479 ^ n468 ;
  assign n489 = ( n479 & n483 ) | ( n479 & ~n488 ) | ( n483 & ~n488 ) ;
  assign n490 = n489 ^ x43 ^ 1'b0 ;
  assign n491 = n489 ^ n487 ^ n485 ;
  assign n492 = ( n489 & n490 ) | ( n489 & ~n491 ) | ( n490 & ~n491 ) ;
  assign n493 = x42 | x43 ;
  assign n494 = n493 ^ n487 ^ 1'b0 ;
  assign n495 = ( n485 & ~n487 ) | ( n485 & n494 ) | ( ~n487 & n494 ) ;
  assign n496 = n481 | n482 ;
  assign n497 = n492 ^ x41 ^ 1'b0 ;
  assign n498 = n496 ^ n476 ^ 1'b0 ;
  assign n499 = ( n455 & ~n476 ) | ( n455 & n498 ) | ( ~n476 & n498 ) ;
  assign n500 = x40 | x41 ;
  assign n501 = n493 | n500 ;
  assign n502 = n500 ^ n495 ^ 1'b0 ;
  assign n503 = ( n487 & ~n495 ) | ( n487 & n502 ) | ( ~n495 & n502 ) ;
  assign n504 = n495 ^ n492 ^ n487 ;
  assign n505 = ( n492 & n497 ) | ( n492 & ~n504 ) | ( n497 & ~n504 ) ;
  assign n506 = n496 | n501 ;
  assign n507 = x38 | x39 ;
  assign n508 = n507 ^ n503 ^ 1'b0 ;
  assign n509 = ( n495 & ~n503 ) | ( n495 & n508 ) | ( ~n503 & n508 ) ;
  assign n510 = n501 ^ n499 ^ 1'b0 ;
  assign n511 = ( n476 & ~n499 ) | ( n476 & n510 ) | ( ~n499 & n510 ) ;
  assign n512 = n505 ^ x39 ^ 1'b0 ;
  assign n513 = n505 ^ n503 ^ n495 ;
  assign n514 = ( n505 & n512 ) | ( n505 & ~n513 ) | ( n512 & ~n513 ) ;
  assign n515 = n506 ^ n473 ^ 1'b0 ;
  assign n516 = x36 | x37 ;
  assign n517 = n507 | n516 ;
  assign n518 = n516 ^ n509 ^ 1'b0 ;
  assign n519 = ( n446 & ~n473 ) | ( n446 & n515 ) | ( ~n473 & n515 ) ;
  assign n520 = n514 ^ n509 ^ n503 ;
  assign n521 = ( n503 & ~n509 ) | ( n503 & n518 ) | ( ~n509 & n518 ) ;
  assign n522 = n514 ^ x37 ^ 1'b0 ;
  assign n523 = ( n514 & ~n520 ) | ( n514 & n522 ) | ( ~n520 & n522 ) ;
  assign n524 = n517 ^ n511 ^ 1'b0 ;
  assign n525 = ( n499 & ~n511 ) | ( n499 & n524 ) | ( ~n511 & n524 ) ;
  assign n526 = n523 ^ n521 ^ n509 ;
  assign n527 = n523 ^ x35 ^ 1'b0 ;
  assign n528 = ( n523 & ~n526 ) | ( n523 & n527 ) | ( ~n526 & n527 ) ;
  assign n529 = x34 | x35 ;
  assign n530 = n529 ^ n521 ^ 1'b0 ;
  assign n531 = ( n509 & ~n521 ) | ( n509 & n530 ) | ( ~n521 & n530 ) ;
  assign n532 = x32 | x33 ;
  assign n533 = n529 | n532 ;
  assign n534 = n517 | n533 ;
  assign n535 = n533 ^ n525 ^ 1'b0 ;
  assign n536 = n532 ^ n531 ^ 1'b0 ;
  assign n537 = n506 | n534 ;
  assign n538 = n471 | n537 ;
  assign n539 = ( n511 & ~n525 ) | ( n511 & n535 ) | ( ~n525 & n535 ) ;
  assign n540 = n528 ^ x33 ^ 1'b0 ;
  assign n541 = ( n521 & ~n531 ) | ( n521 & n536 ) | ( ~n531 & n536 ) ;
  assign n542 = n531 ^ n528 ^ n521 ;
  assign n543 = ( n528 & n540 ) | ( n528 & ~n542 ) | ( n540 & ~n542 ) ;
  assign n544 = n543 ^ n541 ^ n531 ;
  assign n545 = n378 | n538 ;
  assign n546 = ( ~n362 & n378 ) | ( ~n362 & n545 ) | ( n378 & n545 ) ;
  assign n547 = n362 | n378 ;
  assign n548 = n534 ^ n519 ^ 1'b0 ;
  assign n549 = ( n473 & ~n519 ) | ( n473 & n548 ) | ( ~n519 & n548 ) ;
  assign n550 = n543 ^ x31 ^ 1'b0 ;
  assign n551 = ( n543 & ~n544 ) | ( n543 & n550 ) | ( ~n544 & n550 ) ;
  assign n552 = x30 | x31 ;
  assign n553 = x28 | x29 ;
  assign n554 = n552 ^ n541 ^ 1'b0 ;
  assign n555 = ( n531 & ~n541 ) | ( n531 & n554 ) | ( ~n541 & n554 ) ;
  assign n556 = n555 ^ n553 ^ 1'b0 ;
  assign n557 = ( n541 & ~n555 ) | ( n541 & n556 ) | ( ~n555 & n556 ) ;
  assign n558 = n555 ^ n551 ^ n541 ;
  assign n559 = n551 ^ x29 ^ 1'b0 ;
  assign n560 = ( n551 & ~n558 ) | ( n551 & n559 ) | ( ~n558 & n559 ) ;
  assign n561 = n560 ^ n557 ^ n555 ;
  assign n562 = n560 ^ x27 ^ 1'b0 ;
  assign n563 = ( n560 & ~n561 ) | ( n560 & n562 ) | ( ~n561 & n562 ) ;
  assign n564 = x26 | x27 ;
  assign n565 = n564 ^ n557 ^ 1'b0 ;
  assign n566 = n552 | n553 ;
  assign n567 = ( n555 & ~n557 ) | ( n555 & n565 ) | ( ~n557 & n565 ) ;
  assign n568 = x24 | x25 ;
  assign n569 = n564 | n568 ;
  assign n570 = n568 ^ n567 ^ 1'b0 ;
  assign n571 = n563 ^ x25 ^ 1'b0 ;
  assign n572 = ( n557 & ~n567 ) | ( n557 & n570 ) | ( ~n567 & n570 ) ;
  assign n573 = n567 ^ n563 ^ n557 ;
  assign n574 = ( n563 & n571 ) | ( n563 & ~n573 ) | ( n571 & ~n573 ) ;
  assign n575 = n574 ^ x23 ^ 1'b0 ;
  assign n576 = n574 ^ n572 ^ n567 ;
  assign n577 = ( n574 & n575 ) | ( n574 & ~n576 ) | ( n575 & ~n576 ) ;
  assign n578 = x22 | x23 ;
  assign n579 = n578 ^ n572 ^ 1'b0 ;
  assign n580 = ( n567 & ~n572 ) | ( n567 & n579 ) | ( ~n572 & n579 ) ;
  assign n581 = n566 ^ n539 ^ 1'b0 ;
  assign n582 = ( n525 & ~n539 ) | ( n525 & n581 ) | ( ~n539 & n581 ) ;
  assign n583 = n582 ^ n569 ^ 1'b0 ;
  assign n584 = ( n539 & ~n582 ) | ( n539 & n583 ) | ( ~n582 & n583 ) ;
  assign n585 = x20 | x21 ;
  assign n586 = n578 | n585 ;
  assign n587 = n585 ^ n580 ^ 1'b0 ;
  assign n588 = ( n572 & ~n580 ) | ( n572 & n587 ) | ( ~n580 & n587 ) ;
  assign n589 = n566 | n569 ;
  assign n590 = n577 ^ x21 ^ 1'b0 ;
  assign n591 = n580 ^ n577 ^ n572 ;
  assign n592 = ( n577 & n590 ) | ( n577 & ~n591 ) | ( n590 & ~n591 ) ;
  assign n593 = n586 ^ n584 ^ 1'b0 ;
  assign n594 = ( n582 & ~n584 ) | ( n582 & n593 ) | ( ~n584 & n593 ) ;
  assign n595 = n589 ^ n549 ^ 1'b0 ;
  assign n596 = ( n519 & ~n549 ) | ( n519 & n595 ) | ( ~n549 & n595 ) ;
  assign n597 = n592 ^ n588 ^ n580 ;
  assign n598 = n592 ^ x19 ^ 1'b0 ;
  assign n599 = ( n592 & ~n597 ) | ( n592 & n598 ) | ( ~n597 & n598 ) ;
  assign n600 = x18 | x19 ;
  assign n601 = n600 ^ n588 ^ 1'b0 ;
  assign n602 = ( n580 & ~n588 ) | ( n580 & n601 ) | ( ~n588 & n601 ) ;
  assign n603 = x16 | x17 ;
  assign n604 = n600 | n603 ;
  assign n605 = n586 | n604 ;
  assign n606 = n603 ^ n602 ^ 1'b0 ;
  assign n607 = n604 ^ n594 ^ 1'b0 ;
  assign n608 = ( n584 & ~n594 ) | ( n584 & n607 ) | ( ~n594 & n607 ) ;
  assign n609 = ( n588 & ~n602 ) | ( n588 & n606 ) | ( ~n602 & n606 ) ;
  assign n610 = n602 ^ n599 ^ n588 ;
  assign n611 = n599 ^ x17 ^ 1'b0 ;
  assign n612 = ( n599 & ~n610 ) | ( n599 & n611 ) | ( ~n610 & n611 ) ;
  assign n613 = n589 | n605 ;
  assign n614 = n537 & n613 ;
  assign n615 = n614 ^ n613 ^ n480 ;
  assign n616 = ( ~n380 & n480 ) | ( ~n380 & n615 ) | ( n480 & n615 ) ;
  assign n617 = n612 ^ x15 ^ 1'b0 ;
  assign n618 = n612 ^ n609 ^ n602 ;
  assign n619 = ( n612 & n617 ) | ( n612 & ~n618 ) | ( n617 & ~n618 ) ;
  assign n620 = x14 | x15 ;
  assign n621 = n620 ^ n609 ^ 1'b0 ;
  assign n622 = ( n602 & ~n609 ) | ( n602 & n621 ) | ( ~n609 & n621 ) ;
  assign n623 = n619 ^ x13 ^ 1'b0 ;
  assign n624 = x12 | x13 ;
  assign n625 = n620 | n624 ;
  assign n626 = n624 ^ n622 ^ 1'b0 ;
  assign n627 = ( n609 & ~n622 ) | ( n609 & n626 ) | ( ~n622 & n626 ) ;
  assign n628 = n622 ^ n619 ^ n609 ;
  assign n629 = ( n619 & n623 ) | ( n619 & ~n628 ) | ( n623 & ~n628 ) ;
  assign n630 = n629 ^ x11 ^ 1'b0 ;
  assign n631 = n629 ^ n627 ^ n622 ;
  assign n632 = ( n629 & n630 ) | ( n629 & ~n631 ) | ( n630 & ~n631 ) ;
  assign n633 = n625 ^ n608 ^ 1'b0 ;
  assign n634 = x10 | x11 ;
  assign n635 = ( n594 & ~n608 ) | ( n594 & n633 ) | ( ~n608 & n633 ) ;
  assign n636 = n634 ^ n627 ^ 1'b0 ;
  assign n637 = ( n622 & ~n627 ) | ( n622 & n636 ) | ( ~n627 & n636 ) ;
  assign n638 = x8 | x9 ;
  assign n639 = n634 | n638 ;
  assign n640 = n625 | n639 ;
  assign n641 = n605 & n640 ;
  assign n642 = n641 ^ n640 ^ n596 ;
  assign n643 = ( ~n549 & n596 ) | ( ~n549 & n642 ) | ( n596 & n642 ) ;
  assign n644 = n632 ^ x9 ^ 1'b0 ;
  assign n645 = n638 ^ n637 ^ 1'b0 ;
  assign n646 = ( n627 & ~n637 ) | ( n627 & n645 ) | ( ~n637 & n645 ) ;
  assign n647 = n637 ^ n632 ^ n627 ;
  assign n648 = ( n632 & n644 ) | ( n632 & ~n647 ) | ( n644 & ~n647 ) ;
  assign n649 = x6 | x7 ;
  assign n650 = x4 | x5 ;
  assign n651 = n649 | n650 ;
  assign n652 = ~n639 & n651 ;
  assign n653 = n613 | n651 ;
  assign n654 = x2 | x3 ;
  assign n655 = n652 ^ n635 ^ 1'b0 ;
  assign n656 = n650 & n654 ;
  assign n657 = n649 ^ n646 ^ 1'b0 ;
  assign n658 = ( n637 & ~n646 ) | ( n637 & n657 ) | ( ~n646 & n657 ) ;
  assign n659 = n658 ^ n656 ^ n654 ;
  assign n660 = n640 | n654 ;
  assign n661 = x0 | x1 ;
  assign n662 = ( ~n547 & n660 ) | ( ~n547 & n661 ) | ( n660 & n661 ) ;
  assign n663 = x1 & ~x2 ;
  assign n664 = ( ~n646 & n658 ) | ( ~n646 & n659 ) | ( n658 & n659 ) ;
  assign n665 = n648 ^ n646 ^ n637 ;
  assign n666 = ( ~n608 & n635 ) | ( ~n608 & n655 ) | ( n635 & n655 ) ;
  assign n667 = x3 & ~n663 ;
  assign n668 = n648 ^ x7 ^ 1'b0 ;
  assign n669 = n547 | n662 ;
  assign n670 = ( ~n538 & n653 ) | ( ~n538 & n669 ) | ( n653 & n669 ) ;
  assign n671 = n538 | n670 ;
  assign n672 = ( n648 & ~n665 ) | ( n648 & n668 ) | ( ~n665 & n668 ) ;
  assign n673 = n672 ^ n658 ^ n646 ;
  assign n674 = n673 ^ x4 ^ 1'b0 ;
  assign n675 = n672 ^ x5 ^ 1'b0 ;
  assign n676 = ( n672 & ~n673 ) | ( n672 & n675 ) | ( ~n673 & n675 ) ;
  assign n677 = ( n673 & n674 ) | ( n673 & ~n676 ) | ( n674 & ~n676 ) ;
  assign n678 = n677 ^ n667 ^ n663 ;
  assign n679 = ( n676 & ~n677 ) | ( n676 & n678 ) | ( ~n677 & n678 ) ;
  assign y0 = n679 ;
  assign y1 = n664 ;
  assign y2 = n666 ;
  assign y3 = n643 ;
  assign y4 = n616 ;
  assign y5 = n546 ;
  assign y6 = n547 ;
  assign y7 = n671 ;
endmodule
